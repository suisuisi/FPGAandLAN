

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
grYpUA5jzoYp1LlWmdZ2ALEfyb0iZaBlbu2Jn5TWbislv0ePefGNtLrxAsy9+neVRtGKqzd/weQY
1GDOlCD3sw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jJRJFGl+freuRUOkHi4uiJXF1ZSDXCZnSp7sify5hay8gI8WQ5QHE0Kl1tU1VRdOD+ovbKr3K+cS
UqWpgUyeIHMS2fFsOi6SAu6Aoshxr0Vl9PE57JGCyWYxhIS/bFj42inspCVQCybe04fBzJMNWaUp
2qePZYRz32xbymT2jPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu6th/stm+M5ynB/TKpquW8ZkolQD8eNSgYHhWrx1S0Oj+qDq3ifkyYP979H5aZBSsmi9nhkBeP5
00SMQNL9WZH3DTym/hO1AOEB/vZQ4iH5QuRFIKccEqDq2JtY6+UDXXKzO/1rIfmarsHX8ltlRTV/
zcfaeOmCAj7ywQc9UqYmky4qV8fErTo0+Sdz/lesSXUkxz2bi3RdkWlaTaVx6gglEIQd+UT3ZYt3
+UGswd7jIOxS6vlCnneyc3neS690RMPIIoNUnxysnaeZZUGvdfZpjktfag6rjQ59uaAGWliO4MMi
6ToA8bqievgo9dlWIHZ7qHH63+ZPGm4+ACmZLw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
anxX3tP+OSA4f+Zz3xRPWpNr0NFYOEkjWa+yDywi9ewNNEKmVmuybI2vuUNyxHHqdZuNWtw1fzH+
LvHMudDHSvrqUXO0i+yPr/b1uULww82dKZJhMTouZXfSBUYYR2R6eOUHlkc2mpuJW1b0Yfgqe/lL
U2cURbnRhzUDfX4a8/KZsget317eHUxMWntDUJjMnFKpxAe6rTs57ljr+47CKoyVApxpFRtXyva0
iIrl61ypfwevW1NM+dbuq0A2ep4qpKF3QXqu+5quZRKiS9wqmBIWbGIwWUFzi9jVuDlWbiy7K2/8
HWrhgAyLQfd3aizqZge9Kid8TFg/tOAzl3/Dig==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hfg0jhNUSwZoyKs+dkGwZfuOuLOYxt8dUSYFBsXNe53zJQUTW2+PTKtB4x0Xb2iLN7gmIGI0MkTa
VnwntAtFN20kw1KSsvMMJ5tmSswwrxvHJwEQEUQ97ZGqSWO2GHL6Y1M+TGniM4GhJ4MqrJ9nz3bJ
lDbNWHgjFGsf/h3qT5IiPslEewuncdt89+9yjAvcmXEyKAI2nU9sb2+Z/dYcbWohVAJhqZIShNET
j4MueDXbjuGAb3rviJH30Ms0ITe492AtvNh8bbtTcCumEGRwdxdBrBtudooM4fhp1QOulK1MlV70
8clOJrGF2872zCxai4LigCCBOk0uSW3ObDKbXg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SbPUQ56CmxNuuFeULNmdtP4VI25yIuTqRpQZv4fdI4ab2e9QChHgoTeL8pKVO9WcuhlNTx166GsZ
+J7LQgSi3dQSR++PcS3u1e//zfZcwXePmh5ndXtuNKSeOT1YlsZMy0NFnCR74oDcXIAWozlvfa3H
+Ha8zpAYNJlEcIxIlN8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iBM86j8TSZyV5DU0rYA8Io0mzpNhxgzW55YqzBpIYOLzQUiY8G8WAdKhnnqwoz2tPjopVirg1TR5
tvZKebOq9UC6KFo7vKxpOX57N0cp4fFPLdWGp3bfCI0YVxBdZnmmB4Oc+YtxYdI6e+BC82GkMG6d
gVuqFuf9L0mulL+yXuTTt2uiDajwZIcjyq11UByNJFKgZWndCJNV+FkUL21qP0t0BgzJPx1vq9GI
Xcdhwmaqi5DH7ZSxtXWYHzXgMDV5w1iNgDI3RX7uYUR/uvXUFc8tvCukL4SxyVDekPuhO3EOq7lP
gm4n/MB66m+/WkJd04R1OsrCyFsGEkoFVCl47w==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TDm/CaHzF2sRlkHDDHosS/V53FzLYAEPesCrg1+oRNDDuRD9Xb5WpyqcNNNidE9joaps4c7lrYCD
3nRf5x+Z12x0YPF7kaiPnyDbXkFRv6Qy+JTaRUXeoTs54W+jPqxDrL1x6Wv9yIyFxShptBbnNkVI
e+UMuxDyxwcdq81KmTCZc+NgWtBB1VzY7ity43L6Zk/6njjEpAsUd275HuhcP4JW4NFW1TZDaNnF
Cww6OTyrgEG5hWZR86AzBS7yjfi5vJjN94IDbGHICM+1BbHZNAAylzDKaXvbNdWIsQbt3lRVnU+z
u9i9+X1Drqb7MWsOo8jYLXDlib7Gpm56+SqMOg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133696)
`protect data_block
iN4N2HEk3aD4Z34cQXMAABEdk9ZWVivZoeSyOzFDxJB++fI3uKggOpY8u1WT7xc9QwGd5623b64f
avI4AS5vHWLm94bnXGPEDr/k+tY9N50w7ft+SDS3BVuwzFIlmAxyIFEsEoPT5f1d6AYoeCiypOfd
4bD/vzzB/CYZ3Y+mnnViocGEMu82WQLCNrq9d3A9pVKuJ/4FGVhPhpK95hhNditSDzvMckujT6OM
ZM/FYSpErjIS5555jKGib737ISJ9MkeWsW5mLj7ptPzYpcutRLlErsqN7VyHMmCguZPONKY7FPzY
/V9Jc619l/jrYw/0Cxa69ClZLK8vJtUm5VgHrAaSu7Y1lkxi07zuRlcWQJUVVRCu5xesEXC93PAY
/gbMDTZo1dftPiO/ibbXSXXNEu/BRcIKylJlzSP0FZJ271MUEwz31ra8HusQ2PdvkTSOK0SHbvDz
Sqfbhn8iRC1qBpO2F3cNyR4gPGMsSavPjmC89qri2xttLdGbYF2xmU8tPPzPfJVFqAE+481b4gFV
fdA9MNrbb/P+g5ce5QYqlhxiD0gXIpwteULg4Z6+C3F88pj9USILHmW90+zIz+wV8KZKo1OluUQ7
ol0Tm6Tf6FH6O8+3IPZVxF3RVkwHojSHVyZN+OAn6Sgfz0QRN7MhaqKpPQFoQyI0F31pW4IfQw3x
LBED98zHjTMqkToLR7jNU8yyqlbFc5EPcD+gJ1ZV9W4CU+YjcLWNqPcTbGag7ZVyyIn+hhuRb6t1
YGQ+MdNKnXrQbkvrXbdbJ8XrMvrR4Cjknais/sIzLaI7LuNbh0DBQQHq2XG+Lct1kYg4NGcYUuBg
aBCk5fo72OJZwo6tz4c1cZcsNR7wXG0vKvXq8nyd8lM+BKaeCfpRboISEvJsG+q0F/jhHq8Z+V4m
ge4dFqWxHSQV3X4IFJqnaoS0S40kIO8wGqwqm/0kNdSY6yxrfQJLQfQa/cBdLBq4Evc/SlSKr7Iz
Jrm1skOarvzjPnncY822rs4YZRl0s2te0gDI+RSef1ydfWN8Hn4dZdOwhdSiiuGhwfiBQr23zrv9
V5Y6yhEG7vZfK6p3cwtt1l37Cc2NfvQsf6cGjoh+rLaIgJ8fdH+jyLISX+z1C6Kef8uTQyCaCCoW
SJaQxmpvyu0sl8YCK1xrsRJd0yWOYNTOBMY7pPasOJuSw43OqfQJ/HzSCEtAbh9PraudonlmXywn
YiXS44+HJ0dZ/Zl19MI7tc/CgAHBr3bUkOak0lh8mn6Yt+LIRjJozI3YxsuYt76Wjne6o78ZHdu8
YepYa45ARtxf2seIEXcSoTrU0z2BSMCUfMngYmRWzUJ8I/NhFsMf21jU+P3X2NYJqk6tZhXPbdf7
auq+QLIw8xz7qnGvS2FTBrAm6NPA3sQG5R4FQmkORj0UMTTojpyrZJfi3u9e8UlOA0zyJsmqg07H
AuThxkcB21LMXf+xTIpHResvC0gixR+FjejfMiBaeXRNMVf8xunuAcq9YvORUgQ+dZmESEGGrhOC
p4hevc8nZ/pN+n4CRoOGQ0zbduzBcIe9E35TKQpurGGkQH/RHfaOK4kfG4whpG8wWuy/M0d3iqVO
zsgyiCcwbK3er/9wWPIHT2rZynlF+T8nZ50mZyp/WmnXTWn0r8OnawJTrUABqd5LawMuwh6CIF8N
7vyPbhCZgeQ2WD4Jz8KkbCk9TGmTb3sS2LFqOUyEUfTp/Ojh0sWBSrt+WInSF3HN1+GizgN/dKNc
3itlpQ2Ki1OcsSQKEQ+Nyw74JbpxcN5jyuhNbbx5kniJN0qUu2qHKhm1dynmhv+tm2hMOSSvdUeH
sohiM4rG+lSkGgEw9XLK79ioaLlKGYKnx2ubH1zOgZ0NpwoDT4o7DX1F5w694ziH3raODpX9raeL
VUOe/mneLkMR1IHTUe1mUv4/UszVl1ttEWFV5VNkKBRLHeC4J0t5tSQWZErMsFk2ftp2W7pg28lD
U7DVZQO6ZnGfuLX1NAQCWUdo3EXOgJkrMOSvIov/nXmDPkPNcQfUo/Nv5m4YOJX9XH2qTEeOTq0o
URXks8Lh0EMcOYMpZkxAuPhHbZRQt5ak3PlXIVAj4JFHxPZZHIVjrM1UBkv7uukBoSFvY2FK0oP/
FOqsmpL+hD0Oeds2QcUEHyzivYQUBB46HZCU6UefeUe0l8p9Qu6gU7CV7NyFP3MvtN9IkgdlkDdj
McoWWGGu2vf/ryRK9dbyy1BEeZeIlP4PlMN94eI4ESpZ3JExUjxd47HqO+W4V637QPD250TTU0jz
ydsMTuIOqTTIIKT09VQ6sjQ6iydkGTqP5xvVx6jNkX9LElkxmneWgZ8pszCKm+oUwRP50gzcHBKk
c5GQGwGTiFCjd7F/VQFZj0gNUPcyLk9Oocq9IV1h0/gxdrL+kVh2/CrslG2zQMfmoiv/qhIJFUWm
e2clc2fAgUj20bwvqvjokmyX5tLytP1DlM5ay5i6VfiGRtxK4xuUFW8xcJ+LXcCjleyiIv2jc5qa
jfGetEILgvacPCt3ddjgyd7zIYt106J1gW3GyILMlA8qyy9RQJVUil+1whd/s//flzLt05h8jLU7
upeGy9IzvKxZf9K/VPbUahE9Go+6kcs6aP3xk6WSJ77tz/tDwKY6Mb1DpPDXGtnm/wh9vvfmYuKm
A2N9xX6QtbcyEpOhaPo+vG6zrHVBSfjMk5rbQzpwyVCNlRc+6GAdHHNWEgIL6WOLiqAl/LOkBtvV
DM5zpB4VLV/awv+A91IioGTkN87+H4qoED4uh0YWgd2kGNajL+TlEqv3NBIcryI7nQFC1ikVeQFf
Es869lvNNnsrFKXPMDGQhaD+tSD7tScmksOxjHf97Utvhlak3NYpISsHz5WJ0n8PxnqN4ZAiAPF6
yUR/r4Z/g88dFExuzKOWC0XskiJJ2BHNm9kzCifETCwbi+5slALVbIUyNSHb66tym7YkU4nL044p
HHR+htKhQba2fePhmpvW828NNLPDyCZYY4Ec9uqUoTUF0/zx4HVK+GoOsXD8yunHOq7n3NcAJK+P
+MBBUV/d8AAA23JElRRdlN8wHV8sw3aSeqUS65wocUu1xXooBZjigutvF7a3MfCFZumzMH24hoaq
8HCyMPH7q38rk3Ekx3V2Eq7Azk+6ck397fWc6ud0tHLk45GhupBpc/L/CdFEMk1Vj4rCkPQr8mGH
Aa2dYxuqR0o//IUGeZhQHOX+ffusZLhRw3EnC6sU+fEz8bi4nfS9YbPigGW+YxjAJ0v2tIjI+AYh
eeUua2sobzYnzQCclgtoUn8h72Jgpy0TfVabPO/arFaksqhy8pdCITumlKwMguqRSgGRxpxwYnbN
TxSmQ0qNn/H1KWsM8e2Du6VIphJIDl1aU8n5HI9DqTCOl8fFv8/hNelwkTiUP6bx61V+uzSTZVeg
nSECckUCCr5zNayH74aM5mfdt+ejOqXyCjmXddxkfHk5J6dsBHWrBMCtJ3WgHf2Q/8gKL4z3u3Pc
HDjKaF7Z3hM1DUKcs3ljmE+xvxbZWCnDGD75qTqoY+doa2+RUts7Tp3C2L+nk7e4BJVmXj0AMu+a
8FukkbQxk1HcTk6t71qoMPE71YGI2EKgDAoksNGnvoo6T61qtfenTbMYPaLmt2J5CsowSH/bo/2I
xvKvh+SkZ5c8KPKulPuNfaYnaAEJT8X/m8T7T2slrEwqdANdrzYELiAhuudibjDPAAXaZETNsJ9A
0LGA8XcCbBKcapfOBLTd0DMgpw9Wf283RBrkGIMj1N4oYu1Syk3GmsqTVJw6cQiA4mq2e+gcl/JL
XmxsfiIMK6efbUqTwU+g2KYjetaGgaCgzb8SEJ1t+XjAp62okq0FZ2epT3oEhzM87AAJ9iheDhqs
6KLm3xA9NYs0NINmJ880vzzZGauOhc/o8XzWvJSjL/cIsC7/pdsS9msJ60+7pKFfDEO0puxHFEcf
SkaEciKEH0Acyb1mkHGj3CS86vJMysMMrFCDZbvvXnOUtpoKV4oPmJI8NWWemnuuilErKiNwlIhH
4WnhiI6ks3EkFkxgYBFVOOJ9gcQz7XzA+eYui0/hYW9vwbIuC0b4mGyOwKUNV57zssP0vnWkuuqj
D4LEa9mUTM2CeMcdoGJUn8eXY4ktkovuo36FniRqd2UU/SMtAaAbCYdS9N7c6dWcNOgycmD330p9
UnlU0Y2Rf9rBujeKKRXxET/svTQ6yFvNgF2IdHg+EdW7mIh3GxJ5QNrjodghh3KM363MAN1uX65m
und7uU80HKawXz3rE/k6Jpq9hChwx16JUFfA7j1f4L6ZI3YrLd2L/i2PxhOdvc5CwIrMch3ClXd3
/7EWLQSFv2wRqqWrZZ5F+qmeTc3mDiNFlACX8lr0rktcZZqZeQn2siiOtF3CXF5NACZi3WH/kcgA
jQblT5XoGzh/iLb7TvARheHZC2B5EXR/JrmIvWwtZKwvpeqaX83wzdh0LZw+OhtoueA7TElJi1J6
n7nJzqWW7M0UYXD0MZMHWx91i91gSSYLQXsU/Up9Gz4X/y1e1fdQcQ0NS8IkPf1K1JQJpfGjH/te
fzkpT1aqdowT+FCZPVGV4XwZN28YMzzMjRnEdOQNSJRU4SKoZvIBTJn8BbxjQRVEVpile4PggA2W
P8KwY+NL0SsVT0n3ugSDfVcqC3IDHBZmLjpSIFZavUHqiSWXN2Pm6OHCH/Dp6pj/JsAA7jmCsyrN
W0q5CRRT1cPUFA72dtoqwoBkV+YJmKg6Z/efvb6BZgj4NtjMMZbOSXpVRLlH1EUi2YiSyGE30qnI
ZPKuBXE9zqqcrIxnBnjzH+UxyTz/sb4OSkWIa/sLEZlbNWkRcpNcVYEK/69tTyW6gjhRqgM6z2nM
t2f1/9lQ4lq6eYrToasH6xKHCfWKERdSvyIZIilY82utTbiuXccp9iv/KZTiaHC2agbi4oGVBftA
jjwAOez/BQz7mRcDKpa+ERwJJcQF80uQDVjQd+k1AAnW8M3Bn6IQZYydexPD9NnTbKIZ0kwvOkbd
elNQSnL4UmkimLCs5XfMXFbMB+L8y1Q1f5HKvAskEckv3ZHpBnzIue7aG+bEpaQKYkCOClFvQhHw
+lZvvlK1MPTwMDSkqAbjR+vxKcJ1IUxR7TarGYDD07poLtHL4KHhIqrJVnID1XlbE+2cc1XJVn+U
urAtwPYj94dplJcnyugq0++sCV/m4HJaHDgz4GWiyOm68DO+FbEykKKaI0c4hbznRN63LuV0rMXz
FAb8DlGSj9QdJUygnfRESPociuf9/hpsD3MMECcTmyLbpog9ksXsXAP8ZhypzgOrlKMopw7Sypbe
SHuMdtvpfuZknHNFgzhUo10bQ1LybOn62L2lTBsr8iX4S4TOwWAAlU2QT1mmUsqgDjShNvjGhv5C
xCXrk3b7CP4iuc9b/9pp6sMeIMTicpETr3Tk2uyqkTUVJ2M+0Rf9JftCR4VbMIGB+L5mvwjC0QFU
ooUEs0adlNQ3U79b+Ne80DYSuMyAeM/ZE1sX6SeujZEjqOJhDJatYKkLu6nIGo54WWfg6fg4gMuK
20EolCUjND2/ZXEEtILD5J65QynxnRRNXy3rYA9SLYbLjyeoHJIMDzOjM4qW4caPvKMe3vQbEgyl
GVNMFepf7AjYYRgboS1PbNvkXrFr0S4Okwu3poF+vJfttLPmshFoTfpK7GAxz2xD/0B6Gu1K28+Y
o3vS02QU8EdwN+p2d2RdLo1TKlc4KKu5MJwVQWrpNKe/rRD7xqccognWAoUlZVSKO8kavvi2h/Ua
1su9X+OqECkAUdeP7Gel+T/OQg1PgINUIzUzWhFHmSipPDoQJTXbynssSJgk29RyeT/+TV7BC7nQ
luPSQUDEzYEp50xYZua3V71CuAxWcAf6L+4hT+zQmR532NjHNqvMo6AaMB/tz4lAg2QO7YNn0iZK
4DMPzvbZKXTPjQEs1CE0dbqnJ4nKSW+lucUp5dVoqsyfOW6jYylDOnhIpV8xQxy+O+pGKO3MEdQp
IjIxX/JmeYLAQYwxAFNtbDabPtEyazlLGQa+wsv7TpNqX5fKleRL5SXGzGtdaBzFU94ExdMZaLIO
U0tAygYXmhVMd+E9EAtx6jziF7Q4sfExYNIDBF/NKF70OQ7ApEqlj21Vh1Sz8QB1LOQuu6mCEeSM
Q8W0tCZ286s/BsqFlDmG5sweHQ3yrEXmziiN8wcGoCFhBlFCXwcddA13ef7xaONLoKYc9eKKzRa6
6+wTD4JieRXM2p3abXnTGvLnVCD60FPQO2tZAhaTIFM8c3vYbJtk6qG9hilZzuCLmF7qU3ZQHQ4Y
OwsK/aHcRSd8+uAb5Jm7hIm9EDGclTGFLqwcMdbf+rtRWY4Rl4ujv5DL9KcL+X2I3Om6fDHfGyC+
v2KsYuvwaKvzjWD/6WPs8qaNLLFvvZv3CN9LoJkLemxWcKIkU7UfWvBymaItNhUy85YaERj812EA
jDd4E/NdgaZCvz/iZljJzm2rvhCY54f2VOncngkT+cm88SFLu6b7/lVnddQ9jDgEJzhxkcLrGTE8
5uGbziOe6KCRuR34M8FIIw7t2JtKv4anBvOAhYTlc43RLsECBfI3oFhPwq+LwbbqNHxP4xvEE21l
LjRtidWaLBkiFVVo8IW+ctDtM+WToTS/q3um/hDs5SMi+4udQ86GgC5jfkUXx3pW0os3DbFZD+1c
Viftsz947xbD0UIfGNY0KeAd7NNK1i8NVwECn/hHJ+gxbTIgRTlyuu+mLDhRxttHgwq7mM/aJPRz
hm65UZiTTdvtt9YzGsc73eYP7qF4JqS45TSjgR7VTsKITg1z06cE20o0DIYjgAQyo0iGM1P4jEeI
tQhxgQvWiozpjTqryQf1/Wd9VXXYpithlqgpUjTizIpr0HC7SvqGLDZFk74yDnKpYVjOvg/2Encf
HXxlHk5kH9X8+tO5z7+XQOHnziukfUKDGe2RZETwTWqWOxx8h/7PuJn4k86GotsOQOvnVhayM8aF
SsOfKzhg65VbZV1x/k4n6+OKFtY+D2wUM0So9ubs2T2rsZsNszumcqWivVtmoIchkT5PzlFzdpNk
+muvTrGySbWejakPHH238QZZ16cGho78LU+kx3a5zwlaO2CSz6+jdfWcxtMnmck29QHMj/Xd2OvO
5kTRNnKOThAMdX+/sQxJbTkUBrsxPfCHWYPGV5lsgoL3BVKzlK70a0Tsfwc6w3w9iNQKN17dQFDi
VykxRScq5xICDGcHk2Z0AUSshcM/CDXPrv9N8U6jhT/n6BzYFxrQMFuPVeiSlP9mF8Toh+vTvj9g
hbLkCl9Omp50zJnOaDuc469kM1Uio8pT427W0vpzhumE+dK3vMkReblrlaqowrgOYuc1VOk+vz8R
pQQY41rFOkeZcyoGdfsSWwVZEzq5evJBKcYY8SNdMvC0hP2zWMRt78pIlmcT+i1uRzUwfcXZVtER
h9r4/mUiaKTlgWh6g+PuxE7vYElSSwmDqZb9mjh+K4SAwx/C0h6t/5Ki+vkOtvXNvN0CIXjHLw0U
t3sAwB+DOBHa34YMW8zewsxbbub2Kp6FtFvYTk8yafCR2sy7qqYk3eq8TTLyg79nEIG3fm1gyWIY
W3d/3T9KHGrQCbjKKNzy1gQsxl4kFB0oCCzf7svP3zDhiS8ffnJq1WCzubLEGj+RukgF+JIFPf00
MNSTLSdwOUJCJHmTYH+v5HKIeFy3bhMq65muXOJU0SJXcHS+AcejCt3mp29yJ2pENpFI93A0XAER
cO7XDvbXIhTWAFwV9r8QXKFUKtz/X1Npve8gjAhnJX1yjKbBbuU0rvNLQYnd7mpc1sgNGtO8hyJs
QTVHp+DUrnIhnWdGHWlN1dO3IKvq45P/v44Rfk98EKqBwxzjqs44ou+mLOJ5DNbLt4fzIfEHfjLy
bH9wq61n/9n5oBfssXCSEMzPqz0KGrpB1vt6I11dMT+YpiQwFYG4cKi7B3IPgORcz8VLwQPHqngV
yxStnyWKSzN2wtrATTLUhkw4nVAB/FCg+jcBBLa9CBMm0VOsIYh+uXQ1N77La1h9RpVdYIWFpsdF
ezH+qAwwyFd3avG726KXburLIPraQ9J5xXSvGp44moddC7BdvnH/TE511YV3DMGz5eX3kUEXzryt
uFVC2m3XvOW8lFWZnjCG9JaRnXLTyE8+vMONKsyep0CCBmjlUMMK17XZCAmD4sWfurbPtNUf/UxS
nNps449/T9m99qxA+7d87HKdmtcGGZX5iwY/keQfKPJlMo8JkjlHm7zPsyCUBoUGZvoRClinR9+4
8yLwzDznw+TfleIi2WATteJ70soTiZl1IuGqVZwaRGIJEno4WYmFtUmFqqSnPIrkL4wO7wGWm+i8
dc++S8W1p3/Shm6cIOdwZrSRxcMHX2ZYpCcaDkSGxivamOgsNg33Uu3LMAZvsIgY3FNO0xnL+1CT
9Pf2s7U9UQ0B54Aq49Xs11+e2kcPyzh1sr8WZCkKRjNIBJMmNFxiVP+6NiA8irJEv9uXGOP6g1F+
hFFQ7oUhLqJYo7fMb2yTHnNUZzQp7zQzRi6UgjTHi/LP4ZfvTmqkDk99NdnPKGYazrNUJGjpNU4h
PqHR1MC/vLYhZIZoGq3unBX5RUblqUAkIKLObxNhP4K827VOeg191gbNzHSJYhu5aSuwcJ0VBHSq
x353wgMZFJEA9RDtzjLFURX6mWKhvEmPPo0fadIdQW6nJygPH1EQjVxV9Ou+hlxRpbmd/I5CN6pJ
ugJLRWNW4wMuNCYO7gon2Qs5xbmKz69avTDTMPL+0g4wCDvlVCH1Ca0/R+gDk4kwDYGz75ZCPy0W
Gbkq8YkHJat1T0yP+bp5JoZ98Gs9ucKgMQjX9AGn+vT7af8YipPacvrA8/zg5T5uDSEJlAWia61B
EmHncDpluTBPP2iVOo+4l1fyQhWRDPYQiVAtf+fwY7fkW9Zs4emyLNfjRv/uEuZ6DQir3xxGS2Cu
ftjGOZT6lSCb1+W4B8pfeEjCGBKaymfdqp/OufS1eAnCK0Di2lko49LH/mRy7OFDFo21fy8jPfP1
Oo2SvTu5jbuyQhwCPhibgxdROqB44svTXHwK4qlSWpLHFUHUAjkCIYp++ot8TWWYtfU5KDQBptr9
a4C9peSKzLZh7LzGFL8XGuKR+MpvA6n0b9fuo7pFO2XnLik6t7c11Rpk/DEkPuckdVB3c2XCJRW/
KBY7o1egCuD21gyTyeyScIKV4ADlVmm3BdW0cK51+4ZOgETjflFiz6UEEshSnYcZaAr+aDyK9/Ea
QXv8xD4I7G8wQD4UpgT0Mfl8vsyGusUehYmb4xaAwsTSZWsoCI3TU+v5pguT+Lywq1F6QQURA5iJ
kJekGyNTOVPpoLq5vbBvrXLDNWPfWS9w273ar+X5HcuCnZXK/Ym5L++7iEYk8DcsZssWVHcfUpsl
4qt2IBkz3OKUr9D2/xFpuZQDVaGcBLx8GnHlnwynzWvOs7/o9NnH4+IuAE8l+9w6mgA1hHHj/12n
bU42ZS5KmCa912OXbsHqbyzT2PVosK9eNAhicCmFqJXx6elqXv5l+07EuEh6fQiW0xdTnAYk0hit
uJ8aYC9byMKUCAYVEL5HQg1Vl5VZg3mDrSP41kDC76Ne21cFKJBeFE+CbBmbbw2qmT11wWdKeMEL
/7s4ODGGFc9TQTgfUAZOEkSZLpHmIsH2+JiqQJxjajO53g/XcjI3JxgmG/1u19QSPXHntfPYkCSu
JCM/z3cOEy0M/IT/CPYPdYWvVjxi2PM7/rklfhyYQhOemzIxS/5kwvcC4Xcbi/7u8CKOBJcIFQrM
tg22DGkQlwtTvfQQnOPfN6+2iuNC8CtHdkgLsxzpFy6zLcnG0cy7z0JZDnmeyIY4xjRPtUy192Kk
RLx/z60Sd7e2XWaE9Y3B2AZik7mYcXGKj/obekMukdnfiYkpRmYWHKOgxMRwTpnr+9zu0kzrxVzG
nSA5efXWNiUlU/RwaSCqJBnBug2TdDYBGwUaup6/d123l7jJ0D8FCrLZNEclTFBdmWqGpMU5OlZr
8yJNJv8kQB2LTjtlLs8yQqFt4y7c0ozASYOWu0Ikq9Az7Cc3wsrxAZHmN+Dqo46KA8HtPna0TnHw
NbZfCDiRJ6oUYjkff3+Nt49PjNYN94PHFYtrbEp7wgjz6ZewwnlkeMfV7K71aMg35FTCcfE8kdg8
KooIBOP4v/aZeoh7gBI7LURiybhmuOi0twF62A3amylxLW9jrpHy+G2fDr+qjr/iiUNQxRTourBm
NXnYWur303SkFYNzGPZ+4PtfplYoRMoqQm+uGJMQIsvbxP1DzYlN2YfOT9ZUZadus8tNBt4LsyxK
oReMjPF9OjsgcegJwonnOtL+FJp+sghHqwKq9EEUDPfkhhFwisnfuVxOQhOp/QARSTUi47LahIYl
kaOFVnfsuK9GsuZwX0qHCQ84NIy2zj6n1EscVc44nCTlVHN+fytU1d34uMRd644oGipviu/8XJWb
xU1Hsyf3y06ckTLPivLruutIHN8Cz4HQS4KJeIOQiG1uul6ofUezziwgIB+qRHI7omupGKe1UVfh
vrg3arMOr6dZ9DBsivA2DSDJPYxWoW7+ylC3zABoe4MKp3lq1QGsDplkzNYVoGr1p3iUWvDX+MGa
55yRElAI83wVmHNIy0LWywrKvIxH0nQayiH3gdpbocIjii95nZUehh3BMnefgs55D0Xgc8xcUl9L
6Xt9ZZwNh9TG1FCcBCXlQ4ihWJWsrkM7+4BNopYNSjG8BXwrCAi3OQJVBzziNdgpk92YTvbnAtGx
Qz/85G+K/HhzUn320qtZ/+/VZ8dQUSBgQX+fKDQVx9gyBl1Fdgf0igfmsEK9dU2Y/XcOF85YOnLU
EocCj5pBP7FWhgEie2AhJ4X42OjknSRl6hHmvQ7o8deAEd1Fx7xBIgkXKRcy7b7t/7yQvzoxq+4i
ueazhgSoJpJNu3ZOQo5YLFPHRT7mzY4az8O2HrWax4YAziZjnGYL4VwdXjIWkfDj0BbOf5dPwyX6
67FFTRNPGU15ZD6y5ipZQiJfhph4DuwOI1owA+YSz7NMAfaSniHrEJMp8l1882A1Hd4nAplRYLct
96+Z7MuXdVJX772GEVXCoaKFrOEqaOP89WNEpwcbSNLAV3lPduNpWVAQDc4bR9IVV3A330RHWbYb
ZM+dRcH8kaXV4F+2Rzs2cr2Y2NOzoV54WpAtKIY6uP/WGJqZmzwJvFPw/PgFkc2WmL6y8f+xZR5g
7MoMT5XSU9x8bCW8P65k4dhskbFQOvOB1nlqyUAwKfrcWvLWGEo2FoZH/Q63g3a2xYKdOHJM9QeV
RDj8u0F3+0gMjUCI3qIfo8bpFUuqX1qFRfr4zJJaPB2unm34wLS9QKCNyr/9DHvJRlVgMP4k3FTs
pAtCGSoTJMCl9SzRNVcZm7bpSxMHa7OePG4IUemQei1xy5YG7nuL8anxh7lpNHoDOMh2idPF7iy1
s4AGsrUphjGI7Ljexu9nZX0P/xyp6eYhOmHU4R4ZojzmxuYodkTxgYdHVikEU615pCpmhIZ1H1k3
RST5OtFunU4ARe0HpH/BCIsr/W1hkqcMZ2Oup1QIbnbpDrsb31Wd6Y4eEHz6JRh9+cHfyRhYrZ03
GLWqYU+9VOVRP4tB47mUPeRz1ecUS9gv/E2/VP+NVjEsaA7RR2kDCILPuHhiTedtySKxeNvLeqNQ
ENdxRT7XYNGlViMkq8B/qIJYV9jRSkD6vrGBr2Eny7FGN/KqONTXbaBjff0LrM7yYZG9kHjWzm+i
JEtrfnw3g8jLKVow6clJkH44MKEw77IHCCAUDeQnFjspF8BHgEkGRmQ9i0B2CoYoRcIvwsSB4RtV
4HkXwJ9PCcp61HlGQHWsJMqJTNLxRfZFnGNVKyBF2+oWD+KJafZvQVlULCrskxEEOzJ8ycUXbzeP
Q1qUrT7XN9ZThMUgnttiMt+qh9quXTL3dJg5EOuI9IBKEKvaCr5G5guHFsiBrwqNp42Juy0RBQx/
Zd94Ct4Q4jgFz3LNPMHJ1L/2hFdRUr8DOzwbhueoj53vJNaE+vsqun4plwuX/celeXsi4NF5BUj7
Zwvx3RKX4Hadd9XnqWIigvopkb+yqDwfp9qtfuxR/efJsxUuYzZ+GEAUOd0ry36rxnkfBUaUJ+Y7
9Qq4Oxzf51pjcq22eguOjn1ovbeP4xGZvcEuuGGUL0TRU8y+6LslypcaVY+MvNFikXPKuhfiM3lM
Ft/xkCoKwGfCOaAAoi+XofpoaXNX54ONa+Ufo6LBrll62XoVLv9c87OJgxNMs/yO9p9+TLn5vaxq
uCSgPaNjczkN6THAiF6bnk7Qel4mjgbcflsa+bof7pxCmHM3LUhdYohiym4yGro8p5DtjMLWs27R
sgodJbICiQW7jK4UYGHoFiODV+loK3PBKAahJWFED1jKAiuxbNyKXw6yZqfiTNEagSXXPdrZXWDf
bgiGRh6fnIsOYCPc3ZVtTX7+DEOfDCQaM8PrsLwMA9qU1WBIBCsEtH5O8Y57ZVbhpk5neMiaJ++3
Hc9NUlwBgD/poPrySpz+WinxAh9cM1y1CajzjYDMWlqme+OvBohp6rKjJpd00H8P7d2x0EPKaQjp
knkmk0ySAQsPLpAuwb2bu/DstL6kiKANcLwnLNzqQv0CLxUJJPKAKsN36K/El69BlQLAOL1hEwBm
47T+qjXw6vvxEnEPepwxsZ/EGU6zqaIbb7euC7CCB4YPJWiO5tMNtLFhk9YXfH7kdp1Xu0wr9wuZ
iXxJlC7yFf5KnIWo4fnUxMDPhbPo82K+UnoTjmVvYj9HZwOFDcvE05ihEXCuMroIpVsla5MfvZwi
nLk+6PjcHuZZRC3c0EjtGxRSnRl2RNCaqRCFMnkrkNo41fUmdUHdHLQsPa2xag/F0g5dwfE7dPbf
bfi0kyA86v8dpdpT7nYSjUWcGiHQPQR3x/3P0QaxssJ3Gqdt5J+xclZJaCCYitw8w7MmhOrf+RJ3
Bmxqxw4Y49Kw5zvgSaVbAtqStBCuDP6D6xHvVV6Z/M+ZV7bfIRnG2XGDo2cs/lYhCfcRIIMVhbb8
h1txERLH8zWs6oTDhFevr9HXM32qpH0Al1EDErYiBdnNUb/x+brjEz65W9GpYrAPWu/yAuPNiY6I
O+cYimNwswUUCtJetr0/5/vPXIlXq1yJV3AcoIrlnXGBsOSWPTZ6XE4LdjrZEvoRVBWPxTJ4pCXP
J5SMLBKFZY43xzi/vDzvxR/5DF7pj8dGXoYB5y1Hveh6NLgUzNPf2gX44ep1HKnbSHBKHFI/5USW
A3IKhDENaxlf7wrWXmWAZO0u55aY/S2Uz/lUyGK8hnQAENL7+Kk+9AZ2yi80zUI6jlQBJVzqMhlx
8630beUmtyiw5eBdLA8GawpL3f765pc5CvdVp4YfX+Q6uaAUmSWkMxb8uzPbzbH981IuX9foeAy3
QyzCVpkOtJbVFv8GJVwU30CXK2/s8SoqpDeRaZ8JK3cB2vIql+6zZbwB1UoYAozpf4fU9MyxvheU
YJVK+tsvUepY0C0tiE9b18zmdRmsjHCLceIPNezRZR8kc5yVKm+FM6qudaWlC7QgggWC0GNN2IRA
+kWIAEgjcXGk90vFSZsJh+iQoB4IkAInq22QBW/uHyJh5WLPa9ignCgevqkvkpTfXkpAfPMdFPEe
StI47PSZ/WM+mQmccTGxDOsoZdV4zisQ7LqFBPKVBDwVKZGNO3+CY8s3ISDMKgizx8XugYKxaYsx
4ayD+3WqQoBiQx6HTPxHvLsGRcUww5SyzS26oHaklUBTrl6f9d0T42p5Y975SKBu05rErn12dHC4
WbhYqd8U/XMr6h2GFtecp+5euqnuHhuXFYsGQh8czioPXKLKHGY4uSwrWuvTmX06KALMIUKzjYho
zum7zYtCPYGt3dlvB01HbEsaTsRFoDakI+arafGg7PvIivyCAQhHbt/7EWqPl5/G7YoS/dnY+lZq
wA+1tH/FMFqGubk9E526qVBHPAn3K8YXzA1dB8GJxKyzc8l+QCm2GT2jBdQiGJ9ZNdl/js6tssFz
dHNjOK22RcmPMjCV6SatF5itGDYQ7YgOGQkeXWE0j169zDeZDVs4EjDZslKo0eDjDd+j1bs3QCY+
Q53b/FVGkcOaNv82Lcqat1rWmBpcCr6uOP1VXwuBacr1rBYIj+P+55Apq1AOMgcI3bxUtbmpjMCU
0BkP53uTn1YIK0wqp1+rjt48dYvaAhT77eCYA0OkTwhFepOgdemYOhAHSwe6XBFbr4s0DuDfR4M7
vIcIa0IJxF3ifY5dOBNKZaXBgYFeO16++OEabGYCWA5jZb1isHfRfVn2sZlvQXbCa8LKbRUqj2/q
J/07dnSihlOT3+lf/D4XpXsNYO6fxYTm+27JZvjl5OkqEritWSYrarjf/isQdhyQEZmOUZZZYNft
0+XIA6T+tMG3avHe7tt8DEKuKqoP0RP9wE22uN5mTgBhswS/JtO8T2hHej/IsGPNe4EJjmvck8XV
Pl/2Vok+fur7WoJMnnnJ+IpArNsNsDW+PFtie/KTWmDwSpECPLICsW9voReQhJJgmaqcKYt2Vh9s
3+NzrKw6nDl2cQqf65VpzmJyQkiIBkyhuJHQmSe0ujvn/nQhtRGJaqfvmqdI7810fHNqaVle6Le6
I8uyE4uzPuLIGtW88KRSBTcSd/PzmBLteC1oAurvobiLn3/a3Ry/XV1QxI+LYzej7foXH5NM6JEY
WRLUlyQzasjX3WoHmjUtihJigGItBtfbLWyuW+i9UvVmtIPCqRsQQigxhhd+mrVlei9sWWIG2x++
7ZVlSuoch4ozRaA36nu5NiUWX8GHMNBNn5lTIDnZOTYkzgY1FzSQlPKo8e9aRnLVtrWSvuwQQst0
Chd+EQTXkUd865M6C4g3/ONI+dnHR22u5sCt02xIycHRSbSoULZ+m9+Dj47tlVvEtbOsznJ/bkaj
n5bXDkId6o60jXlFJnM2TEmvH5IBkRcoJ9o6pXYF8p277edKSWDFqzNokwNoLUMFo3ikqhE2mhF3
nRfLBw8O6O/eehA9L7vd1CDY6g9xJXxarkzzcFBGsK22BO29yAb7r+lU+p8DIYyikWiBduvU+a+U
PIDISOsiqONTfF5KNESM6rssbGpCAAneC47E8N1OvMHjSd/Bx1bEbJcpFXREDxYjsnDOjCUmB+XG
9PC2z/2KqQHifQm79KXo1veH8rcHNKtqbuHeUuSCrc1xV8jNwgp+mGziZKtO7dXPcoG7mVP578T3
82pzJJudp6lGvFoKWQ25eVqdI+5U8bOeAug1MqMENkt6/GOAJKjPRiz5eqI/fTKums9ypl0Xbjfn
keBanTEhyNB4EtqPA6owGS7WG0lg8K8BsGQ0MaW3DKgFTDzPLhyOTXiLTlXD9q9nmR9RPKsiZvU7
9lzMjfqZ46Xh/HLF94CFq4a2xKEXtdEi372UVmw804ivTCpvN5gxnjZBi6tQcZx3UcQcCIygmziN
E5JWL75aIrqKJHHCTK0GV8mlpd+ZhR8P/ChhEu1SDG1qzV9Bn0qQMtE8vim28ZGbykzFRcQQ+ymr
617RdEsB06DCwWU/AwraN3ihOBuGE49NdIZmYEvdr1Oym4RL9++MjNJImuDB8ynsGxWE03uDnAK7
cckwJ/pe7lkJTRB4Sy1unXSINpy6njk2DGMOXkmhQsmFMZPNE25m2ONO8zXaaC6EGRabmna8r92t
tAstmxr/Y6GBPsPbAFlRWOwNG5WLGCM19bBfi7fV1TaEa3Pud6VPkfIhhlJdDxlfskMLsBAPKm7L
M1GyEKhpNgS8MgSXwnxD/6/D/agel/93brIIARbflCVEllsqHTzLoqzTvY3q6gWCv0mRTUNAgBRb
Udg91mTrkekbx87bDE7p7icUSVIbJkIYLuQAiFAJoL2juOoJzZWsPGWqth/9qrg7JWAqA1MelZiX
1EJOevRfwFCw8gKxep9aNXIPCbTWI2kY6k/sGjNW5sWg6D6gtuWVtwcvD8YFwvuVT//3plVKYROy
j7xIwfkVLZkuvwRBKDeXDwwedVfde2KQjQwPr8yJTDFKdaNnUPjjqbh6EwIxsW7MThXxP6jDEnII
ypGvcL/qguvLZVG5ROeOibuZDw1I3XaS6jodEi6bzA3Fft+5TVldzvfK+G/EEJNrs+ozNyjZl2DV
CS6dJYbAU+wgOMbMPcORd33OVZ6m5MnKxIds/RXOqeJStfSV3ACdtu2DV2dObMd8Scp1CK6DIGPY
j6LKwAnnHpU2VGQtq0ZAcHTcylTFIe4b+O6EgJTEx3ywgelK64aaION9ow9VcDioFGSJIwgsxzbA
buXsjurSES6gqYFeysczxVimsg2Jk+nomqU7e4fgtvTeqkNxwkws/PzU2vzGk3Oy0NsVeIEVvxqb
8xbXy7es+abp+E9SK+bsoqUzOkQjW9HLBrBVrVIOikHeYnhiQDghH+sGcyPGxHz5mcbqEMpGQPZI
RdfsXRmYvxv44J92xy11cBLhx0UmlYpIrxK1WJWcekqo8P2CFlJnkM1dtvfBaN3NQzjMzAiCV3rm
Ql2NxdzyEPOQT4TwEMA5Pz/D9vwExQ96CuGTZJxkwCEObIos4Mknl0QMaAdGAGnxwGRMBUdoQcqw
zsMkMZ/ImFwx4zL/BQfldQGsXjx8jHIc/V629jbflhoDaREsU8L7Vldai7cJRA+wXHr5gQKhOvVk
60mQaPqMUyy7fNTdKiWmuVM55fY1UQEp+T0ce3PGfXDlsEQ7w/mBY12p55oNr7uLED+stXdyb9U4
zFvdPrWx9FUAnvF9aCL6qRsPpPpP2MfTw641pgPvVKQBQ41/3z5EQtZRbQC8kY4YHU/T99zkpM+Z
3IVzEYOZBUTv49MU0O03nQn9Ex/rEQ+/BboJfYGX2uYizhyDFMRY7HPTVpjcy7FeN7Hx3V/VafTa
qJmL3VXJLz82DraIXHi4WTjbjeoxXs3+ahfR/4IkTyZHKeVsTxI0Nw8eKzo1uupWPKuftcI9ZmXd
lOiuLAoBcF4wUao/jUGerFINxickEaPs/00bib2tmPJ1b7+RK3kfAryDIGss4vWA6NJ3hdU1wDoI
RX7C9EGT3oOY7E0VilBlPJxt9TiNFVSeSmCQW3g74fU2Z6V5zshKuTh0bowNFy0dubV/CR2QQGr4
GQ9CkHplxaoHw4thVs4Je9MkhmmAhZOednaVIO/F6+Tzskywad5eXisQptv+FT5Xz7as2iT5YWoD
7US6l5phZDLO3uMjaCcD/L0wffzbPYGU9vodXL14LZOZwzpVTjfs57cl+CtNrjJraRPtiT4cxzhW
Uh8gOCYCEdx4Ue0+qFG+tTToNnHMFjfbFgXzEdego/kumKZRx8M+rpZBzw2VX+N8jkumFsAVpwax
P+WCx6o+5FW0abWa9Fdc5xYleEtxqT3z+y4VsN5xYqbe4VS3VvlOQWxJtQLH5mc34nwlB1OZtHqq
nyRlXQK9bYeC5daJDcWWikzDnh8B7NiHes8H889Wk/T668c9ZYrSU9oz9w7XGwsg/EZ+hpCma5W1
OckMBk7CGZ1a3v/BPRemxwmRZ1mx1KEo6oGd0YsqRlTxY6Nj/GKaKutXOkymoQkXIjOB0gisaf+0
PDLB2FTKEb0UaSguX87qmCSIh3JU3YSZnYxLq+444j0bKVeEmSNcFwA5n8oczb1rTFEaT/HQUYw5
GQSq9VwPqxA6dR1ubCrRXgOBsKKVwBeaToA7nulfKICZqFsT4K/cteJbg5VGcNhtfsoW9GELhPoJ
bt3o4Dk5t+eodh+RVEmFep+FWeiNcEVwyJwsx8GOAeWjx2iSMdXoaUeJUJkl8tKaLl1ChbBvZFl1
HEoX8jQVpkPBoFXIw7QJ/o/TpS2pBExlyh43vHz8ov2eYkAURh4mis8AdYRXeqXlSdXdFn5okWxe
uzj73ox17TbNWgbkPwiFSSRmbVN+k9EhGFSNxkHDcx5BCGMcnSUVmizaVicP0XKDdKysga86Z2Py
AQrZ7TGfV/Z85pyBqjuM+IofyF9ZlUjCit8oggH7WdMmpvCNcoPi+3csdx7Yfomr5HvLblbrIVVH
P4rRzkoXsWOlm1odmmmDHmMETUL56E2ApQ0nwz/ZYWTEwlIY54Vg1LRUJ00S3Oe9FAKgtmERygvn
JgIk2rTS8EqwMjuBZbCcQ4++FMCtuPQKgGrx1wESVrERBzScdSDf4TGNhLglX9ju7DmyoS1dwQdb
aC8IH6XebWm8I2fXKIdg9/9+XkY11QK6XsyXlvAQI38mmcewFzPRhMKkypWxur6YKtvIujlH0bcu
Nl1U5BnDk2sWmvS8N5xuZYkW1EF0YiaH+giIIOPWfTCf7m8fou0oZe9jczYKbWbYSRWFZWJw0a6n
XIF/mzC/u+vs/6TbtDLKSZvNO1UHFmPwMeF38kBv3W/NJnvnc4AfzfACGgRSDr6lBCwsX53ZjnLa
jdzWL+ZGLq7TkNeir/gSSVqJlT73xBxif5St7WIdy0XOn+QqoVI58zguEv+EnIsaj6UYphBU3H4M
bJl9meUbz7E7QtSyVv3wgZ2XFfXoav+AoNsWQsHmomptKqm2sMEP/QYsrHGH0tSuNf4ayFIICEo2
MdKXh57PN0lX+UtHpFo1Q+FmP8qdXGoRtq0Nfs3twPciH/b3lsAyVlej4sSRQfC0B+mlsCPgeIg7
yfgHnUnnHKcltGHfxipPZaWa72LqSvplblePuaUpGeZi9WBVGiXdw8YBfz9ODTD30VUftL3RkOBh
E/GMOTmHPMuSXRW4IIXdA2YtRxPLWtErTQFQ/523584bMz7HaxuTYWwoC1IEu+Ix+J/tqvDco1wm
oxZD4RMwT0mpff70ksUYUqkW5jYWPFi1yuOJeCaXSWqS95yZaaGQgtxyZAMR0Cs5RnNZRwnAhXK9
2xkPQFKbfxlrfGBx968zclTD5/k9O9vbzzFHhTPtLXzf0frqSULA5IXQOQkPcfO/lDBgSGBLFFq3
l+R80OyOLb9q9C2W5WE7+H96DON/dBIEchPIaIJei3aK4fzm7LgyhI+V8DMV0wopTc7R9NQ/yF6j
38jMIYDaYqRCF++khQZcCHJlICWdGSoj4/Q7Uk2PGE+Lb23Xc2bJO874C8Y3wCoOkKeatTrOuXsu
Vj3CLHoTw9S/d8WxpCx2V23x3OiWuNuFf0tOLOCTPO60rR77zZPomAJinteMVZ34kGQ4cCP5tWAh
/yskMg4LbfneDgeoJhsqIr7aYS9eD7P7MoWMmmcaTVnMyZr2jCD9hJ6Q3HpGmmxMizIHFf23bvDV
Ny6Ps08D5R8ofCKqDlaVJgQm4tBJY+VaZDx5c0lvSgQFS5FDAYCzQ5VOARbDTUazr+Pf5sjz4ynI
sAa2GgW6lZPozxyO5l+ZE2pKbdUOdWHwocakzUOtYPuVxmmlwW1+Ga78fm0pUPpSaVugPJcuOnLK
pveASrEo6cYBcL1jbVx6bHGK3p+OykMI3ko6Rh+2XofR76p8ChCCX1qCWKsw0SoC5n76ojazdrx6
zOalhACL32XSTt73mroi37IFEH15tR2KWHKbMMv1+q5SSOBnk2kR+uIM5sINaWkzC5I1mrVHBfbZ
caTgF2WsC20Mt/SzEmYVLvIRM4LeqXr4at6andABscI5Gpu9u0WjQzFSbpOy1rAGTeg0uXbr5DoL
e8SzhctF7FY5fNfOGsWGDYD9LYF1NvSkKSSZLHn6piPn+LUodJdvs7JiAMwptBcOM7OdqSNwmlOs
1iHj3A1j25A39DDHM9ukjP9rTEsmT+zyl+IB3gKPX8z1In4bLHXKwP+Rq3XaZ37Gb7jZXHxSYgQL
AsMn3RCqe7ajTRpIA+bheO/TvXDS82QXxDRT92HJqhA4SWT2mlHnFsRjc9itfyuHbdGGR/RwD7kG
PKgVzkhbNBA6DycYWt9ZoHn06pmcpwk9E2y+FaRoZrNDp+RWI/E5ltGeMdCejUGnXVcuDNqNQaZo
ESxSg1vwpXsCpvY9dizY9d1UTk++kytuU2WA910qSseoCLtDBl+s2i5qKPmICgbI5qjEbYmJjqmx
pXltm/lxAj4tb9YCAunZzXaMHPOXAY+Oy2j+ZyFQexL8r3fRPs4uwLmc5ElZ7Lt2tOtTOs5AmCAS
1SFiiVMh9oqH6j/j8BRg0fxOHvaIWhXPLZ4vEBw3rMeubOg4/bxZzwhsRYBSsenyRezQfytfE3BO
3AZn/18bg3I1XoluOkv+4zUD9SodOeJjiWeFkInlNNob9/GFEjiLzR8U9e4fw1BZLkaeID+8iIn1
lbobgQS2L0690o9fbXhi+lP56q5hfkfoZVU6DRjha4KflXYVDrOPo+Q9f0kMn/o2+CE+lUU1WpAU
yt1nMvFRkleFnzKNYq/xOZHkL5xfsn0u5LdnNMVUK4TuXVtUlbHXIT9JeqfcKsUjwaLxdqULwGgr
w8YVfrTLS92SnWVnuWjPltHuZWh+ntTVV9PjY61vTdclrNSyFaag2VT73WzTBzxpedu3lPLcZgPB
v//cXzaDQ/cAHMoIvefUcDpUVY55FX+Uv2hsIWbAACM7A/7LnYFXxajmyZ/PRf+55hyHcw+j50AI
81bTuJpg+e9pDcyXTPiGnVHtI5jznTh45DyWS0wx7XKyrXAhtnfn1m32ohz8DmZLCTEjns2/CLAv
V1wTzRIvNkOmqN6Meh7Lqx6mUGuH/7p0E14oxNAxyqVKn+SckLvNa+46guBkpwIuY7ykw8EGtK8s
YeZzzujo4JhPsUhT9ZPU/SPkUjnpPGDMcO3de5fy6klRsBXmq+LhxGiGqBRmci6hmVTq4F5Lw7G7
/2Gq2gw/NzztYN8cXRcZKZvtEpKMn8IXZfGTCTHIMSsyOE0G3Z91iYdRQpO6+lOSNeI3Ln1eQGyC
iCWMRP+E0BhN+xE8DyhXh3apOAE6bsqOkEgfEu1z7zqjqeiqWKqJXKfQA5NVsZyfmC8Zg7AL0OKq
NQGnU4JKcPUBtBj37wUScxPN9LFl91IHg6lC2/6YW9MOixH7+R0zf8DKGhoC60y4qTkQlBQM1Fb8
EJV47WzGsvTFxSpUMxpdAgv/aNQQ9yNVOBk7wL4sIkOsGJ8zh6O5RvuTp3CeUcBHncIrwWpF0iaI
eEhqIsLo7lmbdSE3aLfr4d3wAcJblO+KkFj8PCOhT+RCcAht/xcDL54Ya/SNensdENcQR4jEP/HJ
5eQ1V/goFbvqz0R/Fgr+ANE7hkv2tn54vxsP2FXrw47QNRkvcjiM9I3dgvAoLyd9E2mcjeCWVbiH
cpezHU4AhyZedrXxUY3vQc8kpdwgXZV5eioX3iGFg/gCONiO0SfTu6jDqfuGXlw8XnwBC9ruCU79
QaDUEgNm5X4v7RkhgW6eGgbcOqNSV2pEz9pLFiFIoKbQEHP8BxsFZ5eoc0rhZy+cUZfHUl5gVu51
UEgMb/uly1u3eVT9tXF4hHSRodkHMPyUY++R0kleuihL0S8u122kMa3QyunYz3BSBcPhJPet6TCJ
r7L+GZ4McTisFmOtRjQ7BFPBBt5Lgw5lDDOeBr1kEInS2iC0T0s9g5LH7KdQb4nztYHVhW0XtOl8
1iDia6zCHBpElFqMNsfUMmW4xpd4LGKmpCfUhb43fOY+v99XR+L1czCjsaSPQL+FfAFGJ8h92sFl
aHsHGwRUCT3sYL2PcPpxteBmoHvuagMj1fJ6zi9wKTaLQWKU97RouRlG5NS5xluS7kMPwjSkbiLz
i1pZFs9epf5VBFYSgINqaX+zoDhUjxA81kXE/ccuJkwEBHr0yjFj7cKeiGFYtpPMXuBOZf+gZYaP
7vPgSNNH4lilyAXxdvlsnIUgFFlFCBCanlvu5/Nv7mynZ+oAYoE7pixqylSv1p4L3Nsarrgdz1RM
7uar7LhPP7TJ8Qr2Upu80RD42lJVrmou9iFyjuxZjZNz5OHNX/070g2+bZo2lY/frmM5wsr/u2zp
AhwVKRR/2wuzkGEG65lkrDJiDUzNsxbEvamSiBtbvnwLTF4hqvzqI8HDpX7FBKBVPcFaWKqsVJbG
Hkw6CJuiuhedqAlpMWFD+Nv68GG/7EypCVb4LV+IJzucXJoW70GKWseHdvqUhS4mYv7Q2t7uR89M
ztumBiqkBGo7cI8fTp4AFqxlJGYFI/ZSAHj8NDPO/q++R/0+3OaNMEouSZf0pPCjyzC56tydRjWD
B7E/fjmmDXDLhJNyV0NLPhAKceglKzuek93KRcR51GJwOshYLmjdEnhReGQkSc2WHpkL+d0bSki6
jB1xsruzvFYuXxNQVb8FDEZ7/R8Gh+lL8jGI3kVdMynI9RDoc0r9H33M4992GJ9bAHgNjwk7vd6F
W5uDcuRSRdOZDLxFUdzrc3xjoJYhEnaIOJKcbS0eV5txTWEnxwp4w1naa9pKFcqHmiUXRWh+BN0C
POj6GqpIv+bGzKb8j4oCAIRuWGpIM3722NyrH46RnXBg/eM9gdj5vhHLcLMhsDck6UoF6JYoURSO
nw0afTWHBkvh+38PY3hgEjrPmBYyPH23QI2BgwMjpUOSO5xi4FBvnq/toOkU3ERq4UTtR8/tfjp7
A7m8sYZZ9ue8u7Hamg6MnyqB7OWdlpec4ZkkUhk7wEVGI6qiAfgLATPpC6RxDeAIEiCZZKqhgaBM
nl/lmUvYQ+bnU/RCeDFPe1wMKef4vBTWOOKrOAa3BeGLRdite2PYQgeX0X5xcJnNwc2juzt1d4nh
26+I28ZR61zbjK0HqzfJQACYd5lHyVvmLyQ0LU0KOnmqs6DpnpnsRGPL8mNNhxrVOVU0tsYZPbgV
Mq3FZGF+d933fIlKqRTt0bQHAZt2nQayFkQmBmC7pjHP076PJSEYhpnBPf+kKf6jyApdt91MwsRd
qOBM+mOeqgmdeXlW0k2h2awEV1WmEHTyNOjh5GPePEgnqizBNuWYvyF+1jhJv+NXRrQOYi00DZbs
cVZPd4ysMvyREDt6v65rseaqrWu88Zx88Xe76YTL6MkJ0yvzbSveZ/HFttwKHdSrTj0DYntyGgvJ
eEdiFI1ZtAX7wvGzI38tUH8P7sL9llVvsjo+52Cxux0V/IGdrQ90U2dtypmxD1f7nxszUXS0e9aa
jSDf/DpwQ4QRaGtJIQI9b702nYuDfiK+KGl2gg2NA8N97r80gfyM5qpFSK443BI02SvdCYrl74f6
avIuLmUl8V6cJMIf6u1igxGL1IuTzlQOWNWFs4L9fHQ0FGUEUOtVEXMSjVHP17jCbPsbrqlGKMVw
RqjnCn2m1IMiIov/V60rTzHb0leT7/wQJTh/KSwlecfQHTDNH47JMsWSws6dz2qm1kDAnw7P/0CS
rGSOxl49LovKvy9WEdQVnDScHV4qjYdDRZys3lJcHcksr0Mm/ENzQ/sC1PBUfah2DLDEfHMGAnVb
PgIXHagkQGvWyKQAAdQJ/3ijOAARD9BDgMCeK+8U15HZVE6tH+9pTZmREPl2SzW6+fTEk44TLMdA
3SFPKUzkFG89eyH9eA4Ru+a9M46Ut+dEGWAyYnu6DMAEUIByVCf26+DECllRmx4jlLqxGa7YVYWt
b+bk0mmLKYnN7/BsRyfh9WhX6jbJbW/Oau9u3fthS6gn/xXcQ05iq08L8wS3Wu+zyaWLHgml4kaT
svApNRPk5ES3l12roYmbfcrsy+QjuNTjyErxpjcsBpuPzuJZO728f461TSqtktY8sw5N6/zwBZtg
vvhJMcN+hBao4haZqZ4qqHHwXGkN+kpmUKnRfU9FBrSL5w7gjAcwqJI5CXLUatCCkYhiejm1zTDm
5uc6Bik0HiOd2Eg4GxnlsOHdGt415sgBGFqPHLJsryhvZCpuLOdsasGhQKUJpZz2sKElSrlbi2Pq
nIkfvA1lhNHFA2SsNBehDiJfsHRRCELNfWPT8VaqsgRBP+nYGD8PeneLz5QJvrZNQWxADS1NpqNf
wSTJO50PyOFrbJFENstVLFvmjtDZcxz53Hvnv0ubC8o+nAek81dwhATCYqzSU84IyAkJZZ+mpw1n
mkEiGR3plUxbNXCNTBrgczoTk43vKvkMJ5YTJXK4mHNBfECejY828nZHjGt2IWcHbOlA910lN1HN
VOUccKX8CrsAECgGQQmCDUNdvzRPLejoS2g6xjuvs45VUCagKzhbim9CHgbgV7cuGbOckKqfP/1N
R8/avSMhtioIVN5tXsDyFgpvyCklGtKp8x0HhdUGCt1wahIk9frOHJY5QQNsOZD1Ax93mq5fBICn
11x32cAGMGuis80yWbyVnxgOkD6x09cgYQtL2ABNH73r/JZj/H/+DXhfsV6sH27tf6d1D7hFeanM
i+CwQ23lo1F86+D7RBwRd+vTDD6PHA/ylx90B7lW/PDB5MjYNR709pH/T3mUVBXF97bb11YHpL00
lISKPJc1VSax9BmSZj0iNbI7MPb4y2k6j5XUlD7ZKAwbtFyJXfjQVia5/N/Hx5nOGMYgmDB8GsRO
NoCKt0ohqet+LkN3Lqqp3YJH4Ch7xG7C8KIlCQ3d84BFOhSWAzUVKzQqF5emXrjXTDRPvBqGIoi5
M9nmamkKLoFRUM/Pr+gwojuYlhUnDoj4ZK0KYlZBna3EiwM76g6rxD0yNGaJFmMIvx3gLK+MGTJF
qW6tejk7Vtn+kZb+BmR++1r5jqsX67xenrHP3NaiCp6faWOXhHDS8JC+HjvubgNUNdAx5YG+14OX
jPRBnbY5XpRdjSslRVJq42TZLIvB8Wp9PJMapbMBUDlHA+1gnhcNacyawtyqPbc6fASvT1cZxJ0w
DfXaiXxzAWnuCM9O1ITMDSp4XVK8BREKWgd+YFQUR29OmgCYHqmdCxBKGSVuUltjMwxZuaRWWUeH
QczR+zlbidU89n4Xkta5ER034LWF5dXc1cDyrdqZgh1hlNexe0YHHXT+PsSGuiO1ed+7yny7SnNU
Atmj9e5nk6mgof3iZOkX0bQbLwvqLvhbphCX5voJLKnJvyKd7LR/lXgl35tfb5ndsneFlEjmil9M
jlz8XJ1SZ6vSumuplQaycA0d0leq6T8aQsWSmK3idbOI8YoTp2ZMYumDpnsVDiiykZ3sMn6pT8x/
mZMb20MjddstRfW6QH2QIjKd1QRSbPhP8UzufUZ4TLgmudOC02AYAYZSt2ITOt4rkY71E9DCBDtY
qaYxmPAxjdv0ydjGRsVX/4At7CNiaXtXkPvMkiVIhHnpfDlQcT/nE0hfAV+WIaBI8OTAUIoHUdEo
WSpa6fwHHELhF6ErTJeWu8sX+qw5YErGpmdM7MGRIAmwyJqlblRcVt16IwItW24TLEayDorJ+1PR
5xudrPpQpK5luJntFyz8ccynZ1t3iyxg81hximVWgb3D7BNUYwEPWVWxH6Urrftl0sRRfRUtnowd
+OP8OkSFvNr8ZrSxOenVAXtF0vvExfOf8+uX61fZa/oS2d7yS9rkiicXHkP3oTc1JiXVBPkUFdLd
H3zjgbJuy2ZR8NYn7KZtToWQkBO2aa78OzdTcuqkQB2Fe0XLHllUsZrJ5m8WvJ8ROEDB2qmmmEI6
g/BVlM7fQg6a9oeZyfp/S9SKaOIlqUk4yQ9NQRQWHfsAndPKBQtd5CTaXTlp0cXursuptPeEV97j
ToIjy39+pTSNJSTir81z/KXlXY2llOaG3P5jN2kz/haguHsgDX3R04Am4IvXo1jgD9SyRDlKzkVC
P6heeeh6Ps0YbpCVSFWRLD7AWMW9ZSwMfoTPoAVnsxk8NwGmfRXSKExPFtJ/jwy8Ax1FuPSGa8uF
nkj8mMyix4i5Mo7OQrM6bNtjpqpuGM5b4fOOYUC5wsr/LzPeEBYzrU0ORWfGcTjCjy+kss0HQTKh
LA7Yr3kUNc6W5YBI/TJ6MKLhY/TZ3CPkVnmkFq9MJqmczjpE0guow/YlaTYxqpWMB/OrvbK4DnZ9
QUWuWngWNRTbN3Sjav23tCYSPJA+hEMpdrkby2ZR0031b2OSW+6GukxOBYD8LuNSqT59iugWdw7b
le5MhpiKJqp3ctnyhdIOBFcggt+8vOjQpBEMjFYwBinF8w5VPIvZ8pyomDEhG9eOn8TnD9pgSnBP
t7csaHITMSFFLJ2PO47nVvhLSca7QZwHSqIxGMGSeh/a1UbkQpgDp96R4Q+s3fJzDAbNOTGrh0KZ
Za0rVYrUNazBACVKKDqulZOlRZCTdd6hfwRP5FsGbhazeI24Kawm0N06GL+i/Iz7c3WwoqxD2HIl
8UJYlUepFvuB7ewxopR8xSfDAFEfIiNQJRI9G7FYGdn265wduRTr6Cq4JR1sitv7Mltcslqbsng2
KYNIWAhbb6Pw5RQ0zIf4TwMLLXZQYiBORSYFADd5mKRnPyaKhf+V3+BPWNAx/HW1khxB3K51AzXY
ZqBgluiDhZujNDVGuN0fBotIGxzMn09+jY2nA/YFGVN7RimbUsRwuqh+9YbWHLOI8otjRBY1DayZ
g29YE6GDy+m9LHTWAUY9rhXjp/liuOT7F+soE4t6OxSpw+ejA6C19XAR95KxxdWAn5lakZV7ahlc
fwB4/IeiMPiELCsNbE2hGkgRsPbf6v4s+OOJSfo2ezWGvlXc2qwToLQcIXctK11nzSSVpspT6ME6
oLYdUHEI5idlTaKh2aULX7eac4pmb0nntlZu8maKLFxpaU7sW9sGTx4eJ0f+kctDzHqd1hLN6N4k
DTBxkIYiSoN/RhHvlPhOXVHmM6Q9s6mGlBF97ymbz+LOPCL6tbg7GERlfz50P7IIkyTRFDFD2c9U
q2ykNyyLhb+w9CSwQkimMmOk9S2msfULj4amqGxc/J1NF9YpOZOPrLsbXUbu23rYjNxL757j7it/
BmSIBVRftjFyk7uFSlurX7a+yt+j/97XCBNfAblzvbN+L9fe2lB5G12M0qIDnoV1mtdvXCdGJ63R
oF49dS8p0MUplu0A7Q2svvfL28WZBGiDYL5hLvEVcU+o2BWL6iIKEc09p6JQYg96/I3cpbnSSQ9U
PxvtZLf6AuNP4y7peRrNsTFnOVwUNQr/Jis2goQzg0XPFnQESA1J71otN9mcs3Fv2hrpc+auWhBT
9FCUiccLQWCvuTi+S1NhEVFsoOK2UxdQJsRZgxFXfA/IiChG4SDEuhkkRWsGIjGv2Q4mCyAv6YrV
CRd4mfrDbWGZvpLSgCeWIyDSL5h6Cw1a1h9aW1+B7AaI3d8tfGr6KJSyXI4plEj6jmgpgaL8n7c9
kcBu7+p70WGNCw3N+ObdCWc6UiWeeqMgYzP6yoi5woLdg2X7936sZer4zS6pYK98F1VLFKz1+ZBM
YlJ5JvFCA8Z8KzmPZSShjoK7zV2LxeVdRougGKgUwz/8qSrqBIOHEMozv5crdBrcwK7KC4p7f06f
zqBLNmgyxndI8zo8QB+pEICW6huOxiEfdCW1sk3Nvctp6mMR+fYCq/y1n/X476/9W0p0kN9bUnng
LQrnnMyNyNBxOKi7AG3paYepulWf2DS3hwQMBys6OvZxcdS7eOUrxg2/zgWwzeIinDszqYmii5oh
IeDipDInDt+iHEyjBpHqKNXq4mg4C9cAFol2Tu07ggpyOkhLVS6IARF1HQ1bhZgHMcG514Bd7OA/
9wMn3UqXqnJPuRuGea4UI+1yZW1QH0yU+TQdS1JVq+ANbUH+mfxMvdNu0YLwhbbvr1yZamQjVkQG
sEqEtC+WXKY+UR1hQWNskn1k3pDEjy1XnUJyxmA0JP+LLsPpoICkJFY+o6bwcPL/l3tGBlMFe6+o
XVuqZ4KJoDwuw2isS23+FC07yseSRIoByXbnI7PuAFXcCX5kHmR+88eH32z5oCpz4QJq9OFfCSVG
sYOe5aQMGHhMbEwyctQWOw2LPGD3I54WFMBv6Lt7cx21WXY/3H3DiAlswsJ+KT+Uk+NQFlHa0FTK
OZzIk2yGsyzfJdgltluZf1Gjh8Mw0slxAVq/Qd5kCNpIsaKAQwqk4fX6+WLcxrT7h/K6Nd6AgT9M
VxXFuh8AFJtA023WYXwRwMGtZnzYgc2NNzEwOJJTu1donaT0xChldaq2QSVmm1n1n0hz8lLraYgG
Wo5T5+eBrZraZzuUXAW7DR3jMUHuMH+5SU5pmiE7rtWknDmBoDZ5eddwS6yxM1B3GH24dNczJY7Q
xsDlBAJ3HC31g6of6lc8TsT7AjnLO9XdoKIz0aBlGW3BtEtt6M4K4F0QzJLadhJw0oSA9zZoitJz
wC+G3jBsF3HslLF65rDijmdpgUqFP3zaWIfDTr89/5xjPHRekDPy0Gk73BqKhaLuaUrKzGKb2Ive
uIX8BZvEr+aRkYfiw+nnXJIbsDO+q1X4RkrKfMbqR5oJtL/eES4VztvCUGqq7LSNcUwjRYDZwG9B
/3S6y1i3omkVlOFWu5vPMTwJcRBNiSXyzoaQ4VYUlJKoMtJCJhYhQnsMbi77pLSzpH8bEBGmquwe
RdfTWSF/g8nFNmEFFeQaoRI0WIoNW8XzEwld9qHYUKvPZi2+aZ4MZoikmTHvWFrqhlM7qKV+aMXO
h/rWrG2zOGDXHvbSJ0R9C+wHEhC4XIQrE8Kp1gjSek+lDHCebhU+AItAdOiDTM7pNfImiAWbSusO
PRyzrRHN5WHHj/HOnH8pev4Wux+xcuGhKmFq8kN++vd2cD1t2UdZBC6Nziu5KYKQDqblgCxHxuPG
JpHRaXNFTWbpjNDJmSYBM4ruPxVaZWhPF3JXRhM3KoBCjs3dvuZAu5QdYZ075TQB+YPXW/bsuZtH
cRcDNy6VzZ7ayuH+WpDYzKIcowrEYgWvrLljEetkSglUYuB8BENBoAKJzYjHCA8P2x85Z1NsiZW+
b/Kp4b07gLgYxb9gSFyMw6/CC8Otbu/qzbiZfZ5Ot12odkSPa4Fsvx8Cs/QP9qFBpYiGoAcrSUqJ
ESPKonrSsrrRiVjbOYlrC3zUG9AwnNIPVf4MfwP0/FlCBPSRLVDtoOfjdQbtnDQNP5/5isDnSL8Y
8WtzewlEDT1i7UxCXGpwrLJ4pPiiy9NOkLCeROqk8CJRr1vVjkbmsH2K3n1/B7dboYWuhigZOtdo
JWC/psLAubQxPranX+kd4iUk+zO2ngDRe+4hRCXjzclDHJen3YJQDPT3foIQM31khhb70DDJUTFm
KzEDXKuKJ0N4oU2/VgQzrMObN8xzfrRQ3z7TsnIZo+mVFnVcLU0hl7dh14E6BeMtPb/BefWqV5mM
o+hw8uJEjex7XhCMVMoaRk7HWiCfKAVXliHimrpWegb1/dH3IU+AOguRMWaaI9m8xDTFpOn/SbWE
UDSq1XBZt5x1yTb5VKl220wBfBFIXXyZbTSA0FDSWVnlPOllH/E/kOLalRYMy7wvC+R2811Q6wfD
JFfBZDoAytsip/C58Owd74+LyvXOvDCHpWvp8OwOG4hqROlL+NskdQje8hk0z+b2JjwV+m6CrkPz
upfuYI/qYccaG16MIGlqeaU8NV6GxDc2FtaP50euEX2KR+aF7MJdP5o9rlyi0I3RleHOlPxzSEaf
k72ANlP/E+avz8NWRKFq0qutt8vKfSoBndFBvC+dhmCLXLKDyxSt0379i038J5CmLjA3UCKluodh
YVEMYnebnE+tVgOJh8PI6GWXyHpV8MCI5M8zB5Wxu/SunIloZU6mGJAlBfWedlpY+igB7nIXsEVm
9+ag+f+9hSDyKNzjAc91s06sgpTFbK+ELgesKDgrDRCj3PA2775eC0iXchpGUzCLHp0mgJ/sgWqY
pVB9QThPjcQbfkBn60qJ4/vZdM+0iqy7HoHkeq5M85NTFtmJUV0F5YRkCLKqHDA0lPNLux278v0r
8wg0QtV+e/8h0ppcUHo/Q5jgzhmtC5Fcfrts0G2fk2rQJkkiYVSLrkgSh8SFz7IwHBDh3epYftkN
pkBFjwYx3X6djW5aX606TVhsNjEA6kHe0NM9OUiZBHgTMkt5hiPZxnO1YOqhIlPvBkeashMMGtBZ
ogEXoLdI1SznPxMiyKXTfbJqPFOF84Q4ohpzx8JbmG5mV59/tZHg9uVu8FvaonwR9AGLL5afne4d
1CxSIG79izxtIoVcxmJlTmR4LO9yMZfp0aT0wVwS6cijsw0yUiZlcXQg/xfQGexzSFdeh+JDR0bv
nHDyNZkYPZ4P44DA5I89qcZd5KN+TuEn+ElJ4m0TMJ1l5Z9+jhQBZoUecBTEDkTox4cfs5EMxUx7
07CuF0uLXdukHy9naLaWQJp/fgEpay3y7rR+JTMCMSYiW2wnUUnwykUikO/v2f5BQVBwhaVz6/3E
CG8UV1JVuQvUdCfEoyqdH1h3M/bEABJbpS0iZoHJ/vd5uSHrPYvxCSzAYy0iNTfGqrHx5g6B6R8p
5mJbvl3rlYlJhs3rwPNGitCSlhuLQm5BVW+c/vUk82I3aGbYE5rxbcGhr8264/K63hbfRChcGEk9
dxn9oATnh59utDsz3lQjYFO0ass9AeD/K5zqyyRH42P0F1w6foDS8JmCQEhq0xbV5c1gmVwJ971t
ltVhxUYLJZ9yF+m3PYPTe0SYF1Pao9//Os8BFe5WFpFy+SjL/rhjdy0JjI1C/cF8xxPsv/jBW26G
kKZuufqmpIvuxv9Xku9qNil2Sj694wh3e5i2LLhSErxJrYaNBnrAOCZAX0rphduA5NBh0T+2aiCi
Uts3NcvBYoTUp7OGKX5XilsoWlu4Qkriw3OM8k+muzI3LUUqbRE63fnRtLE5C9KTU10Vy+UFzk7o
NAbYH4imD+kBpb62RywNSGsSm3KgtCkejKbpAVgfDDChOVFnxiXO6QUyK7Fd5t7vdcOZ5OA+Mfjn
DFpArQpMcZq/Ou/kIU9ZXsuMZkvHbp+3G83cAoRu7iAD++v7bcTbt99dheAkc9rbLryFtCZ8nGqi
/wmjVDNBiPQgyoS1sHZLuKzMvgJ1SvgJvQDeGlMOtDAiMMh7ZYmVwiyEGI+vMxOlpDDF4Z+BAqSO
oar7WZ2GkJyKTVG6LKkwxqpi9C55FTH/TsvVwh52oMEW2dSWu/nnw50gkYrIhY7WvWe9y6v63ox6
WMyk8lmw8Geab7eDUDIXHKvQPWOyin6lt5miJd39DIJNb5ZZKD9tT0h3V4q5MqKmyMsyy4uys+T2
jsZZ0H2m3/6TvpBkqDhGzx82c5sjrMEjW6q+C4MA0FzrwVyNd38MNzkP/OR5caRKHIZEczaByMJ8
k2lh2LJMLsZgm65oqFW+SKxP7KOqANTFWG1JMkfty5qGZw08IRlCgjO8I5WDpMEegKnHB50H2uTW
YzoJNNZQ80mfymWsCrOXDP2lJCcsYjSzrOpmMCIpZ5/2xXkVgBh0D0+DyIeEvItmwVZePINxQe/R
UJV5sL6pEwWLrcZ90BezXLuwIh7pz+7h058EQr4/7emmHT7bb3WEijHxJmUDnjqceixhFmaXPWxg
A26amacrw6AP5eakrwTdmfaYXhudPLGiNapZFeeSzC8SzejVHUiEocPEVWzo87J8qr0pejTZPjo2
/aerMuThHILyUSVzZpis0gGvMrMwXXpP02kZ+/s/4X/CUaSBJNNQ52nTU1bftyqvkdKSVWgW6Fto
CSyI//TnMKI7/ANKjyD9Z4O+96Jy8Midw+qaB+J+Z320ms8gGBaVRO0BEszTCWPh5yOUWpsaFpMx
cTEvq9EyC8GIv27TFOklpZ3XYaat20XsR2MleNGgZq1nV4N8LwtmMrgHn6KvA44TJoXfgvDCxg6x
N+7HtZKJi79nWU0TJtVA8yKZF74XhimQwhrJ7mP0j5N8BxM1mrZ2UTC3q6/ido2FaxhTEL5yYYIR
jteHMXZzfRrNnw+24wpR8bSWxxCHJ+fCx+4YSPK1DE2EtVhYeh50mAHwIHZTNKbv9mBPO6XvWQaR
myluZwWDlza58sh5IsDNFmmiKPiOamSTq39SJK7QIYv+qGf5/2JiVK5+BmlEPXLb5laOw19ELrjC
3hQ3gk3tBVaZabvaznQa8kaRLIGBvgyMyiZSX7ZaDK0MfasXWk+K5nqVH+/+C+OjFOvQ7s7LThxX
9Sf+nqonw25U9ZRIsilUwUHZvUzehF0+Lf8BBu+YIiiidMHtCXrDGJ23KNPqOBT4xuqZmJeMqG5O
+UQdVctnL4i4rIacE+06aOYWYR8xxP1WXd64YTMpN0duK9aLho2BTYc8Hoj0cjdDCoRjMo7nJZtz
kdtjfotEVniiWjVbFq8anMIm8dTUq9c7TKrA9meU5LBIuGzcQWIrhTzBoKxGJ/uujzWb3JctxURN
oW5U0E3DMHn4TEuNCI0BEPbQyO/E4XISGEEzUOld47tLyUjqDy05Y9XI3eB33YZWhIwODbo9BUtz
tMYWMOhYl45mWQ8EYq5/TtTaa4RfCv2oyQAcYS5GGRGtiYc6RuF9PKy94uJ7Nb+32BeqsbhFhsXF
n2sHRIz16yb5UURzAkAqMlwuBCzu78TILowH8Bhp4bxgdmikUTxePWZoJQzdTVlez5CRjhQ+LhxE
AYiverUDk9LA1yC2BSogP0rEp+/o/RD70B+WEx+vCPcLa3l35q0wlgobn/Qb83RJdcfYgjLZdKw3
lR3/RSng7IgdevXzlXdoBdhexhihcQ2jxiUMknPcOvN7j/pBeW0W8mnKxFzvxy/mzNRtB950THwV
WjVpuoUzaW66cuWssSxZfinhStWSwrZP6xZoUxf2BRZJXp7vfHv9Jj5wfFfVgZ1beIARlwZCphDi
OEWkyGgBMEcZX8g/oG8TTWp0WCk79BScAzg6cNir+CGJmk80Z2oFN0WD7y3TWVBnn984OBxgoVww
t22UbIQkDBtN25wLl1+9ieIkUn+pxqiUg0LlFdatgvWiUQ6PO2QZQczt5NBnasqki0m8COxWCgsN
0cBZB+5BYIPGKXxq/gryHu0Nu+whO70goOv23IJAFqWL9tj9sbkUWFWiudEZruJfvAZjidGIDJDW
LOSSKkGzKAX6mcAzSo0c0NK6cwqNWra7VAPRm1/231j1Vey8uCRulvkvNx2VX9YZOfCUN6tKX2xs
poSbMvO6u0dgNX+GuqhkeCaO3uf/BS25N2/SzEhVg5R6bTtC+gh3nuD71j95jbmqk4idBE6fCJNd
t/jWkmDLT2FVYFrsO865LitIDpo0k+hH1FMPou6HT6Gtql2J9n2eqax1brGhR01BYnxLaq3ut73i
pdzQc+PyUhswJmuWfBnbBy1A/aJc+BjBGbvxLRbomHdj+giqh+yxEBufOTzsWK89roQtYoidcL9h
MczfwAeQFF3opeNc80sl0kCVhw1CKqt/kPX7jITzY0yb1upzLiD84Ai6rWveABsZVitkK98covZD
nXiKRt1Be7iSp0RBlai8KXi9JDraWSruCPKnRTaNhyt4Ab68AYtPOyw51oQcxEkYYrupTT7xM/rm
69lltl6hMczcdWnl2D9TyNNtFUv1ogf1nCd/v5CFJjC4iZBnCmB18+ix4UWUpLQaJ4zkhfqvfPKt
qOXCRwerS0DNBP8LkDP5CjxvCVuEH3WSmD4FD0OQojZUJGB44/PAibxwjNKNuQKvFP48WL0x/+kV
SjINB0+xh8ExWKlRx7vw/+9AP8KZYykZiwNuXKxnvKJjnUOYRnjP2Sym+RaCG8bD0uSVkj4W9Ls9
+h2y9jGZbtrufhCXzQdryAG7m1MOpNdupT8m9jXt4vBD5hNrwWQA6O2Vis0/YpVRyelLbFBXPU3H
DGQqcgZNVVGjXPfJg682HiLfU52VdknELzBXzYfJmvrql2C4Da4LqFwm6B9TrWboKgX4cOJLjcJi
HeNc0HCWwWWqVFZKkgXweGPCoOBYhPpl+GVy9F+mMDnlWWfx+a7bl539PxuQ2XtDxSbWLQI7//u5
BJrWhjVSUQxo8Dkbq8LOmyKiQXm05yAFUJcPvhq8UZfYGlsH8mpN2aH212kBnA8JGnQ7CATPtg60
xiLAYa6x3f1Zz9AcydmEq3ayR7e/MpvCXFvFsUZ5VD3IBkGDtkBVvT7jS/sMB4fd++Dp+v5PupHO
WJ02Cqb55PNLp9+qnaYZv44cXDF9ONrOfYfdmCTo7KJmxzfkS9ZEjPSW38b/h8L5QSweQjQMYmCm
ScpTUgL3ziNN4DTVCCAlrabVfdf4MBBCOPMDd+altYw0i7QiQuRmHy5Qkgh2ALb9caa4cblwEag4
5LDBheWXrjwEVXKlJA1iTLkyTipk53tfpzGZJjJPdn76p0CqUbj7Kiecn6FrlzqnjO7ROOmCAjLf
eBSSkTgaoIi04X1O2Mf8W7a2ZzpTLeYrUIS+5rQ1hfwYzRXwjo/rvjQWyhqfpV/icxKs1TsMEnTr
QVCkpqh2i2jbyihshNAv7Hu6fjKMHoErpjbz7+t5nS1lyy8fMVlRfHJQ5v0Hf7PQY6TggwXH3Fhj
enAYoD0CBfSNDeTAdROzAKdGL2hB+mW8stcRbUaCdOyA6XwgCb1Xe9oUpQF2+JE8XWM/SJy4Vc9p
yo7Lbuyd/ftYzhiKBKxQ1Fhw6uSXn4s6dOyLKq6B55noHpOjneJLtFc3rP9S1m63BkzAN7N7B2RJ
OgaDR4KGhMWmwytGxOQM3jH70FKZkkTNOg0oBcSSlXQXfLC4hY/3nyOw4uamyh8Zf57sY40I11Ny
8kxwMYWx7BVcxd9SqvPYxWP8LHtEgZzgy5qO00/iTAK95XxTFkBu4GDg83v5drInbvN/shGQC7Ca
xJbSd6G0kp0de2XxsLQNL17r+GUQqsky+xJ7R7mqyWFOLW484dqz1O8URqznzCu3Rnb/+7ZAtfuX
RN6FinVX+1iOuu/zZhJFky9NlF9D8ese9ZHSkmVhinbwWjj25SZcHwOSRXqjpSCeRWIV+XKMGNq7
vPu1Hgx5PQw9QDSD33bbHHViDlBT4krXbMn4VQWHlS6Ih6FnO3zbrDthSSLe0ROF5rGyk8OYvU1M
95GvoL8YOeZ6MkTIRRJ3FgWXA+JhPngh4bGZv0Z8gzsgsEBGukBv1Rzclnv86oFtH3JCBY8yKRdp
0PydeKtgFZDMUxFAnoLi0oVnxuVvkrLqw535cIPlS7u8CxrzZa1ADd7GZSGmg7UKvS5/7wq/S/Mh
82nESYozXFW92dwqO9y17t4rnb92OtVagFBkWkosRUm0Oo9rK1DNdy1x+n9+g1+UZpgI0bdAsAqC
FHfhoatvebLg1Or/dc+pwqQHGHxqHX5pHDHR/BMgk/riOufvqjCtGxtxK0dKYEy9tOzaNC7hldes
cwffym+R6ymPkTv+EiWqBU5miIZnP2O9c4DM4Oz9XQl32IVtp+P5eNauCK9PanhsEOySvAZgaxRe
5lXOJm57YPMv06fBuD6i72mATL8m2ShNu3qw4104Sn6LgoQi8BTF5Ey/K2EEP13Wy8ovddmd52qR
EAwZvNNB+up2pD64NSLGPrksCgkKF6TPwNM5ySoqCJjgTnq4Tq6Oi5KZgqUwhoN166wluUOjnPM0
pHckyerkr1jAsmclo2Js+JinzhteVzNmQDrWA91KMcnx/oxFtI0ivggSWgwUBjmicskU/JEp+r0C
kWd5hWIvetSh4Bz456en8n7skREL7wrumP07GSUIeD0V79NUml8lZzWEAvcpYsFW/RFyPujN+7rV
9lg3u2NuW1wG5wi2/7Hf/fIYO59IeXVkW2rEPr2jpCoxf+WMC3RqoXY3UDYqeraUdi12hapEd0YN
ZY7X0UaVZwBTiFidiST6nRIR1vIS7T1Ckp5ER/H+kWVMke8XU5etLfSHu3tGz6pS1/MZ4uwxX6fr
lyk+XcU3h/GBDd6ZaqlwCNu/M9IkOT1q+X2UWveV7eOk+YtaSAUxjj8R2jQLQRKcOUBrLb7/e0Ic
PDeiI+a42zjslpwh/z+H0DCn9YjFC2EZz+vzOZXwlb2wv6x6Jo/njHaPGyn4EKQNf3C/c/aWLIjm
k6QVn06iI/wyagce+I15Xr3PnBfHi9RB50vIGQDypduQSoNTVOcsa4wNtLTLCu7ONBWDSo0MrfDy
T3i5lJuWYSaIVe4NDrKraq/zhm4m3/eJtOlqf8yKJVNuWaIDN6B86QJoy3lPHO+RvP+WdRsXQzaT
8Ldvn2coPcgmUdb7jsRFdEK+WXLv6h7JOK52N98UTKGXciW2BjPSQVMIpMj6+JPyjR9QX3FcazhY
pp4w2dukSM/VGuQT/71wWKLWF1+qcQye9Xro01KrKp2KfeIFIHJwVHnO4oHphji/gPnYZAh37ILt
Ha4xN5CwV4IbnOj2rnw/p/iO2LwDlsEsI+rBNZsG2ZjSWd3hQarGZO/wV3N+yMbTB9q4GP/TET0Y
VvaxyVNulHdyAyYcKIbm3wa+fn2yNT5JODKCi80GY7GgD5XScjP0OquugN6yFKH9YlBJoQ9a9rfh
PAVtqxPqSgLh7LtTGcgZnw0km3sn2AG1WZrGMg7DcbL32bjv3Y282g2zKF5aV+T1HX5us1TerP/h
2/SgRT2rVcPF3h9/PPAmG/RJ+N+DQpyygvDpcyJQPODUoK/9cRwEbgePla8jaT+5o73PIU1YiDbU
IDtIA1LUq54tKufDDS23b8x8tjaM80gjkDQKcRhT1xfV+UBirKVm3ScGGxUuRn+Edt+1c+bAP3EP
WZiA5/EMB+WSrPFrwJ/M0U33daVwBL36vxnBOFcp8EN7KahSCRR1pGEI6WCvsfDk7NShu6GheVvS
1S6Idh+vrkT0pkt5jIH9C3nRIGk8RaNSchfy28OgAFgtG9+PK+JfGbvGjvMUOE4VHi7y0GN92Vca
gLbrjHFsIg4YlKzHO7IQrupwRZxWJIzZzbHyBCVUtSucsqRgiyx26Ff7bsCYwkqut+Z4uiCf92To
be4he5IgBDmVs29j6JIBINDMcTvy9DRyMXWN/36tlFMdDSqbXw6n8Kenm0aQ838FlsNeYCPV7s9P
csjpX4jYVRTJbYgFEShPhW7qbLcEYdBJtuOqZxyuR/6eJ4QUlwJKLmFSHMqIURjheP+fXOHPserK
fbgskBjmffQXG9zPfnBYgDETehFZzhDpa9omANgBB3V/iQ3FjFsHFQy4TaA8t8ptVX2gSUIgH95n
usQNWaMZoN+lic20LTIBL6UgMNSOFHNMf0fiO4P5gBkRrjsFWCgEaoNXqonzKbfd+Q7+wbNUL7Pr
RgWYj5ztpIw3Df6ALrDW0Sou2SnBi+7Byjy3sl4hg84i7tMwz0As78W+PHCRhEwK5aspkczM4E0a
Qu305ZLRme59gd76QtlALpo3n+qCjldIG7loQOiuPvJlAxKTV/LWlV2sOE1iNZz3SN14mlooAMY0
wVNH2xCPQ7xp+1jPzUC/meW/8DZaAG58sLJqG5GEva2uVcV93Hr/+Xdqejm2MUOSkBfa/0LhUlix
lAte6JmYYqcMDYgtlsm1W9rl9NoZ3sevGyq2Lwd6Ux5Dz3MSQz+YFR4NxHVbrl2YNxDoDyAz9Hjd
AXJlwjy78DvO2QFMCPkNu1CoEFATacwQCXnQJhTt5b5BZ+SO9QRgBy32F4uNzuNSdl7DrxjcMx5L
72TFp8eFRdKaqN3aOVMQgPkAlpLnYO3PErOKd8thNv3Fs4x711R+v2oSmSydUC8WFeIhnue/uUVj
88k7PmzSBAvyiDIPLGzQpVkeX0KK2EWnKcYSoetEbTDQDohAdTvrEX7a26XJCCmJ2YoyARv0lgvr
qWR5e+GZeYGwlnDsgXFEaDG0Wsa/AIJ3c6GAaCZhj4uNfIsWKT1tRSV48lt0hDz9LzXKeWC6WFYe
Ie15V2rx+blEyszEZjABBT2ES2TpqXY+zWsvk3c1wW6UCe5qUxKUcjzhN4Iu1mSgSF2wscGSE3sQ
JiwdKzfPDqDgxvrVNJTrLs94V6QXy5C6iND3tJNI/qW5kHjFqKmDwHgdFf1gl/qTdbr/UPSRg3ip
qJuwIsFgw6YiUa5a/N6puPeNQ0oM6a8l1fgyQjUwjZM+u+D0uEroD119sWCs32gORXVDHuPf/UIq
m2bbFIQVL0qoPgKBKCzjpoIPbnOhaAbgTOkC60kymkFS1TnI9T6dNWfM3FSl/zGKYCAVdAaxCrAs
aGLC/3FPaERyBFij2m3RA7oBnT83DEQF+JwSGIUaZ1ITJz47J/vrrTHFUzFEIc1SGAW/AVcHq4Rq
04ekEpTZ650DmwHSOSHnC8cmPhbYtR1d4kdc4gS1nM63M1G1uYDnfkqeVp+77fDDP8YVY/5CwCGq
LZJ9Gyd/NxsMnasLXkxqEhOr/JEweJZelpuf/mZKDBd4jH8lcn0mrVa9lhe9Euyova80JZCThaDr
EutalzDJ4CLLLn3ysNb97gt78QGOsVOCsfKUge3NTTrZ9eAYyecLrUQ/YD0bBPcIceJNm+wF1VxO
yj9wJvU43KTuNaQ7OfwX10fDs1xpmG5P0kOkDzVtQ1m4tTKDdxu4xYDrQdR8W2QUpYQAplyd9mER
l4Tr/I0ltcJxsmxGS2zxqqLBp1xs0VFtbcr6k6+6owedTKHam3E4+peggNMU1C72+O+5Dx6oJhha
j446zgDuoydl6kX2xNLN4WFbYlww3kr5Ezzvn/bFLyRKnZ5dQLnWGLNkEc6HuAQgy2oo/BPu0jXq
AGsEfXrfrBO3KRplcL6G1KubcBvzhBrKi6O3VfFXzpRrVRvtySEjycFVTEpe/XiBRoonq/ngun5A
fFGfCYOL7hfX4zyeP48od5MRHAuCtZsPx0z+3siY9HCENQkpGv+bJCMbQa9ow5b+TlwkxCr1bEmN
bOoMaiuq6tHXOAiF3SRq1dW9lPWSdlg0XMRn9LJnwxQltQWGxj6oIeNAJX47S+EoaRSjqBdcNrkJ
9IwoV69gt3fDQnzaGCw4SM1ThzqyVIi4p5utvL9k+K8XdaqWryz0WZDnTNwT0gA7PuZ5NtDcPMSh
oUkYmYIiaXPdDtC7slpOy2OFBYHKIzvZVMBDzJF7bR+++coOykmTMkQw2zs+ggL+ALu3b9Vm5yoi
9OglSRjNgjaEe0QCvYjTe5w4prlA/W2vE4aov4agQpIXlJYYilz8aFXTdi/u+FSX7mdRmWBYicNy
deGbEFTxMrKAKFZN2fn9SPBNxjbXIvRhdUKVB6h+kQMOmL3EvbL1QRkmDjpPWVosPIGiXdUQMXmg
7LFWxAxl1ItKprPrTZpPK9c1XUIfIQrQalcQSaUo9Z65u8E2gw1aLBW7IlCmgSzDU3TmVFq4fLZ/
higS4DqywQJUgAjqfVumO+Qnc1MtI5eImPAYTdSsax7Pz3LlefG+ZAYzF49rQR0fHK0OKj+gFRT6
8X7LI6OiKqo4WwNAVI2B6WXAbk39axtmBBX/qiYTn+oWOgZmcNBbVvdOGJ69+3tAyUsjVN1FU91h
5YQ7hxhgBuJwO3avGG+12WvAfJ9xRz/1V8wH5/QK8yiiEpT081f9VBJy5evL2NhoxLOKUL6rEaIv
BHv8MBF4YOknAwrsTYKd36xdOD973oLLJ8ZQyarO+jTfb6ZfD9aK7glYtCwr2HacIrzsZM7lqpd1
MUUfcwqW2SlR2U1R91ZIU//UEXYHJZzuKh8LLO+0MG4Zo0Atrz3mKyFZfG4R+7EWcmSRz4J+3AO7
e2WOiXj9vfC1KXch9fa66VKJM3/6okVl2Hjpo1UY0Xhyakll8IXDgExJE8kEAgKYP9dzCc7/scfE
+qNJvZE+6KzkuPvTJgG+IqZ3Rpg54W2aqOXWqjbk0kMJXPzu9IDEflNNVf2ybUDYaQCGLSfpQnZ3
VGB49w2SbyJIEEpjja0sT7QQB5Cup/X4ok10uGLES/gfZNLkwX3Ar4psq481r628uhr4IqmKejx8
zPWzEXAp6JnpaGFUhPHAwfo0WtDPJpT4hf9iT6WGCbXhqOo0AS+J4et5SBskqOSVfWSLFsqFA7kn
jNt0BvSrKmRos9dtzzZhbmQ8Y5MzsSPp5rc2uGEjEhEsM3w3F4z8SIrJ+tTUQdp6Qa6kSAMk2YlM
qGyRNEBdf+upQJIyDCU19UCrqoTjq+tLBmU2Esa+YHOVbYdJPO7ytuoOYx+5uMKC7IkI70+SOcmi
lCE2sxuQUzufi4djIttPJ/ilabFVeB7AKT9/F+DKzoC2PK9xbUXgoUEEONHMiX5qrgU2bsj1uNsT
h5obFcKTbeOxiYxKIcUJi8i5nV7vDAKC7NhqRFry0f15rC0lza4OgkecPcfT8KF+lUQTXbwhJ/d8
XmLVDEJ+s4IHj6plWjTaL4K9tjSJcOQj1D65y9julueGUCO2defJIJc0rF+W2CJQtFlqZNuQlLZ6
pcneKolp9+iDsMfNMS/0A1Sk90kSVT53uHuPMaBUclxJMY7+upVcKC3WZxMW8CMYI8ATQ5xCXICw
vlalP7BIwGUOTMt/34BnnZFZGc9sx4JGzkMkabMpCFs9+g/RWECFFScMAzS4ctN2g797ry0ff0HA
mHCOSP30p9YIK1PwWyORvo24dBwtUnnDFGnaw74xqt9iOCnmwfFMRRX419y/iXYtgb3mmvaFqxDY
MHrafuLXviSW7NR8/l9T26qBzDhMOSLshUwNhMN5rwPM7k3TeIg5YIvZOT4CWOJlqhxla8CxzJrj
1llMOPHrlntopoVV7ZAHQpaT5Kr5efS8zdGpU2+B8hwoiok47NWdYzl4laMepj4USO08bYghH8ZR
7zkDebJk6TpCiGMw5VgYtN/RIXcWaVWxYkSESnpWJP5P0T0Eb6xMTUkn7I2+/+E0xiubxrLIy8qt
RdyRmTJLBNDNcEs0dxFvPMYcT1mJp9WADHE9RGX1r2mXUSvR6JFhtpwdNfpRlxRj+EiOpkNr/dVB
nPfItGXfaUD/4WKiaCfzIUps9Wwp/G9wTzU+qzYBH/who4IEr8GzlI0CKdvFivux9XGyJlBno+kF
mjPcio2GMp6EvFGjBHOhHaFPMVxJZVY3a2/x7IU9qacyhOEmGk7+2GgRjpgYz1dNMSJL022kGROk
k2p0L64p+F8ysWo9i+jMp+1mIBNOUJSVyF4jfIq2ND/yZKT6vUGrhmYoDg2sBm16NJ7b8jyg9u/4
yqMQY+AxuwYfXIKsm1WvOdQ7PJHpYxM0EbU0ohk6ruWaentLkh90k7g0CEBKcYPRK7ke9f3mFnaS
Sh6mI9Fv262ylhX29QLZaNJUBzWUVEath8gsi7fgAWWjcp9VtwJVNXr9ANHfw6rP7zOHFeaSC2Sx
+YTFfKMElRpHObZrMJ4W1rs9znaW/zytofoIEGJmgkKc5Eu0wTi1GXZVDcyUZ6VZg5cJP90HhPtd
TdzTLkSt882HDsBBlmR2hghv8PIZgfw54gTIG1uvZ/MUdir7p3w/81HF6L963C6hLhfqPQ0zZ7gn
oF0hh/joGG5s7q2DfW7vPSPoO4gLwRXtlMlzHPL6B3FIYcwcEJdtRCOKHbxhJCOCg04ZPBtyEwTa
eUdPmMtGIsJaDWK9MgRyDILBwnHA6dtKNR/I29wKP7gZwlNFJMoEd/t50Xll0mm/WNEPb+pA/13b
pfe0BPwPLTPDQ9eBm+HLWbkb2nr3gu2peOERHJliwlm4vyOJiYKpRd98ywrMvrFD6FOjv7uO6owf
w/3WhYhW0r3eUIzEA6cErUJvzXbLQX6kAcyqmh4JnH8QJaiGkatCU2DlOfeY7+FCR+TZs9X1uEDm
mo3ThjjFzNetaMlWedUaoPmFDpouHtyIxDTX3/s1n5JJIzzYO8SfhV72Ke27pFog1xpPhFuizN4t
lp234GwpRFbXfXeqsnuJoikYHZLrYmf1ZWszybxJ3VTkw4JGzKNUZdRwzPDuP6iSFogOoMX5tvHx
aYmEgq64v3ETwYOjA6t/RxtlSzyWEIubKKkExE2xd7wStvdDdVdzH2Y7Ze4f/0c97g1T9c6T/Cna
kXtXqPeED/xsu/Tjuo1iOm1Rnjm6eUJKth/INYUZF2Cjgi4Cb7Vnyfj9X3hQSFBbpel3sqtwVVme
3JNhCW5isgOlchVvo6OCF/FamKOchWL9dB15LuvECc1DRYTztW9E5TO8Y4561Wc018XleZQZztah
PKzXD/MXmljtcx5jKXjBBLrG2ryBrO6HECKyn82zIXlkNjOA9l+kSyUhRwJhQYWhCjv8LmbLXxpP
13JdO20I2CVBV8cEFe3aubgOLSto6Ul2CLM391osPjblglA0BGaShnYOE4Grp6NDZkG+l05Ns0Ke
bvlupzd1JO3XFNLsxr5yPEIMfGf2yIjQUs6ll80SICI2CDmzzESSuMlYSOzQpnNrPk1HEcEBfCvy
efZBCo8igkrcjZRYPt10kUp5hprYvRB3dp0uUpRkIrBK231LbCz0JXSMkDhV8ag+VZThivz4etKO
8wkoVcS6UWRPQ4A+Wf99DnRo/R4+ytZ1Xys1ZXDYE21JS4MQcbnUkNY6hWq7JeYxTN77zN7Ygqje
JkL2Ngq27k9oHpDFLGid2D38y/3WLUncgqx6YcSdfhT7t+BHI6hF37SiTC1Qkw7qBYrGwBo9o4Tf
CBWCgHBNIc9xdUYxq5zLA4mdxbtJPsc6MK0cHH/hMIMoVejwaLOETK0Skq5xvrbQxgV1B7/vdAfW
G943OYm2O7v85y02aQGAvJNuDtJ2jg9TnbZ/GzhEvYW/Zxv2gCn5wv0Q/hWI9SJnmckoBPkskWKK
Hciio3QuxJhI5WlmvTwLQpVA9hIO/NffTSnYw4LZYzdVyke79EwT/mVpfzXxcpidBzOhJuotpI2d
hzoE2nACV853N81250vFz8cTMmS7Qjal2gJyfIo8mQYGW0kSq6UDTUaF4Yeig8wOY7NFeBux2GMa
FYl4Uh7z1/iifUxcsB05NZBfCR9KUdNhdoJzOvMVfe82US43q52euV6t3k3e3y1jTg3WdfrQgv1V
sUBySnY79ZfvVkg8sS5blV7frFkYtclidlpK8wj1ZEy06iWviYSGyoFXtxrGrfpuUjXae6TGi8yz
M0sacTyuCHOa1pgy5OCBK9rr9Luk1kdlMaJ/VtHXdjODD3iMjj8J9tanPZHknGtScaS3+MoPVUci
TC868rgzTLM1EnmAwZ78QpowWQr00hXN6RteF0fyOKE8vF5iWRU0aJp3uOK5bXBdNlT6Scu36EBx
rFFrP6oeWVg2MUwDKhioMPiOuqCeGWbhTON+Nn/ytBdbGF9DRH4W+fgYUzvoUklfRVUl0oL2GQF1
qOxqKv1wTyo64JLHmGLvlsManKQv5xrRnHy9TbX0YL+1k/PK7BvjKCGBQ47+TQJvEW0cZylUb7pX
FYSV1g8VUtoV0Euwgq4jFZ17dgDDeOf2uViBwqSgiVm5UoxTuekTYFPmwiUPmz3I1a9eE24l8Wvy
wD8+9KVKdjuBTop+T00GBZOtywyHfc3FfmbVXtoQ+4gYAE/rHvd3W+ILtIi6+MGkQ3WvpgD6NQHE
NfVaLj0CWb0rFI21oAd3yQVNJks6RBXr4aM2S0Rd6bxgMTW/6OLb8goGHWUgPpYmYur5Lz+fg8NT
sjdgKaT0Xrvaynyk+QIkEX2FBN10TivkMh1rrCBMwPkA3/JvzRVYKxGqUf/lTIrovtAs6zb2dNxY
YmkWUY84zp+EuFh0GOh3gC5KKccmA0TxHy9dMfg06ZMAJr8dCJRPD1Nm6jfXTtcUmODy+QfFYUeX
/DvfNPEPaa80MeVFF8s/iYj4tXHzriPWaEnX1IYQ8bNxH6OrPRvoXBeeAurdQ1smpsKDN3deHI1P
rO2UWmqZdFBXxAeM8gffZSv/HpRzRrF9kgam3ZpCm7lCdvlIjeNPEuJgtSnfhC1Dt0TpllhnOitR
7v5QVdMIFQYnJLCf95GAhliQM1o+c47KYxH7G1Gh4S+1XXgX4X8PFtwjJ1mz0n6aRLc82Gtj2qds
9+cpABTA9WzsbH+JWVuXgrHxrqLDIzaaRshmKlAAJR0jJS0HewQ9VvUSByzKq0qGY/Z+yLKQ1hN5
SmOa5mSLt2Ul9iTcqchoLhPDH1Hiomq9mL6+cwNvKt3X9yLy8MrrSWK3MQISYmo6ynoAYlePQnwL
ZEoEztq+FWLOLpecC17VwSi6/iGRZRzMmI43iyYcJZSNBupAY4QWzJomY1tSxaCKoX/QABq3l0jD
OgOsbDH50z0PZ6ql6YGY57K1DYlvlEdIcJHETYOhsVQdSFq3dZITpZssojWub5oqXoyX2wFZbsMj
fDOWZO4eH9U7b6b+0JxED2oQJUqOpmSmOHofLNA2gW0Ekr1eDhvri3iK+Sr8J0vP+xBzWE034Y6K
oDmwe7x/6YBljMVg0I0kDp/BuD7m05ty6N1p6UJ1zDQSgMk/4mzy3sRdsJwp1MY2VkXe04Q+VlOm
TqByE4sdH95mqNapABwngJLRoFChaEhJoDNEQ50Br+BAz3ca8A/rmGBKhsKFOnulYz5wwptBdeol
GTGKSe7g+cXdA6UJF3CVJcxxfumn0/qWT7e7ExPnuzI/zcov3AzLInlqTD82c24CC1YDWBlpzsVF
/SrCVtkhrT5BDG0vb57006tt3HorjybKDt9k2UOzGkR1hTla2kObsxedPJQYOy1PLrci2rqMlXPR
DgCcZurRCRfiBhWb4Es2nuNo2te466QTlr2YZLXhrP0nvoz+4VPIjEaTslLbmvDgTMh7BfaRteUo
BObyNvb74uQj1fomnZSrb3RwtRbFBArIJW6SCwanUuw5D5BTmqeiN83aAvjl6UYCCtcJD54ZjOTU
G8PdbrcyNB1NaSgkGkaO+iGxf7oQJX4SYbz/vLN1MmQiWZFrp1Ua84OjdmoBaCAHQoK642+Diaom
BbbENn5z+9WkUtYgyv1GPXjLTTJGdBI7wpAeluvjD2h4Mj+fcTTW8qoSOpN2S/hbggxsbiElmJtM
jcOQUqkkOtshY+NNsbwVooh3H0wSOhc7CpRlWefKzPK5B/rHY99fQcvoXO4hduD59k6FSEhdesIH
nS8CvxeT2jxgPVdavesKETvHIbDagMZ6tFaMge0O+O0y7ogrrhXI0R4AXIIWBG6pPio/U9UuB355
PuhzQlD0S3/dhl9QJSqkplnqmgNvVKT05fij9I4yCgi/BHxPnX5FXfn3YbKKG2TN9qbANHZSx13R
x5XixQusD+WlJ0/kheQpm2/vCWLwUyPAazNYnfrB/WRaGKFOsQChE3HsMdZhAddUpOV1/B0jPxgC
wtmZQVaAoqkrqGbsqdWi7+NWLOZZrt6yldAhv8/mZVneYk4WM6O+/XCwH/zN3h4mOswDkn7kVLSr
XhF6TFsbJ180xy9/NFoOxzZW1+pu1WnuIz3Hch3m+1RP8+49kCzOainY3vX1YCeUB2nKD5tm2IMT
7PBx6SYiNlvN8KWX5Q1SxKFeaRKGcOGjfQlucRAo+WTa4hO55t/BUwlI+1BxLjMxrDwE8IzBYcDb
OEivqZ4ye0xSm3ElG85bn545FdtKh4WCacR+ZKhKg3WAjeCMjpsIV45DgWagoyOj13zGacNoW5sU
rO30Yt+8T8aKiMHt2/U+W+Xyex/iqPZyv7OKAlYxOxw63XpKlqgd5q+5gvY7Fj7O/q/M5L25XPcC
b/FZ/xRFKmGxu4+ZKB5BImhoQOfGXaHmqV9XzNPtN8Bg2xZ8KEpIXnQmZWEwV4duC1Em2nf8mnrw
0Wzqad8uruUTyMzH+Zo2m83iFSO9MSYGTJWR2gh4ypMMQHDvCcHkZstDYsbEfexBI6IO/+oLFMQe
GmrYgFYwOLaUlcpa1h0rzooNaQxA8tYinEvTk4MvhEC8BZ51NN7uWaGpcovFKINVqzyX8tesxQ7g
lZiqDwTVStspC0n/HEAiCQlChms6jGWH6gymESRtbXDtIqqvQ2NS2QvmJQMl8dmCMTYEzmawD/Yy
qguDpr1CCpZ3abYclSHMhfUQltaSOvdc8acJhI0a6762KbziSoJ/i7DAYxsREGTN73yASY6kbJhB
DhAWPmbp69L4/V7kvJgkBIpZpUBivqIGwi3wWWofXW9Coh6uKj3w5lOqSyNqQum8+VQmugyszZRT
p0BvHJSzJDvtdYFOvEjuZmKhFwKws0uRsZPtrL5fHljeqNstN3PjB9oMgRYiBHBvw1wHyK4rht4v
tD57f32iHNZtQL6zpd5ICbzMU5VWr/kdGf1Gy+7SEDvyI1Pfe9NzY5xuJyRRrCpBp/M/gDHjLc6Z
oIXNQR84CC0OfeuM5mb3mvgnAlh8esGsSaUJZakibeBUP3ZvfYb72TCX/DkO0QYm9xQO0I4NEukR
UaNfPSrnq1E5ZsKrBQTOQwBNCyg9uQbGe0PV0CwT7gDyMKD8kkW2ELfkjk5XoxKsH1Y9B85dUYtS
AfThxF2m//o1cO8wJb4Jl/SDZpoLDLledJ419Vhh+7yceNPtqz3oBDv+JP5urzNSntZcNvHJ0tWI
gFWFvZzvU1IEA+LA9ufGcpjMx8xAxCXOk0yVK1DoGSjRhdSb3NTyGL245nzsUWt/I7i16iA+mfPU
1IClu7QxDIpOquy6NOZH32Jvu/plGYBuiSIXR3u+KIbLf/SBROWGa6pZmAQOR/+Frt25OebRAuqf
3204iY36xcze/A30O8TzBeYeeafeTBx3PnYvI7/m+SKi7pUEMPA1D71rBRyItKHzTQnvtW1VyrZd
rPz+9fmCTBTrTjeVP5nqCNXzxsZ5o2S/cWGLUj3/EKYQfQ04hhMTAnjgvnKQ5mfewg68q5AGYlUU
Vq/8vdFSUerd4rHF/0e9YuofPKjdQSnIOWluqcLHEJbVWPnf30tuP7L10JT2ZdYnys4T/pkU7SJ0
LKK2KMVTfJIwCs4/xO/iEIq3MQUrICLdMwE8mMESvaAMmcZRI3+ot88zf2iJBYDmLzgyqmeMwvUk
7Kq58wryT4w1GFThu2+ne8Tr6URxxKoBvWUZXNDq1IDCLQi2vWEWrCoT2Ef5lneN4+tKbQKsDEox
vkTkIulRiemvi1OTCHNJfbnNImz+ZN8vl3uvbOCVrsBw8Nj1tYnPIPd5QoHrbZ3JIHrnIy/qacQ0
FM6U/5DR0GbzyHtD3KH0hl0IfgGyuzCB8NxsZb2MdjicUrzz7lWX0PbDRG/b+X8+sOhOWuac+W/b
r1Q4p+GuIDEO+Y1X+Y91cSOSXngrfEzaMQdFr1GWgG4+iIgm/VN5zqrLIJl3w8lk8dlIGG37e7J9
PByxqCbPmAIIoNfmhr1tIVfk7HurdFIT6Tel1vIgwIw0SjQMBWpNqPhAHyyIrs7qDg9BzhiTyfYf
Mr0qM06Qe31oJJQnPnzKTJKCWqkA/bDj2ZacECuqJmC6589XJGZFymwKsGKUGwq1rewIpLVZUF+T
7oH++MLYFExhk+0MwBom/dmunD0B8i4+QmENigf8WqtlMyPb6rP508PVsPDWrA7n7iHTiYWJ6sBs
cyhjwohfcJxYp2D8bjg0/tabsbLet5+4REalwtIZ4swX7mlnZ69ICwpstZW215xoIE4YFjUHYKQB
UOf0CZnseEFYkEkP4okiONvDFUFwhNpkF9xCPhvtF7tlHy2ridlUlX5N6rCCtmJonPqOQcECS0+x
zJ7gKWDIFFNWKS/oeikzE60zJbfuVFRGIqhcQcBme5ozhI/YVOgC6Cdl597XW89Fzz0xQMj8nHBU
wJxjCZ8NXnV6rqvfQ+OQA1KeR41SgwQFVG9nN9fWjOFZmHHg/s+tcv1ISWdEUz+GEpqn8RguIBzb
UwtzTYU9EuL99eI8md7kgjbPFUUDgSmngxuNSrzuQ9Et/yqUM6Bp8gpQggda+kq+rNkf10i/dMh1
3f07qm7FD/dmIoiGPrIz5YH9xXuPYvUoRMMD2drF34JcJ08a+9Dbzv1Vj61sPMN3MfcQNDdORCet
qCkt/5GRezQjAaTzLgYSHU7wOJpeJdA4nZ5F7ZJBJzuhOhyvwKABbMAGOHlYzT3w0LXf12TsRVU2
t+SH1Z6M37/Qa6vLXjxGiwAv0utFpZM4EHEOxJ08+JQUvfZH9evAKTGfCcGpX7v+dIGI2KKDU8r/
SxEZtcGIJwTb4g4f1TOZQVimKwoSq1zKSUgTC3B9WgQWLQO9XEZlykKhqs02LrhoKbOl/5NmV1nG
L3rVonDdCHqeKtmcpuWWXYDsfkSKAYNTrSOKCrUCexvhd4GAgJ1fY1DTfvCHTL3jHwCPzTKVGPaC
V62ZgLCIT0E8Jp7OUwAZZRnPnmVlSudVBA0TA5eMBheBee0kL+1cjqXeSkaB64n/aZ1JQrHIvrap
R3evsbCoCViSAlI49+byWHWDrCKZoK3InHUj7RKwWdyY2ohoCb0EfewIfGTy1rEbDn4lve1B17LV
d8njTRAOvWE3Jh/+W2Jl5aapX68kJ8HTQOxBdTgNiM2HPpxb3EjYYW8/CziwRGEOIRu9KYy6cCWz
XRM2QfF7mwPlTXtHJ5Jm7VemnVO56INYxZGpad0dW6D8p5IvtLskTPkZHj+6rv3zUySn66ds8LDO
IPcyn3ryZurIBzmRykX8IrWfILx8vQVkEgK0VFTj/p+f6npFdcef1OsWCUsnBmiWcUPV7sRmUss5
3u7jG6LDmfDOOD5yFc8pO569ajnbColw3Pq0AoKssQppWPMoTzyMq/XIoxLq4tKZ500Joi5VfT+H
VVQ+cydQNhoYWO2tsDwJzkZ/O69etCTU4myvRo6NWZ+B/B+fnzyicPctkgu4zQV2h/ct0ZM+5gDw
Q+8HSrauvKewjeCdAcqTu1tsP0bGi8Q7qdC/2JA6c0JQPO/kdqHAklGWzPgir/0iTPPjZbbuAGYY
Ewpxuz3+QV3+gbqUBHi2IvkcSSNCU3PKrhD7sqxuj6y3TxJiAUv/XgJbrDdpFXCQneFvXMj1UsNV
gkW9OsCY/iQMQX1CpjYKAP3SNZ5gHKVf814EyEgR7VM4mA2zX5o/Pr/xsytF8Gk4QHQ42xEKMp/s
pgDr6HrHLFFvKCz2B/+wLIVf+7HdNUTbO7LAQlr6I1rfzlovXXwvPMv8ARWSQNZp8fU8Dfm5QMNU
5pr5SjaR7+qOdEAJiAtgtgwH8iO5cj0u2KUEUdIfsAllW0SMT4fCSjZagqwdVmGgevchm85i5+t5
R7RDgkLFZKiCfX8enBDj8iAnU5HNTybly9ON3D59oVov3+vq9dtzbC+2A2O2Dz/k1FqimSOxmKtc
bMnlqagAd8t1iMT4nZh7kU2a08ziUCMzm5Y7krpfmxkM3v0B20c7O/ddw9uXCQAQWgy2Wt4sTdbH
adS9giPhf+crFAEAK8rBRnxN7q+afqfq0Dtp3kgImAkxlvY1MrjbSTKjfuMiCJrD1jheK5x5Xk4p
gLHfA7QbM03jgm3627qXAC6pHINStZgIdmHOhJDKupohtHpDybGg3pl3EOh1uk6wvEgJcJhzRH+Z
+xJfAzulVM0PX2Tq2MSs8Bl7FmsnC7IPyFSN/4daKZsBdET8H8rhHHrGUUk694+Z8RvwKrYwvHkO
tfb1DaFdWZ1XIe21SigiLTKPJ94GbtJowcgNC2QdBjKmkx4pblbLqU9jgGxoRmUy3E5WmxgjjLmX
PbhT2Qv6j1QroOjOfBOLV8JXDg/bciccnA45HGtPYP9q72T27dfRRexyz6fct2Glre4JgP625oEe
2Wnie1JjB+DDTj0HeI1ECHVHMR1SX1VJ28nzCucgw71QuVCR3GH2ed0YCmcMd44TLoSky0Ze7IHs
5FSjj2PwS8K0ZAoDPTjUdXCKa68LqYQLvWqUwbpUjd0LC9LHLSKjVtBE+xgxWDJD1MzragONF/2A
pfVrx26jtPtVz8ek1aUnUKdQVD/O7P1tJyFIWCzL7pd/sQslFiGcl/N9mkHL34+StpmWcw6hN7Q3
kXS/FRihB9Z2agwVu6ROhe3mcGloR/LDJ3ci92rfJjQCRztcyp8hi1u0PRTZCIfIVZ7JTnbd9EEU
HkPXMWMWDQPipbg3QZ5l9iPly7ogwRJNRUPWgCIkyBHEfdSMHyplTmf936J5UAD1X8tBwAhvjoEo
3OfAm/C/KC2CG9zRK56cTacEQRybx9/2eJp0gAvNZbL3sP5iw0IYvZr1ACHXFoUT63Lw/lqon1Dh
4nVAW4xiLWxQvq0FSNCr/xljzzGLghws1vwcXcQNxNRKSfW1BVmnPFwIURb5kCmiv1xwj3GUDd5q
lHeEKkAhYbSP/VNiGiz5H8djlZHZ/+OiHQs+qs2LIGJMY6MKXcptzvo4pTI13y6y6b+erTdhTeFi
sl0Argbj/xfi9K1GVEU+2vfFvsRwP6bvVw770IItGddLMMHsZStFihjrwkBtUx9Gt3qfJVBU8lk7
5xG1/1UvbA9gAh/5Z3sZMIRbIJLKrPE6fn9LPkPbXyC+jnh0cVLDlfWOgDoblVrhvVYGbh3ok9vR
xvBl/tLuKagJshY6pBN9gToke0m/agMhnjS+PHHOn5oDqBMPF8A7SFkRL8olF9eHKFjl9JgTtnRC
I+uPpTcrvUshk7cDuZ54qcPLkjumhI3Hc3xj1X8oFsdw+aMqkpVr5OoOifHPcjLDBXg9Zp75YDsJ
3QStuQBlA7DJg68iKJcDpGIyEDJMzASZyoc97kE82cJxVCLALheBZCPf40hibx3bX9i2sBUxwhkj
mF/E16JYNkX0B7LrwRSiLn0DlrQD+y6++yaYYyCmtKUkAIOU9Nq8I5Rhx7rOf3WBqiNeejk+x8Sq
DN3XDNANFuhmXtL99+xikUbtsLLe7KjToFmV+0GYWnpPlW5SEwhGYUfn1pXRUKlABRFyxDFnAA2A
pRScgvqZRLQbv9oLiFRUo2pkzMMrixq26066tujBOhxU4bSsk1dF8qVOu5Q5H0HwJfn5PzorWXeg
KUYGNUAn3jpyWrTgAdhbC5tjue7rpzP7K83eFvvJgMgzrwhqjz5Lct8z/o1dW0BAKOn+HproqSSj
LmFUXzabGZ/1yFn3DJcMOKAWKiziU+fZPmL6ai5u5nzJlVKbLnya8/C7vmJUYyKQZc9dRncvhwoL
HTNnA97irWQbqmwjtDB8kqjei0FbFCTpTCceTDPAd2uR+P42yZu8r1D04TOHCNQazfLBRodgwUCO
gAuvQ/wY3C3fGgeKaGLaCwTEWgPfewOqLT3uRhQLr2a5unZYST0GxnXoNh/Cy1wBsfhN4p4+INQP
AmMLmX+9CNRfivjepiPNgIptlgt7NZaxbpEQ4/hJHbY9+/uFYxxaqJbq0vZnveRRUGzfkrI8BaRy
Tc4a3UFodiCEOGC9CCntvxOqvIOZtpQ3bmIAjLsNg7+hVG+tIeq3KGAYtdpzETveFfq+yo1YaL6E
fEWJVsFfCJiuDPaGXgnEljN+qa25vbS/VELFw5835tDEzGNdlvSDEJbrKDlplJr1VKdnf3QteAWv
ascKUMzsayg9jhBEikvBIiaY5rJ2M8g4vOL2cG9m8nlwHy/8y/h71SRBle/pSmhafm6d7FDF52NU
qZjpAWiNfK9uSTFXUVpOCS4j242HPwA3UzdFJmcmVMnEiUsBb3Lt0/FXkjFR8CFgsn4SsA2Es+2x
elPPAMvnp0rxoRUnQ1oT+dnnTYkgfesog6TuNum9YzmWcqwXiQLwfK0wUt1AThSEtqapzp0iuk2n
9CYk0KJhpZv3l/+avh79mMS9ckv76DqRTZph+nITxQd/CmEhvedejeoslmU7VF3OGaHI/njrONQF
jhVkS0tIgc+1RRdYkKdvYMGoLqlXFFp9x5eDkHnzaOiWOn53DpLy/CPPjA93i3+X3wedqgqtKkpo
goaQeyrwJ9KZeqmMeweA4YIh789eCKNIctQc83np/B2GRjPFVN5eeDassx3NdUoRCdzQUzHNF+dr
sL9UvVCt0Mwlg8pEDBuWq0iQduRWV0SwL6cCHfMTVvC1ugIDDFLac+oF8ftepUU5dlegPPNQPoCh
GV/3phLsSr2MxHgeIsSido3QQQYpFLkO23CrYjEH5ZiFlPls7EIQhP18fj70e7537f1XVbbtHjZ2
YrzYzmy0FTsmBIj4nxreHmB79/yD4E587rj5ScMKgcZi71tPYQ0/vBU+fmr8LhGnDKDjP2741TNP
uq0bpoluoCJNF3+kLGR/X90rT5tKYf0/D8oBWuUVHUh4PBkS43KdRjyrJslxiZmv8iWbwVitUoZG
HSQIt6dDeGZb3m1kfPENprEIIYVVBnA1WOseBuujqoeZTjC8w3iPKxuBUylYc1YN7aA7xuue7oxr
k/7DZGNF8jcNkPfHTG278VQNP1ZxC+B7xZBB3SmddOjMqF2idSotsZbJO9/N56vD+BKf2S/U3Xm7
eI/RS7ci27J1Zkef0uVSDz6EdE+R8kYR+tMFLy/Tu+bjrohySyinA/nTb5/pVv2hi/Njfu1Oqwvl
+SmMPah9vUdHwC0YkCuapYpZyYWBjA31WzH1kDrExLMIfS83DBZ5SpZusp36Z4xuWq+H9kZ0liyj
Jaray130Fr6c5U/NW2meaAvlGzbWNGafw/FuvCnJdtwphmyuzbNYTU/GYRDR0Lc8aaDVJdTEJQ1n
SeJCB3XZ7HmSN5NuNSAO3tQgoNKF9lzfJ6CPppQzKvoYpB5e/hghxMAvguUYpsI0sx4mTD9jDgz+
H+o7fwxXg8jalZrrvMIp3Ut+BRxyo+UU4xy0Q5uH8DskH+lJTPp/3tkv+z5oxm8lBQGs0Gir/QE1
0DQ/CWLo63zqtz6M+8HLpahreJWskQpr+DrqN7GOL1IHlrY+7kp+osOq7+9hWm1bRAxuE5eNIWWW
/gK/Q6DRykWC0aa9zjXx1oWyiP8qbvLH8qp6DF54EQQdfxf/LL5Kp3sFXntPoxd6KSSs73R6OicZ
+3PfxSALK2v5Lwmt6Pgq+4501oM/Feg1+0qefS1XRFUa8a+32jN8jtdF3Mmpp4IsgI+8sPEWMgxv
KQ3aJFSCMeB7k/jToaXfx27LpE0XydIZs5TzsxyXgffz0wHsi9Jz2VZi2q1ydEAyQRZ5pN5E740a
ewh2KGIIVnfCjrcIm+SJ3tACNGem5tSv5RycBhTXt+B/ETK6VGIu3phwAsCaRVm6E/9DYhzCEahR
XjLGfSvU62dd7y94gKM+rzwLiFglH5/RxGSl1zUBOwMdwzTwJGrwGR+sx+/EDwiamKpg7TiZm8or
Vkvc02yklHjZ/Ra3ld7jDQKDi4PDA+fDDYPpf1nGcmHQGn/waE2tu0j71SX6/CQ9+YACzvRa1Isp
RFpNV2r5pZPuWtKp26enaIZttJ2EAbedn1N6GN0cjQ6C+/HZ6O6MndfbK7u0HBopUkblFD3nNtvR
YkCxoPCHjXJlRLjP29vzVj2zXjPlIoJVx2kQlTtKyOlfgXVJsxVfrCeG0We2PVjAr2leTF0RmzSO
A5tS38Po7SnkwvYY34cr+I9ehAzZfBpSGvaXUrZ/2sCIjqp8lL20PPrc7SfZl3QqZIIApYLrVT6P
TX+KCUazBmbwMVFB0XYoyj8P+iQFEMTcbkf1z/ewmgstfLYH6sHEPqwVOeIf8aD0lazmQecQTLyA
7Cjdjnfq1Ncz8UTADZn2LcYFr7eM7r1jkKC59OoM377AKG9a/zI5DW0A1ykj0ltiIWdIbc/kTIDk
4ErkvNsai0ykWzVxE8fdEjdBF6j6SDUK/Oci2qn+2AOv/lBZsKL+WpMLk/AyJsyOxRQyNm7pyR60
FpqX4ONPsoT1+oyNvB/bvgCC08qC1LzVL1t0p2t94bKxff4JLP5GnPPXlZ86LCn6KM9bhhvWV8Y2
KS2yFsqeFyAR6JtYKCXVzs4elXKJC3SLWdMW90qNnaJV7V5cRKJSwW23DULGAtRsCzw2FW6OcfVW
nsAImfgb0pfkHYEMRrBpUMD6bGUIk7hJuQmi7TICawO1sXcJZxOvaaclIsOo/SJtWUyA2cJkJKau
iPGmxWgvl+uPWXYFTC0gEHbOgD3QDsWj2pI24L89i0yYXFE5bIoYycjXudVrbJIysMKTq/k04yRU
JhPq78SMsxjxjjhlc4deqswhgGRw6GUohERViENZCut+McXnztughFv6ggSl3mc8RrNrOgqRRent
AVHo0KRAue7OdfVw6296Vn0wjbfhtlJqXRTiFIGoXoswzZSxOHp3Ch/PSAjrZi/cVoGpHUpvzG8z
I5VtMgQ+CCbmGwLV84vbxVIH8/KOyXoVhaCs2w//nWlCQy8P3s38A2PV2lzZyMRI8rZ2z4WYjGqz
ISx9z7MamOYlbJHQ0WDPNUzg9BJsCb9sDH5PGE4VZsV/8LdDeq7kl0oLdn4c6XiPMX1EH195fnDg
HwNAc9Jo4fnqC+lMjm7n3RhpVlIxg0I2NJeFHXo7vG56WddZLvAHa2hvFPBwZpabKsikm5IObWjN
o5SzP82V6k5Tg/I6Bb9BBq7DgikIC8FJIqMCT/xl/XeXakZyDTZ9757BeqkgRkp5sADf9iMP67D8
8zAeoTVgxGTgw0z1qhO+s6wGy4annHIrcm5EfxnnU3PiosrYxS3/bLnnSc4WJZBgwyZ3MLfHx/RK
FTj4NjOoJWcupn/2ylHC8C+6SR7o2y0oDBEub0KQe9J6cOph4FJ66aipbs34KJzzoUD1xeL0p7oV
PXngOslGbKkmVady/PJBJnTkaMMtLx6ejZlnUrxzEq/VAj0Lxct+l54Iq73L4wY/YVIX18oHx5PK
jl06rh5dc2lq8lpXCpP7RjYyBhNyfKp5Cus9nk+XpqwwRhqOdiGFcGYyMqllW3BXAwuyzFC+QZMj
hf0ZKYKsvW17Eat7Zg3Omo6N+VLGxTw+cTRYrUFYLnOQDr/29LGz5Xl+0WXxQs14+kDZbM7qPt4c
cICmc7tPYnOOBse8Gl5H1/Ufeb7GxilZTl1AGk+MtCKbaDvagcAaKQ6QRZo+ZChZOYZCtqVp4biO
JJV4EXDQrLsgrtzdaWmk0VBigPZhf4LTVM9VA2pW7eTI1DNsshkIApVJ7KMthBsXY1U/cCwzTBEH
XP80oVLVZG/oRoo9Igc1mkHYx0uGGhrNDfdn2R3K/HR0RQ75v99Vf6N3wOBL3TCc1jk1UBV0KWdA
o2sif/0aMpMEWkDKOjoZFQYMZKwYz9+4b+XFlBLefvxBfYVeeFVpyyshHpAKBB0S+5EumzqDrubC
7HPvvwxH9uXrDBNjFs6JjvEqoff7gocbmQpnuwS2R+SuMN2SnmP/uHv5IoCMHZ+Qnzn403zt3VUk
L4Qp4wEK3ubC9JNO08r+nTVnvCvfBwnh8ZdQ+HjItHGdU5a3jIYM6GoZeCPw34BsBa+2ItH1Z4qn
rOxqllEJoSdsqSvbgz/n+nFXUyETYTxBlKeaECrcT7CL2irt+z1w5SZWWuQppz3+ulm3Tko3oSkG
6LLq+P8ZpFUzu0+J2TwSahxu+CH6EJbJXowoXnkDNqo5IEU/z9Hbv048hyohSGJKc0LatJ8qNBzO
wkzTIa9rAk9jJW47Wj7Ao5IjhPNP35LoWH3BU3sMJRxLeYpW/JKJFgo/CWBw1dp4OVCdaZ/EH621
Xu8dF6hb9XhAdD7dt+1kPp1nes0iypoInA8kt37UkiRfcItzgpNvlU3nX6qO3Vse6T7n0jtR5nMr
PBpAMHTWMd0KLLVoAclmB1TM/krSrwUNlF1GHGiMncD+Yd7+gSFiFlA0q0S08s0GebfgD4F0ptOE
6ok/7BnZHDIZokyK44/NoNmK++HfmmuzOaPpiCHPet3PpyDARtJHFGRggR+HeZjzXDOvVjxlBES3
ZsAk0dXb4bCH37EHmsmNpaSrZjWY436MyfnGWwlCj8EklimxQ/sy+SHfV4Xp41POrz9TxmwZQizV
yPbiZAn1NfCzVffxV7CymOe7+sDPOebzpSoBnAusOhv+RjjjnOtZJKoIQgdt7SbMXrlxmlmWgPk5
nBPXLoywBdeTwUEp68NaKsZgnSoEAcJlSmzWWWEUHKc8ADFFj7bwUZzp5PVNRUM3iA649929omyu
p3N1sfOgAaw84QPkvqlEGy9aPhdBnIuTwMalXsAQwAe3Jno7R5wMcLl2mRPoq2dvv8t2CE4iYEpL
BLkf6NkZjPCbe9Pjhg2V27ZVDKllGTwrRStkPMl/K3Rmeuw9gojqCwup8RwDVH14fwQrrgsEusry
Zj62gxWP2ipLdnvXUF0ZOtoAFzhx94HgL908cE89ssngYZfJEHLVlBIlZN1wU9DhE8l8eXqHdl0D
oJAhwUTjuT+jrQspcE1qUgCyC4OOS9GZzDMVn61zspFtEsLiSP/+ZboORTCRzItSuU4h4exeqlzo
Tj8XNxVtAOHeAC7UjWAxI/J8/qT69nHOI67LZkug9VLjkzbfwBU/scU2NpsMKJ2peqXvbv+sWnWE
9zKib8cmt64d5L003066iu3uThpJ0ccg6poK7iEqhyh8OJ8X0MlEGYEDP12ZdmXnyaPqeA2cuwlg
D16L227xoi+G9I0G15Zc6J4HNDvW50gT4eYR2rVOSCzPFZArtN//AGymqes5GaA2lBBQd6bFtCC4
1+tCG29z6Lie3aVfr4i5rYCGF970RAvpUEe72REuDyYPS03Xzs6b85CkPxtJDP3JCHDjCgS0GGyx
8/iZcmuK2wk3/86KS2rnK4MUGQQusW/42GoROrbpGq0my0LorQUnIhYNdNnvOjS7bcR+1BQFz9xf
Vb6DkW1ImxKj5XtuIfKOIUVVbfg6YSrWc7I6Nb7lg04u2ueiptn4R0TanIL5xpO8y5WqBIZk8Ohd
zt0B7dWgECN6mYP0wjFPyQxjOEvKP8cMK2ZCy3wS9lyXEhct2QqfuRi32ad0BNIMiszErug6GC5n
WOJuwLn58ZL4FEk6lLUXFJYgvvOH7+ba/RrkQJGoH64R5kg8TrwYyRq3B90Oxp2xuZNkNMdmIubA
L1cy6N+fe79dH2M5M46+YpS1v4vE+ZoG75d5CHapV5Wo4ryc9Cu+1PSCnbk8vR0xqY2gdJSWoGEN
WX81MjnO1F2bkSdrEo3Is9BQLS9Pd2H31ekmNQjvt3tI7kaxcLUmNOon3SpCAjyZQE3rO1rPEen5
XF5gtd9W9mgyofastln/0gXtWsp+7EWFo1q97kxmNOjGxd/1mmAmYLOJ5cbHiA52adiEiwAoZzUW
7ykb06LUfedFw/WIdG8ELmJWm0qCVeyvlWJwUYO3AvIZxOlT7AD91odI583S4QpWZUC1iC2mzU3u
twnJrZjin7SkmYyLBkEVJSbIZzYv1rufnyupLHXCuJlbA8+tBcLOQKftrt1OCbvQoxN4eylvf6sF
8GPd1XZZUGhec+TwZ4aFh8UafD02LKCO5Yf2BBdo0GG+ROyCtXGZL8JOoKcBeQwpgzI+532hNOpZ
9R10J3PcxWmutQCkE7WxEwXO/xX9U2NFmZe3OOhmeUZ312e53oavpQ3P/46mE3zt5SGmHFSacZa+
q8nutBit/IjfCW/VmbrKTBGGIBewRlxMG1xbz/xNUB6jgjQ2XtLdFr20T31KUSU8jBjGcwUv3CsZ
tMVWj05gL29qFVWnIe7uC1ku7mPMpFzynPzmz20knZobAUzmXIqzNI9YGfdLngHhGdTLCRjNsCxM
ozv2o23vNEYx4B9mILbv4A917QfjvHFBSLxyi2clHE9q8LMXa04IdvZnhmUuDUMVAaeru4Q72Dh/
s4FZemtfCA4Ok+NbElAgcdw+DvK6XSoLbyUd2xkO+q9KdWOsk6u9VvZ6l7ad/wUfNjFYjzIxFqSd
BXrdWntCz8zbzJJ+PU3RkcPlhO5HHTeGCGFwlRRmP1gSdUOsUUS96t55JYMXp135uAt0nSfo+Kco
3fzZJomXoCHHqIRDJWrOwX41zBE/lV7tEZBgvCfrHGrqjTqhNggFEJ367AGyY5kA+XK70DmVcco1
d96K6o5jSeZ0Y7JNqgLPKygAyhBzR4UCu+0PNoJ4LqMbBcg9wucMqWT5yjuIP8/7/cAmOJW555Qa
I/F5ixpiMHw30HymGH1xPpABjYa2naSCloPt1SUMuupCvS6Up6oYZGXnlN3nwS/HjMEJz7HNsgvK
vyNjn36YJZdHcnnlf0gafB1QcTm8WKkptGXIpN1UwiMhF22xjUB6B0oY2r6OHXOPK5Tx3osnyQuz
07mQQ3teY8plC80Ez5wO5jy0KTEe72oAWR7DQkO+Jvf9vzr1s7F347p1jDc8zFr1miZbzKSwoLHc
+ERyJBjEmJYHS4iKfCJ2sQ4scKBxoyNvKYQk7SnadWiTicFbFL1fHmUWMRp3jV2SrEc4VUx0RtjP
zWu/MkDAqpwJW9HHqq91hSn4F8lOvJv7k3bLpnutO/lSa2dkiuwXGr9heNPbxHpA5u/QwA1G6YYJ
EpIzXi247O7C1TEIuQQ6dqW/EUP8kjeoN3iL5uROmh42ukPvFnoIRC2Y6fMYrezKdMcwggz55JR9
KFZj5aPaa1/HXQ4750ojTYT4auy3q1t0NDsDoZkw+7foefzkBB5j7qCJO+wTpIxKDHSOK8tulZVQ
gs9MkKLYYfgW/PqKlOb4kmlya1pSXc7/Hw2AZorJGtav9o3wTbA0ca5LFyWYynTUFZG0mzHBqIEd
CPDfZxV+a0IJRkpH3wVZAJrN2DVCJyfOJ/G81Lgf86DCUG5XS6kJTucbNBObSRdbsOdm6GmYrmNZ
idGrdmY4RvyA3k1FI9jxT8veeT/ui7+k2btfMwpNJ554bInO0IJFK4syEFmPS1fnygvHumlKiJRf
lVVh9f4ZXozKYCGtIV6p5qnLXMSYjh3gTscNWZbx8F382AJJG0ekxzTx7LfxyZIkHqASjlGeO0X2
Rpv39FTYxIfYxJW4/JHiI02EMDHzEgMHfXogiduIOJbcKwMJSN3WK0jAuEK+yPFQYGyruFz/rCt4
SYhaza4xVdufCVZtKCs6p1l2t2K/8xeVRK5SlQWVonmZoeXv++O7zV8Vk5QUATk6yITY3WtqXsCr
jN9C6ScW67dt1eDJAhMZw86u1qiDjbKm1XY9yhwe0Cw8eUWfK4PPWbPTDZBQzAokEdyN3YBiGYaL
N98MGh6nZyxMVVMu5SU5zs+K2+scQFRn3k+4S0ylQEe+eP3GQF8+RjFIqSpF/T/gZNA/DrPn+5dO
L4+Kqmcq5uc73bX8KPJdlLyYROrvIYOO73LFdB+KmBSymFZWJfVnSvcRMSnT/LjYfXkYZ/TiTpUT
Sc3D8MKDD6nUUijgd7Upr1Z1wzPME2YrcqCIocO6srCua79V+d9COr8//2hHXIjDBo7nwoGaU4zv
0cjXITcFlD+HRNJBcaVP/v1XdOSoEjQAd5k3t3DuaNjsmYl1mwscu4GYYGj0nMkDD7zfhODjMWUo
KFcQ55TNZws9ZaUKxjBqeMbLAMmGsQdTpTdoKmdkr326sP29W0RvCxg42KHzGrNLSHHNh6oxbZDr
NsBmtrwWsqtIhzwQGvrJqKjNUKKhi+qOAfAPQruJwj95R6G4siYYdzfnWyrun0oK0xkA6ToILs6T
hgGesd9Pd48bT/RqIbB4l/qp2E2bDSSe03gxjdBdne9fHXaH3lcxhuZN+x8xKZdHgOvwZjufo9q2
NH4x2ZHs0HrxdEoPQJ1mCQD5e3CfYHIPlzVmPIY8KCZC8dzLfT97PXORNRw5zW7wuDOozert1nGR
2YSM/xhLcc/SSbgO9T84V1rfk6SVngCvioIE7OP1dZ8s4uRrF77vN1p/8i7VsXrpZn+3WaOJ6Xvv
J/h0Fqfr4kWsEaitCnwLURtxhxiSFhHl7+LIOU5PWMNt8UReQbI1mOVfphwSKvKDZjMlB2WrBqu8
Ho0CqfKAVtw6FOX4i6j4EElR2WHCkfAnmX/uPBkAqOs+gsClUqdSFlbafck7sZcF7bz6sHnals41
bt1QkVIUJbXuPa71XlQBjlJ5PT+i/2LZEzAOYhST96aI5LF38cND2w/ZoX1WSlmFMHjji4EZas8k
eE0I9rRtYjY6Ghhvc93J5aznUVlsGykTq6tVmM9jSww48LqplVK7smjNQpZG55CawJMa4NzExYYR
3bXzolGCxkAtAGxiBCBUg+uVs+ZoSo+t8Gljd31iMLNQ85FRGeLmFCV85LeSWswiI4y2hF51f/St
XKMsFdHvmk+k6i4VPZEENA8w2H6St1MsT/BSZ/MyYVaj+iTXO3nDU+StkcehgMGUHyGL1Vfj1Igs
hDHWMxgxD7zDySeC+uP7icwAsP3jJfO5T40niKOKYpxwGskT0pjqelIV3txOTWAu+/rrGEJ0yH59
FZB/B0NkDeZlmuh+iEwWuEc91drRpYG3Bd3k3GHtwEadz1/Y3N8Z6WUDOFPs9jv9sFzhAh/hZbZv
YQuzCOn99feSjhaGuG08Scvck02mg31lXbIl3ZqDE1b/gbsF57i6uPQpFCOvfM59MO2hGrA8qbJD
CtHcSxBVxQxOljIdcJeE6F/TAZC4CgYCBXen8vm7pagQ6R9sty5+T0hKPA2K5t+2hrpZsHu/ydjG
HoG9TYMxD7qMz4Ul8ICRyOKaCAfDTnvGtb7A7IWXdmWLQy8HoghGwAcGCBPGIBSPoLsalGwysI2/
4vt8jrnlciOhalE5GXmaQwYLvplNp7zMRbyU+kDgDvbimyLBRX+6brsZa6XWH24431QPBA4kk6Ro
Y5n0gpAxaNz5oZzDsZlrIFTBY4VE9baBm0EaXrnrGQrpuyZyHWSJ7L3J8j52eYSU9cHGUQr5MRfk
JSsqllPV3783cJgNF/7YRSjJRrOddsbbIb7GBNSSHNtKEf8fOnqFz+Umbli3tostsoLv8+WziGlE
VJHxcjco4C2lIqEAPPgU0o/aG2+QjAgtFK6kqUzCiLcamaZSl78tPrVrCWI4xGG7k1pRuR2QxwJi
JmV0pHE9qwJJ2yapg4+jrTBYVG86g+AOsdpxmCYJTksXiyUmG2AgWvU0f1DsnSXDZElK5yKx5Mi9
21wUE4Mvu1Pc4LI4z7bKaf3Ididt4Avx7jHgoQjIX2HTf/GrAGeRXDEEDLn5cExEfP39cxbTWFQa
LMNsuN7MYS5V0zR2LVNrpi7cJRKSUBGaeSXgnSaKupi6IC2u+cSq04Z42CaH+IM/34WP1jG+I82o
UUFzXlcrSDmEJNkIHWxBJCfC6qNW9qMPrj5fp2739powQ7sN58jaj1bhzM+8XvOslnfwjUtMVI17
WoyGSyFLXAfzmA4aRfq2fFU32ijnFpev4n9HWluXhMn8nBlX/BD/w3eyZSU2Xe2WU+9/keBZ2fML
odV/uEqj6BprOVEm8a+mq3uSKaMv0gaXlfTzXXaueW1h8WTnxV3Nv/4klYjdzL85TQfhYcHVnBX/
F+IWKZye6Tw4SexPeNXR1vfLbKpD9rewOljL28HVfDyvDEsOyvL18mQv+9Uc4aR8wnGZIwAq9qqb
UEAz9DFdlLblTBFY6P9yXCXR0tjRsyCAZ3Z9L+71jwVgI1KwpDDEVFWDaYEvw8Qk3hBHlanHgoWL
CumBt6fUjc1BO8aZPqvUu4xhWzYrr/UXlN7N8B7Hn7bhB+KRLxojcTncaBxQZtNxTLadCibonb5g
57xG9WGVcb+xejM/vCf5mU1z6B9rVZZudxU5MW9Vf6+2M8oJNUOsWYy9zkdz7YoLjJodEJp8ySFq
Ea+uRjdOlMQm9Ao36OFaCWAYy4gQEuq1omgg2nix5VM8sSw0vxdeai7LcWc0bMOqfxgJxiF9LPZ9
Wbxp9QDrsAzvule5OlVaLBZMxS956uCctxxg1sEg6Q1NGWKJxoi3T4XNwkz3ICy6fwL3rL97z3ny
O5B0+TFpdQCalAYMeWd78rf9xRYBSlBdGYa/ka2xKwPS80BoQjVLqgF6MgjOZLyZtlQodrdcvhBV
WhbX8hzdQhgDG592zVi6m2HhofLwbw5BlBkz3akhojO9/9GwhIcLg3vi40pjvgrelGzTEPEsm1Ps
S56KtoEDM/t67lopYbd2uBpdMSPgdDFOQtplCSxOuSCOEZCjizPrCklfs3bqRok/5XhC7HKKtL/V
Fl4LcO5ZeYyrmZuJLh0H3T5eXfH2qm1C7GlpJnIv8iASbatxn0L5Fg0jJzFqQp7SQt5Re5ZolJMf
yCDTnnLYEiiQ8hEnYQcvlOHSv4uCrqnW27oenkID5JUxmfeKdPj1BWpF24M6WONiDOaKenDccBv5
sLu8ORRBdsr5mrMnNnqfT6evP47DmZUmP6WMRJyqQCMrcaQnXjUp6xV/FVLn1vAnpWdPPGuYfrvd
v9fownMbcpMoSqKu83YqgkeXOKZNei8zMkf/sOujIoqUs4x7hEOdjDetEWBR5JATrypTAOdK60k6
+27qIxmXf9mnOuHEOWSJ/IPLSELT9J18vephhWYXsYmVk3HqEgIU+s5lYMtJ+le1P6xgDl39Euh2
Xx80zj0PJY7Jj7PNbYV0si5OS9PZe9BfPIeqlEgiHYxIybMdrpRqLffDGozVxve5DdKLqvsWgq7T
YaH2+Er8ItEv2dFNT8ls4ehhT2RGPM+OuqT1yvysH4At3o5yoZuDQtUjH9VEy5UtBo3Di4Jwf3wy
puN3W5TSW0AHiDtN0CA2SIFW+V6ycyrle2+fuYfTCGPjET2RzHZ7CMcHc2aPpAtc21Zq/cktSra5
tRxJj2Fb3x1rCj8SdwDxYA1oYB6QbeptWLZLmFyM5wkELI69IdOtpIQW2up2CSEBs7EW30nMa/Al
k7R5zmL67AWrVrNqCPGOE1NYsb0618Tj1VyeMULncJ8y2tUpZRLdMuOWIapMPcQ/UYdDosu/Qnj7
E+4nGbbnsWFVM1NKAdwCGYY5x1pog61/ea/Bp2656Il4MGf/44bGsfzdb3rt+6wY1yLL5k2G/YpZ
a0Gw1vu4NRSS+B7ZtUAu/I3azc+dQhTS1aNl3Khfx70tMrZnzX1GMA86X90ES+VGm8j/apMY0TKg
fETEWhzc43KR0b4H8A/4Y0mxy+oRte0euXA5arhLwrAulB5ofDs1bgxlMBeyqFThpsz/r4PojIdk
01a5QKFzNOMcDWXU/DMufYw2MBYX7/8/hqYQpcDR1foDbjZYwZe8eg3lzjyf4kA8FTr/JvHYV9Wh
ue5hclmKC9yTWvSfZ3lvwPKRMWUZVzaj9U+9ApGxnQ4Nj6b0Q1pwSB3WQcSUIjcgTJFKJjvLGpKW
s9xSnuVu3YebJw68qbcImyZ+V0yRBZtph/gIUBXebZxOrNID9mvsdkrF5vT6ihXW6rpxubOoLofP
UyCwYcjDYHaw18ckvc6bK9M0opPYkSNHs9AQldz41Ee08aXPPvGGevZganXrJoPEFqXbuIxcjLhB
zxe0EIfDxQj7QTN9kaX/tKXivwrn1oKh5lR1iK8GAJ3oaXjQd0aQr/cNih64migIpUuqQm4LdyTX
nmbzCpQPSP5dWArvSa95vBfsw8pe3YQAO8OuKbVp3gFFxr50Q+TH4jh4EwKI69KszjUyTlWftEyX
9qhKhNWaGK+0E6S1EL+cm1Z5U7/hQgD0fOFcVKuyKQMdmE+vAZu5NI4YWEmOx8G6eUdu3+1XI4LU
o0UeGAxpWBdWO86z5wHT3T1S58nmAKKybj4hWP7BnFiC7jL+1lTBuRz5hzBhNAJfLqg7mCewU++O
P7w1TiYSxa+TgUQISyaA8e49+NDusXPk33ZwHnRaGH2kMAhCxMoIOm9CMguU4Rs1tfw4dns+Sd6U
3Lw1TZPb0ca0L2rYtjAvLn0GnBkC+VdtNQqVjZg+4ObFzFQoh2Xu98iyuRBiPQh/SKsbhS9IWgrQ
J6OdeqDPoNKpCK3Ow3cmR/mSLGkCJrT/PzqwMV/B+c6nX4JZKMGKuNXNXnty6awNbncd0bHBWzNM
1B++NWDWr8EZTzVaMatE02yIncEXbfpdzTtLj9E9NtpazY8yjUr+IKWxPzjNTT817JxjKpz3G5Hm
TPJkBzEpPr+UDK9sNfpzSIMD8xGO7lVXG8IK24SYR1x3Ni5ryV/QKSzoV4es7+Io3OA6M8oTuF6H
X596yybgZtU/8fFg6zO7A6wyTUr5lOClVWsu8/PQBcLFZF6cEq0jp94RvEwLWzdMa7AIOZJtiYuw
OihxscZCBSJysgPWkffGyAzVcHoQ1DznS5PwUsm4/NXfMAsCejh9qXmP/dLweGzq67hRkLnh2vIl
DMA2R/lkXSpj/v8wjXqF99aZjO/MCXNOeVqr0//5WoWq1jtToAdXecUmOTAw+k7O0xDMosS63QF8
4X4MJqCWxyehDPK+llT1Zaj+MItSbqrAbGqCepEfhs9ByRLTsNk/jovWo58WB1e15RwrC54X0FUo
dFyTkAVEWl7OOLtm6cTCNyP7jcS8StRML9k3rPJL4IWJMPQXMuuD2OL4NdB613FcnTx8HYEvuCQ/
ghA4vju5u8BZJab+BIn3OwCm6pLOqswEYYLImWIXmbtk69aZPX/EnJzWyoZLvmfG76Mc3HEGbXLN
MqJpmABi6KcX5gwEDYyGu+hnE0xZbyPRaXwfnI5Yw8DlodcX3HqCcUJzQI4FqoEsGt76eW1Dv954
Ovp6Oi8PLHG25XzXffwOkxsomDVS3qJ2iQGdUm45mCD1EHr7kQG3JxcdgxcJA8xW+EXuhSWofCQy
XvruNXftOQk6EI7EjqhcY7EowHwJJp6yzjDaxkhcJ6CO1XdYM6aVz45Ex7JUFlW7MJKvnf6acpdc
9iPWmkEZkE9R83wLjFSDSB0Lh2y3ecxW6M7mqGDBeHw/c9Q5+lGDsmwyH7saWMh45Xe4LGJPSs2w
9GXBCJ3LJYd3kl4QU8JCQ0972F2tpRimb9T1WkZHdHq2dytKX22dOv1S7dTnobI7RmBc5bJIPO1b
bAAF0UaNFT00P2cLVU3cx0HvgSSEEdR+Cj09S+u6wW1SGFi1sbE3FSQkJuuSEhSXWIk3Wfcte+5B
i1zvcQy/g0nq1VKB9z9zMe3PRYo2uqX6CbTnwk+19RESE/GoWuDscZBa+QX5YXs1Z3slApL7be7m
SJNYJBrZdYFmEBClSpvSVzRLRZxTG1rF0iwLFS8+9igWF/3a0bf+uMdCgOYQ8vFE0OmNra0LyXuJ
ZJH1d36A34ms77rXY2CFTnfYWmHqnhEzxsj/AzwvY0amzaQEAEXDJFZblAz747PkJKGf3mVBlh0v
j80gpQQFC3YwiCQJNDYOSIImfaWKv2a6m2rWylrxn6B1PIsnScAjRUcnXyr5ERd+pIVD6fO5xCOq
7fEItpaJvyqQFsTmLQJLapl8HOGmpy8WUyJDP4jIpIWNCLD7aqEoaJ05f7CTp/RmxHjtyyIy6bUQ
9tJQ6XcBYXx0Y4Fx83zz8wJ5tNlUmpPoXkllmm1ypdOMy9CD8VlFlGMDTYzuBMcAME2CfDV0VEAb
tpU2rLF3RItQ86BsS7glwIfeRXvlmV/S/6VMEC/4GgId+c0Iphx6iehQsrDNVJdE/HCS9yAvJzTt
vu7oIy+I1/GrNXq8feASC9rC2tEkQ3fRPzOqcQN5HzI47UHmvoowlwakRMQKZN3uoQp3JmMHcs2W
g3lo2dNnRF6OLOY1sajVP/deGUWARLPkts/t6Lq5advpFfRA1bjtarD2xpWODuzeMH+6DxYl9994
VUwF4kDQ8QrxSiEErPeQpmHdViPKw1GsnFxbCgUYYed3pgrqTbEt8U6C5woJySgRekL+w3gvmWpn
xJ85YnRpoNr6YCIObxip5hrqH/WTHba4qk/F+11nhJyJqLJl3AtVtBF5ogxwGIHjvZ3JqJbZiZaZ
lpgjFJxL2hVrJfZFSAtimzTL+jSAXDT3UO3BmlmNjnk55LqF/BLLvlLP/kDD/JYf/Cm4yGgSM4jD
Q8N6NwBuCYeL6znOgExchOf3dt6IirBV3+pRuCoAQVjY2HNlXGQEiWFQrjciqR2wgg6O/6tB2da+
Mg+eTB+OLgzsu9O7JkomzP0JW0nidRzvP3RiOYQDItAqaqm5wnSSl1pj7tNqyfyv0o/qeeHYA1GX
NdzdJtop3wDJs2MbwWE9cSrvI9kV2mZLH93TT8QYNuxYNpGH1YtvcIR7Qs4WMK8sR6tbAxr3vU6N
cqGByCPo2o7kac/v+6596t8+ejS6fPlLazfOzCJrmL4HEjsIV8jjSFdiyamxfk/A/IPYQfRWqinV
corscLW2YfvaptzQ99El/DNwGL/0+RTVONSoaBrP3RmuqSMYhyVrnUu6Z0lwmHaa9WzctGwiGd60
ABd+uK2OwK+Kc9Mg6YgIexXIAbkRFnhEhKjdW9hGWiLYh9KUnXocO20yJfqOa4bptNOpIkBWD9DP
iomL6noF9bACoyVAh+FAQCWfIx70vM0yLuuqM11CT5Hh5lwwgCSy93i6yi85NNHRIRext86nzGpT
/jeXkYLtV14ex4wxkLDVO2qxh36jBGAT0NSQIA5FZfZA6BeTClDCI1/7fk1ba4cp9rkzrjDnb56m
BoSADRrKUSEDkSR9RTzEwJKHVT9PoW8FSaMuUUHTjgKk98w9mLTfEP4EAG3QjNPGE87dlORe9+xB
iHbOINQT+n6WAuSTY3Bt1RpD1e1KhKsxwJeEXHKipjaHCRyywcqmGQ2zjN48VgiCsrPK/VOetrw4
Z/yP9iqqRwZZ0C8Q59gL7EDqjI+s2Z0hiYtTNeKxhK3t34gDnKztIGpx8Vj3i2TrKhrIeK4b/NfZ
eUA7C6SEvrAa/P/1E/nt+hLte0vqivNM4NF6LRZ+vE+1UvX2s9r84sCgyPx9ziRwUvVegxdcTBlv
wglPgURujxrIgLcecVnVa5+Dw+tYRCHhVW6prMAepyzTDQ6HWD8P+ktP/OKK/9sxZUyHfZcYTKEw
Ff2V5ay1gUUCgKe0DaRfB2j6L2AWdlqUdOL6AUHLhzRnlVG3SfwMvoVTOVZvrr/3gvyIWrDGn5qv
g/Vp5cWKx5c4qPkdHiLaGbRokGLOiIYTnvAbU5U7Nk1rSLbd/xEt8rTlRKL1zlfU6kUKSgGNJm7h
+JLq1yVDq8yA6jtq3hBlB/phVZT2QXcl8L4iXoV4sDEjnBho4eomVSR72tFS5O64mKoQDvY/qAvM
N2r2QlS4wj346vSdYnlngG799e8SEpFuw7+Xy5F8r0OXbWlOBszWt14CfnM1vAQAYvpAzbzzTKQz
z1ga8+vH1Ggn8TQxKvPO1nP8Q3Kt4X00uYi1X24psjKMLJMT1roPTdo9VX2ksBB+mQHkKfN+rKRL
yrkjGAvkBoOZt7dib3AoNylbWlbItSfxfKVc9a1KB/KyOWvPM4TZ3e5dgnCi7flS8k84u1RIirGj
u7Wvqv3qYPmJYWplWLK9cHC/s4+Nptb7CE67P6Uo3xZ6y1PPZSMyWq8IKuyFJweGwGtcCATa5jBq
sGCr8IdwlYje9YHJy3kBhJPzvN+djO2a1z9AIuI/yf2ztdOmiMQQFZTIgGPftqh+3ymCHBSOAZOr
eOgM1VvOyIdWI6PkiMHgaAHDfcEuMQPRByZnaTiRydcUPeVVMrxfrx7/I36/tOdeLYhlMfaXagqH
hrNfcilyb3q1I/dia8ZGJSqKGe16QW89npnTgl2bFLeliOXHgYijfa+ZiEcs4LsqFrUB2QWiBuGF
qveYUCgG+u3tzXTHEE9SLXu848FSIqvx4KL4TAnkhp628nUHuMbnR69X3eeGq/+lXWNxdItzs+VJ
S1KyDcrtBa6Z+mUI0c62cvH0NPDJ3xJYK+B4/MrUoMxYsvTngJ43JVYMvYpBMfUvfkzb6mcZ8AC1
PIQ0JVhEaQMnx7z1dlaSCXxdWeKNwssKm3mN3iaJK3t9BSz0Xz+RDEi+Opm2YAAk3u1/Qs3oAoZO
8/V2W8H/d6niSoSwiWsX3Plpll3vm50NgFGZOjrv/eLCBA78ZAHXciJI6QxPfKi7ryKKCLdvK4/Y
lAz5R20pv3e4p+g38foE3nl3hc5vh40oIDG5TFC9witHJmLCVkLXWkWHg0DnQEjlVBcgVlV+B7/4
jEDfIAzNfElFCLW5AB0K06FrWSxPNVhh24MIugOg2yLr6zvAXxSXGELrxSAeLt5Y7Bzo7yJQ6WiJ
bY1PrtTMuvOYQrs9scGJeChiFUrfz93Y2+fJGoXFwY3Hui9/tnZPLUGiZ0gfmKh3UPR8WcrFDalo
qJLFLZ/t3NL8+LzH2VDiHHyNDnoaT+hpIQ5GcDuDk+CTfsRo5+lxbLCI6KNryqD7unXTVY04WP9f
6Ly/JbNX1wK3lLTSxcilpCcJ7l8QSPAWTu0YhXcnKtApz1mB83eZ59BPUTzxI1uej4qGWD49v+5D
Fax72rMDdDDtr5xHzO6htzAcrp2WtD8Hj63yZjHEzVL09sgzzbtDnKDSNibr85XFKnfSUO7NXZvv
DmrSiklVvQWYXa+0YpyYVHmsDYG5chZMHLWUxqeV4ahXIYrJQibZXFV4NOVtZAov0d4rTO7J/kTa
5iVjzZx5rA7puJHK2UxEqmnr4mSBdoQdvEjfELGuabCTu1lbTD3bR4AQd3DfjWDDh9fGD5E+ux5e
JZuxcVkDBVwH4HQ/rCLinTPwzR49to4OegY3wV+b9lfElf2vjU6ZGjrnbW9rnyc8yJOyZ/LCuOoK
6/VSE7B5KUaJPKYwLpdnKJi9qrl8n1eOxMo8sHE2lakfdIXCTWAEAiWQWN97ogbizkbh9BKWJ/CP
FH1Rbxc322mOEQmeEyScI7P45BrqLzV+S4wMhdie9tKlfEt3EtpWqhExHCCd6+z37+uI9DEFM2av
LYWspsxV7yV+h0u4Wizmt94ARPfvGNcx0DmkzApIu5yv1s3Dfy8F0ZBo3TPolICjytlcQcgg0nCf
AG7iTUyssdp+8UW8tE6TUXu5z/iIBn6t07uQ2CpmesSwK+jQwr/ZmTCmlv5bs10PH58eruOwu2yh
TalHrBGP4KZx5PiLlsRL7r8JeLolWh3dijc22HcBTmnwnJoQYMo96cmRPSj7SDrDaNVIQA75zCIJ
iufMQ/sqBgIPYxY/VUFypPO5okFfQGyKezo4Ko3K643pB04QuBZLBn/wdTq/Yo5bF6etmNulRMLl
JVXPWwIp2+LrD1IbbXDpdvMsphkEW8/1oQR5/M2gKbVsthEAXF9u7BbNv336NYTlmLf9WmtYCjMg
oGvZTje4y27HbgQd/oCpsJH+glXXHK3lzdbkkpOIABJc7GnqtjLGg8DS7XeDhJIbKfE7nKPeC3Wm
Uavm8Qp++M0iTf8QyTqk8Q4bf5hiaczgMJgMEJWLP8hBfIEsqouPGeSXTGE61LciKHtK7CgggrPt
ds99wfeJGYH7RHsuw53Z/EM54LizBLWthKQpZJU+Z9zBt3MgkLx02IY4JVvS7YE5G/l1Cnx0zThZ
x4UdqFpevsJn2tbfFBe2XS/y9Yyulsqyg97nG/mx0c5KMfwCqFrpxT2cmlyv67+yG4Kezq0rbhbC
cBsUaPIha8q9sYN8aRiYlUYZC/xDauRnx9tCD+GJ34+qBQ7p6cKNBPGG7bDbcXI8vryfQF211NRB
H/D8hZefaxSS6+v/yIDwkspznxPEFx+hQGvNpZa98u0DJ3dAMvPLynPFYxvZe+unx9QZ/KveS8u5
anlhns9LpX9p0zjDS8B1p4XKd9RFRwX3jo+Foc/E6yDTn6bWJxDdf+O1j9d3USizgTd5CkB9Ynk1
wvVO/065jKtqwcKT3+lt8nemrJofue/0gFMogC0dGmJ9dcaK0OTL5ZLjGQzVIiETwaaJON8cm/vE
DN2xmT2Rmpl+Y4phUe00EyKdlE6n4wvQ5h3N34rx1xy7wry6/bWqAasaKRseDcgrKPdOl1sYd4ql
rmle2f2swG96WYeyZA8nJWUoBd47mDFVVumPjqsPToowj3O9+pHirLnYmbaw58WonN/5WlTSdu/w
Rx+VKuM5jfjK4Ug6SQ/VKTvr/3zNsytEvxBoLLtEJymJekrL6Ybb8bQ+lUZ0k/4v3uP/zZMhZvl/
CDEcUv0DET/kSAKHJB9V/NnXv2LbdKxO2O5JQP1TBa3xZx3MYMRzJ2jQm6zf+xr24O1YcTmTy98H
wvd36mZztljHEyc6ZU34LK+sji2lWiSUouP2Rhz8zswl/errj4yK+I6ZjkMC8bQpw6hn74iirMVV
DIej3C51oEZ7dj4WOg/rr9rfHaUwXazUw41u4SL75POWhHDmSWvsYn32ktYUecFGfL4AC+hxudT8
fhx7cHyH5eve7Z4YPpzblVVum6S51fhXP7jdAWeN+PCohJEleOOnOSxszMDwxi9pv/AVPK5kw3IQ
QwsBEeQi/gIogCkAjHQ3hk/nd5LUd2N1z9ejvrR/RVi04g5W4WyCGOKpCkzdBN2kfLRTjYUytvoJ
N0ZHbtykQmZOE3isSz2+BQjgD2mPBmLuQvVmWi9iVk1GLYF9KVcwi9JTiES7+QmHYxUgGiCujUad
G5XkHDs/7am+1o94JAknnaiRR6AlH09/D4ltI4wY2AU+A8/6wjsq1PqZHwjvh4Yu9UOO7JMyBuZ4
rM+SnnqAsudH9h9Ca6wD4xxdE53TrP+ms+MaF0QJvfnz0GxcjMK+e3mSLvkNNAoKtmfIieeVG+7n
XsIm4+mF3UUE6yZnZ/DYwCWwjy52OLThZDL1/O1TWReCV1Dh/gl7E2gqAWe29UUCJ3ax1XGliMBQ
idcx3HQIA+kLYOQxWKk5+J9Xgt1/g01ZueH6s+4GWZr+ygpoMYxRXYuy5A4by2RY/GjKaicWxNHg
TKSoXQzUqFoqcEtOqDQ9H0qhwrZf2zKQYd5FKFqIVc7e0kLSzyyhtxA2YAfAWzRyYuXQ5LIUb8uI
IHPEP3Xh4gG7jqS6WmdCWN4DOQtYqvgrDhaN1r7Aud7UFNhb0lyAtnjwKDC970P7lAV7nZe5s6Ly
PxrmsTz2OTm5RwbcF74FbrHGciWYBm2xwIgYaClOg912rO6WBIZNjoaFALPzwyplmyty11XGxUMi
yoa3ovXSN0/0YvuIw193qQ1nQkHpS0VaAndKfy7aczBT9t2HEVyo4L7ZPHAEOTI5j+zS/e70+Qbk
MXzVpVS8vq8SSbSbMtQlfmw6YIP29vfV1e8ZW9PwE4cvySNOLA6NbcAfOkDrephw26P97cqpHxcs
jgrGbp+xT0RKykK1HyyPhPWEvoSJQwkxd3emZjbjoWZzvTIzZDf0H0qV8jKjdYp9DV5IQKy9ujXD
jjHs+fH1NMNd2Vmxi7npQ6DZ04KgkqjZ/IJYZnQubXXyzbKytVSKlqt7Htqsc8/WPUp4pF58Ltub
TXwvl+k3UgKu51Mnp3if+hY9IUd5bB7JXjKW08fIlkgS5niaOHfl6PDIjWWvF0BMSyCskaFQwbXN
UDg5iwHNtnA4BHHuxxU3tvYwLF6SZk38T/DAGVIhq+QrIo/9sOj8Lp9j+y/4Sw5vqATrAXvbxBo9
3ffADqFwki6CWKDwe71dl/XaaVgxPM9iYPK2mtgkZCgQmejqc7F9wzoVvG+qw/j+abPDwQOcHWIr
yBMf+SeApmzQAKZ/ULQ4dzBYSn+OmicqLP3HJED1f9C7F9DlmAXq0ZYJ+y/izzKNUEL/TvjV22GR
jAbgjOuibxA7vBi0qX/W6t0GFIH+aWlGwBHl8S2fD5tfOWvIdJvKR9Vx37wHNjsAiGOMoUdV3zms
NjUJfd2UfKoGj/3jzZGJPPkMp2Og+2cWkwAfAIioM+Sxmp+abFLUGq+qIjIDydJek53+9WSK4UWc
ZoDw2FpgIsoy/+x3fp7twt4bsI8wTcR7qXrm4DpWnN4zhHFXbKH4VH7IP24tyUeRf9jARZ9ac9LQ
3IAH9Sq5xJducZMbuyuddXZWNSdmoTlCof67AfjbNjkbXm7BdAUu8rUoaWQc4LxKb0WmTV749ZxQ
/0F3BEuVtfuRCjEErrgjT2iudaZM3BEzLjG2KsCmrJQfK0qNg811xR2QhzCGG73Xpu7+O3/S4/ht
GCLYelw69fQnnLXoFhQxdO87hKQi9j+iopBX7u/bZyqaBRpNhqhLslQWvjMUeOlFaAWaZ5W0wLA+
4CMN4GS1Z+qSe7VgrYl6NX/qngOX0LAa6Hajrorv1xxooDKRtv+uBK5P6pSXZmE15HO6jP9/rsg8
zlsnOLBQ9rfYTOcTEs1z4g+mceRST80j4viSX1b+gIeYhjTtOt3qcU7sRODjqeFbxVDfK/QPSmdn
f0Gq7eJtra8xcg4gBFLjA1fxNGAx5P1pHuJNf+TVjTo2CmH7MmRijWvvTXS5xRtEo2jfBFauAk3s
jwC1vUJiw8pre5mU1VjfSTe/kRkw38SJ4n8yc/vLyZ9uraRL6ln4k7M0gYoylKQD5f+1Fwn3UN5l
2cEoVR2C1OoDycAcTAtm/qzaVWxTZDbplin20rkBBUMm9FKw8rmL9g9D6Fzbxg94NUMUqT/k6dY8
zEJah6C11Ury5uU+0Lh+xR/IcRChIakLSIood6CSZ7Poj0emq7mAWYy4lVrlBN7Kfd5p3Gh39QlF
huxDWUDDeOBr4GlIkIn8fiLxYVmfb5rYEX+dYaWcdZKrVGSUHLgaLiERdqA+OaieIyLVWaEscE1n
q8dLs5V2ICHt3ZsBVFRq6qiCiW3omOd+S1X1qH7/C8mYkecNVXLjr9n7XW9MypmPRToZIBz9rzCo
y3iElGemvK7xtHIfnwY03BfofxRtFb708nUcXFAUJD2AjUcHk5FLRfw3ZEeDo0QtUISoAXszyWBp
hmWQ0IN00UPzlkro2eJOAO1a3V405hEFGIgE05VwB5fRBf0N36G2nM1LlmaI2cZqQmMeEglE7V2U
/pX6VaGJ+8Y4c3TwSTfj+zMZwqg+BVMSCQsYHwSWIv4SqJBjj17PxQs+m4C87YBEgpWjEyUwJFmh
c+LCZfaC9ov/FgHBllP0hc0zZwlc22XOjtQXf9VrT7e+hTDrh5QcEr7BKFfThDfp/6RTmXdLWqeU
dWJ2q37qdn66w3DB77llTK7gq4glliKOi/gF4aMHAk8i6e+G+Zxiqxv5/O25Jbw7sHlqeE5xr0Iq
XgjX1bYAEtgecEFpq/l9MdsdF53p8zTwshxc7koLvbq1ItyMv3RxFhATFGHs2V5SMbyOVX4d8pv6
Akh3RNFaZxGuEfljjYFGPWHbbOQFV97EAgqnfIleFRoJegdm/FZTohs1skb9j8k2tTXzncjmbM9v
wVw/0iXOjw/LMpcdZuFYrQTHYAHNwdoxt0LamONQj3ddRgDz97QynvOpeJiPpumXjT0fcxU5wnl5
A1f8OGMfKcYT8Zz8DIUoTu36ePyke0pjdi9sSq1ttf43fjt5rsu9ONn5ep/VEQ7AKFm83yr43Yq4
IEh5bqRooQF60uVuNQ++coSiYDyh8hIPIX4sMUjfGortjit6CKOE5vaIwnbI8JB7YVnywLY/SO2S
srP2f9fWdvb7yYeQe1MJeDGFdEo6ng2l7qLUN2YKVzpADZFEtB9K5FFfxdKtbzeaYbAa7+w9Alnm
0eRhtyC+ZIcsODQYM30kUdt0d/Xi4Mby/u1wWNgqVabOfu6b0x4YwVGhtYVRNy4ezeaKRW5QzFbk
fBDR6e98+uSQZ0EWH0Nvng5C25CIyDRQAWhSjDvpcFWe0TqLdYFoMEC1cN9EzGaSpFOiGJij+PQM
0jw9y7WDCt780Vk8O1o7GN+uSDfKtLLEERz3VqDYHqHu5ip07otCl2/qDwQiOeesgamZTvzwYAbR
XlCo1NyxAO7HWVRUHoKZZzM9W8iJ9HyOxSTgYlswLTgkclP4BqXI3b/B2RD4z5cCIIsKPOGv6rIM
wByoglh9KIkCsruaB88RI8Jec3VvoQxwPxEPnNYkdG9IMuKbpq6H0xpUCumHY0DBW3bd4pS/GlfK
9lQZosd6Fz7YOyyqrchrXFzQ539LX08IPLwLYi6CKSRp5MdgERMuC8AaVsu9SAq6JeyrAWnGshlM
FQIkTp2sEeEPSoG+i+yNZwWu6vJ6HsRL3r3fQWf7OEdE3TofvkD563rXpkeaPL5HtNPFLvRa+1ej
9B2GyYB06jb1wCNzcoHlh72eAzG2BRgMCa0U8mursXYZd3vH08T/FLD7Nl+LHnmBdm2FfG1ykXpu
SbV3pJXBfidnl9I8O6Bii0spFaagnhIqGwQSSUB2U16+m8Q7VqWPxklWXb3z6//Aj50iE24mJMoE
l89Wo47oIgNIae1mzEl6RfXWwabm6A9lg9rRC4SLiXaNiTYP3vF2hfnrrSqqj+az9uGyNc9z5aJS
/Cx9lwKBPTu2izQQp0GjXTup1BoD+bChl2ZTdtc+DKfD7TV2omCLuQ1UdJRS5dWbej6aVrKZKAuz
LxyAd6L8GHp8tRL7Emy7gipENUHZdgBzRpFWqPPpMR0oDvhgD6V6mJRxNfkz9gbCe4KZpKjLa2uF
Er4wg+uJazsT1J3rI3781RPB7wuBeHC3VPGj/fjKItPH9KTYhyG4iWXPwNY2J7GQYFmBlrVNL7sg
45TI1yCS4g/Ed9M9y/KXn6FsyXw9APZ8xx3Rf6Q/d6flim1OzRYEaLfgzmQxyA8oLpmNuc1xYc6t
Xm7GJ0Img50eVDpYp2asBZXmhnCELXoXgmQTPYMQURIfnaJ2Dugy5fNBruvxgtA/jePWrDuNj6pN
gLSJahqcpu3lDoeNtw4xSqJ9Xkg5IbTGeYk7LkK1p8nuaCj+w7R3J94ddHGglvgc51MpzE+tiVqM
xE6JaalR12XcClnCDrC5Y2FK0LyKg9soLBBNrj0tRRzce0R5FboziEQ+K2wqHHyMy27QTuYX27RS
RQaYojjceuxBp8TLZUziI/7ThTqTaALzcFWCr5WCfAnVaH+vPoAmNMjQdGK9kUowv0Bf3aW+HRlF
BryepQy1XBsQzaw1EUEQXEZMKOaNUlFEMtnzl4azgsdYDN6hEKg7WIlhJ7Sxf3C8IySVgTLzDQH7
U8NaeTMVZIzl7IPtI1BxxImuOrqMiDtN6o4ROAAxqiVhR3f/Ht69xMkq5bnRDMN3AT7QlgQmsTTX
9RwaNUbSKCFpqvHOEksX6s9FF2lFAK4s16yTXYet2Eem15oKVYhBmpA1phV962pvCAPth7FK86VB
DVBtVgxZ60bKuyBSFXpAYMcK0QHvOFcEbCQC4xu8mhlmnruF2TU8Y0FE1AJ4jl4TXjb++bi32RFH
xS17dd0BbbpcVsJ6DpdMGgOC3b7Uwen1tLRzG0706tXfUkAXC4ZCiitrSaWoELPGdn5Jh9wQo/7t
v4UFzWxeC+9p9eozjBQ/F5YDLJk6J43T7OrgzReub067YPr2ZCGQLIqdV4jLbPAkSjSsvx4iWQt/
lcPvScAt0I/ih1QI1suEwlLSJa0DyqPeOnuR3+GGrinb0TjeTtwLS+32WEp0wyTwCVEzmsdKuI0p
svQLpq9b3yw7wWTKjCou+D/CEt5mNWgvHZFkCi92yVm+8Udbn8db7bFXWVEduPyvSfeKNGmxj9T+
aZP3rv3SJT5XO4FyMcOuNqomY9LhU8GQVh4Jyxpv2jDYIusH4vqyRq+jJZDAhUMjbAHe46hMqqLJ
zIZjVSFiiVLoMzAdhzGep3zzu793MjxavvSAsjs4z48duLm7CcfLXH0IEkzLQ4T0PRGZHQJZbitn
xOUosE1expg/7TA7VEElPo7SSHmr4C/dVpKzRt6yaoxS36GCNGJATHD60AauQOXUWpyb2QppDwyH
uvjZzXb2cN1mv4uUWNNCmcd06DtxW2MttXm46Y+IKzUWT2aFndaejzGvPdvUOrnKg+Ax56nLAfHx
d92tI68SVM5WvdO1y+u9wJ5mS7JDY3k38/vysQ6q3r6SYy2mVLMZa9Ll3qxMOtgJvLOQAAjzjNEr
lecWS1i7zsx7JoSDaplsi3mprAL9Xa6SwF3BT/uvkUw2NiGlCOXwyNv5PjyN8qbdCWtD7ZtgwDed
tyYMpwU1TBOsvK3iDYsSFhF7IQq5puNmDxiD7o/fQOn36yiuvGh6MbTlLP6IG9WfnmeMY3hK2kpA
1Lr4Ya8AXckuJMgD30KRX9+qYvmspK4KOqB9GdR1rpBHBcPxTXlVRSlmxYg6A0qZNByPsFA3eebE
WLxcclSWcb8zaIJVWVpGdbVtPOik9y0A725K7TlgSYNL+cFR3Z5KWrXT0K5vVTm7AlJCy7e+cPhB
EtCjXlwswp1Ao0smOSNcYO0bz8qg1WcNYpwzJ3Os39t8ype3mxSVjsllOz6I/KWWPzoI3GzHzGPT
G+iyRfcZwmKB50Jhx+FjhLjH0S5ErZ9pmIa6lOyIl4JwVTxByaf2rj2wjRhR92c7awkX6XyQ9wqU
pYtLXyLpFTVq1BshJUuCecH6x1XR2MSFp5NCAvNzYXlTFQ6w4mtnzGNPhxp7Bihv+ZzkriLXZr+6
vhF0nGzfEuFnvzoHXlyMYBLWIsqON6NAV4+2EThi3z/AqAjmLyQ4TqBJqGSSy+cFBPsKkRgHdDQA
DddoYChdbuiPnCUWqs08yNlfj6yZA9dCRJqhdIuFCpmi3uEs+caSp6no8vbFapN78oOgtpdZsSZJ
Ts1I0C9mlUVST5860Qz4SnygqCD8Wj5yLFuDXsWWTx9kS3WXwk0/B74ai4B+rmFThVLU99VlzJLE
ZjUMJzTunXt9nrJ4sy6EaB4/9Nm5zKLqHCscD0GEi8SxDvMlvYLE1wP4ouoga3zJFT57N3ZbZPiy
yTVajxDIxN3S4smhQsY93kT0GctSs3LrIrR8cL8+BpFMPBWm0Qhw0PbuLL3SPtDiohWyUNR8Iv9V
qQlwTMPACvKkAaNlkPr7JKaUqN0Nmw7KH7N8YEE90HwnqSyNSi/jQ2ArlF0UN8S1EhFMaGChuUPl
vjzaVJ51kgG6/8awZUo0UgMrapm3gkyo/iQvM5ECYN62WQDhZgQk2LSoG3T5r5YuhIh+D48wCFEB
R5zgOff7sEJpY0uXSmZjD41oO/CfmO9dUKfcBRJuSNkHkgzZSzxM7RBoctRuvvtkxNny6pa32NsT
TbdRsnN3pQBEbEdjxSwj4fhDgcusaKHZwrZOzEB/jU1Q6FlmDALDvqaJJlFc+iVhhzt86006ask7
hFz3VKFAfZf3x2HDoULom/YsBMYlkSwPhaU6RgI2s5fsuBzNsIHZWZ49a+I0Ov3kAF/1p0h/YpTY
3SLrQpclKpjg1vOTFGbM9KJaHaPrhPNtkogXoozUV9d+5vBXfyOy8oC8oCrHZbgbkGLjpnoExOab
oLW/b9Daa11FiI88ujSJKrtxKXUtfLohDA/WHZasQwk2ualB0VgS3m/1d3S1abm+ZqGPH2YVc1Gt
koaaixhG7F4M4rZIXq7x/hwARIylz3crh0AZEKiC9Fr8BgGwK5OKvNJe4J5gAhWWFni7uGxtqy+R
tEosSvyN8+NMk1Yr8NPRoSnRBUGrpIX9pfO83vsKlivID/6mvdwlRDrtRbJyhmpeCvIUNLjhR1h8
9tN+ybwbskQoEr54/F4ENxothIzSRTspwxTrGvXrhQFahFLomvLzcOFJBFt1vEyro7RQ7ftTd8S8
mZPgyXYSWuTKmeWrglTkJS8KLviZKcASK31S5ydgoTFsxFgvUZMbbqMlp7Tf+Eap9eBb6ASSpICQ
u7zcdZEThkQ1Fb/h3wYhTRZCP+1rchuZSKm1CWb7KrO0FRgF6A+I+uFCbIrWH8U/WtefASpUX/r+
7djjhBxyVjEKk+0iqASxlxPZdhwA68UU2hQ+IhkF9shECNK9X/+GY63QH/hPH6X1ndtMkc/D6iuq
BeMAjhRFZQNzDyyt4wLB9VPKBUOZqlC019x9DWPIRMiAYryXsNTaATuyyRosP4/D9rR0gD+z8lA6
K6IlIhWEaASZQt6QBeFvlnVJqZHadMYAGA2PkFWQi7385D+UISA+ukfk6+p0nktvDG1Q64xS2u4l
BVyeo4hhIcO0Bw4bZhab/Pl727DWo/skpPIl6z7amVt7VkF8VigBvT98eRspIdYO4TECrIh3xgza
NG5Fvh3qsfia+1o1+X8kcDKpTt8B1UCoohea6nlNA0HYhqRhUpmXg3gb9tt2puNeTr6KCS6Wiqd+
varB4eZyK/aocJ2Xt2RBDIyrehvIR5P1P1Vc8lr6dLyKUBhsEwOKHH7r6X6ZSOJV2W76OAsdzqgQ
EX5a+jC2NLlnlg/CwMldnbloIO9gUrYkOPME2LI1tC0R6jZsDchINcG+wK2mYVWLwvl+/TPYOx+E
oCrrhhid9vAul0lgcAhUvp7AsciFdvtRn9u3XABLHV8M8PuxM0qVeYrtNGnalr7GN9KagRWJpeWl
+zluG4Sw9NNeytNY02SRo17hOmvpV8wfaGlu99YR2678cyVtBgttvxnlSnJCOAZaRVPWib2LW7dd
mXj107qMV+xNvsM//i78Y/33wXpv0qXN/F5P5HkmYERdLOySuYM/kSMXbajFjsQxE9CRTfm9FYpn
ddSoACsj73RrMTTHdQpRg6ia1E5Vy+xSC0mCtcYL9TMvSEr/BUarJF2AYLyDvPX4advpUwQNn4Fc
3l6Bef/IkZmvkyEkvuqCS/wTKs3M4rufPeWXAD2qALLxKsxhHS8c0Ruj4ScwgJ25JTGL5Yw50ZCf
18j34GapThcyEwtoaooZOdLTF8qrr0JTT9LIVM2MoLqoUyvwIhZEvi9wzLr84gXaiKBsvgTu67qd
Pf+145xu5NjQ0DmyDs/3Z/vZBsnp4cURSi3jO46Sf+8uweAtdwzNlfklo0fM3ekUh6EqOUNv7t46
g4lsRK1IzQmQL4co7aJozBP/GSagVjZgYX2gULrvjAVkNK3PDOYzdr5bZti6StdDXB3cb95r6zW0
zWvL02fgdjdZzggOlZ1o96Go4J0vB6vOMjNmNN1YE2PWpQLnoQuLY+h7yUo9qavaHfVLUq9lELjO
CTkLzGObKWJ0Mia6cfAQy1PeJC6HiUo79KaZthhTUW/VRkr9Grv8hdrPgYertSeeIDPqcZKhaFhF
viuS+U08VZdbSjzUJ2EKzL9BojWfqt7CS6FxOPKcuBiuZ+AqhTlgLo3vjDIG4VvbiNlAsRe/Xg+c
6fKdwbtvrhl4oGw2KuNs7PFwH0p5Zpjf/EjT9HCnIKAhk+rAfrNYNfM4lbSJxLJU9IQgPqG6bhal
45GTeP98TOUuplQ9mXqFMNJqx0SD8LClj8Or5LMpNkbWOJpmS3zj5jlEeEnW4Ut0eB8s4nqWw7l8
CjvJ13UrwfDmXXTjruNqbzydLlUmJra2xUyHPH/HSQ+AQVmzM0Xi4UKGuk8I7Wi+ngSn9XWRB/cs
pqtd7JzAG31rS+XzrDGSN0iw+QkC0D+JpA8RVBGXV3mnW6QbtWsmMFcKvlLnaY4cxfv0G+W3A7mC
Wq5sYbnSV7hKaT5fyPb4Uj3Ed1J8yxKGGS6f+CP4fjJhAy/F/hB7/0jRqt5Din1V5atlizr1nIMz
Kxl/pgnsw2AM8TR3W+Bo9TRHdc04gKuXnDO+x7QcsdThb3okxRrV1CsK56VoMt854hrXaqrOe7+c
Wg9GW1o0mdfH4Ig8uJsiHtwDaSuhxV6FPGCMjtuJquOwzpP9DU2YkyS61z5AMkjEdaHU7Ff9ksmU
xhapBU7Kpy2x5IJKKYUAyoED/SYjLZ5vnc35+kV5WIgTjR6aULopqvUqwRqESyjv5zQVghjdWxut
SjZIz7UWH5kxcFwe1vjJoLkixnhYMHNfXFv55QUBp+1nOs7zkPeHaQFAtv676CMGl3bVrhMro+57
eGJNqU65nqy5+/OpFlGIhrNiPaaKqAsipK+FHcW/A2IiRWCF2P0LeZ3bIrA2Q/8zyUc5Q1e2PnFv
9kYXP3De3UHiJ06qT7jfZOJsuZ+PrwxXo2zG62X02sh8FOBdqn/TFHCWkQOf+HfL+szi9YIb2UQT
Y+yvKktymit39dJ9KkXY2qots8YY9lc76yj4urkmHAQKcE9w8fOO4o8tKOfQJLmKxXdQPpJYKQ4Y
ie6g1g1es7H7vtEpIvpahNh0wETcKv7/bJFkmsKvXuNi9XotzVgBiW/ktMAl+yzm5nBual96qyoW
26MyYK1RWzT316CsuSyMSwjmM0M+poRin1xsR6E6ZtC7w6SsgUi7jj7V9W6YDD1ZYX11jqgtKi3M
Vm9RqXFeX8lJuWP0/BPP2Z3cbn+DBXthHLIsM6Zmlh6zmGzaQ8qDc8Omw7cQqEW9hmn5/qbLRqtv
6XmHKgSHCSiqALLYhDLd1VodwiK4SlpIQqav18MDbUvH6XD4dHH20MSDgLmzIRpXvAd3zyTSZ3TE
XYzVr2nvDFhFJmD7EeKIpcP2MJTYTmq/T2ogPWspCmC1/0DFnG8uZq8688/owXtUNoo69Ehnkwb0
ilVyBj7WQnlUBj1UNvEn98fr4VNHq9sb3JZBDCJ/vI7I/kvJiWrRqgUHWK3WcgCk8taAC1HEHUZN
iW8M+AEdaRABXyx1i7vhG8MjllPOLkObLMlxNQET8Lgx+LzzaWIDVDh2qSwbXXWHLdPe3PQM6rhI
YmnBsjmpVv44C04gggcFTZd+B3pvT63o3y5/S+o00jV2QkwvMXHeXdj1ZjBMaJnnG9JLrxR0mJZv
anXGgcEMrhWbbE3WSE5rCSsuDUy14dOv2Ri99YwWJx9AZxea+d15raVRrOiydYO72dViQNPF+GnD
MnPy17YZKOYg0HmtC7c/9EoN2qM9QMgoI2Vn9Erx2E91KtIHsBzp2OnWcT+1p4qWKhJOFmkO/KrR
BhYYKvIWUoSc2tPYm/XcHWrlt4OXCGhJRBXuEJhSx8yC6mc/2FlWoG2zdSdsNHjiubGFsIuBwy8t
XLlAo224A7aZYASXQtFra6z+YX29lxf2ZRsapAJ/dghdZ8VhsIrPG0BKcbU3AapHO5Mx3zpKtKna
cotvxSVTfdq6Ul60EyMBofENbV9DUUvXOb77jFMt7ollH9pTBYfi23EC9RcTvQt/2Usv8kbW4boT
WA9D4HuNovm8rq46rPN7ra0eMu9zCr+PbvTPjmqXQSdQaW3QG7UAwsQSmqGqTyrdTRuEArOopS0t
UMrIqFaRv0XA/f+f8v+BAjwxZTH4A4EcX78ZnslCnxV8hf3UUYCYFlItoeQIOALPiblUAHRdYgaK
fE2nbUHY6rDTMsUjzNXQ4hTblcyZfUwgU3ygh+ZcWHGbFdbYI1mLSHR/bzMLxHSBcY/uWoXwUYo1
bk65V9+kIag8o20rhOfo3GCZ+dqeo38BKMkgngtrRd0osYc3CWUHN8nBWWUOpfs4GFpJIJ+urCmT
WFJso2azeci2AE+p3J9Y4adkajhaUZwYLWARlmKYcQheLOVI2zsqaUFPUX1aCoto/3aDKh2J1s4c
wnG/bQqZ59tzN8CTPpR5fpMTh89cLIGHvmObm2+66ICuj3fF8D8fZ48VJZPhYH4jEL335CNLNrlu
HKAwsmNLSZGZ2usl0k7Mj2OrO/CtUx6DRmX+CFYcvcXX9awHTwNpRdfXRHCcCAmb0o6hl1TWZvxN
vOKp8uFR2QqsMRS++kMY2p9iXbgnbXcwCe2Sh3fK/6qf3QfZCOXm3Ghacn+h8N4v8Pv+Nyf9WKAl
DWEfYLwy+ZCgFISGgePQwwYfFdA0dFrYO86EMk52napMPippWKEhtlHGhegVimviF6xF0h3T9zd5
77JYhDA9d5ewZilrdKnR9nzzuk8NOasa4j+WjFkgMJ8ROV48/N68fziAe7Mlp6dpk5erUF2ErKnh
sGLx6he+lIkt6mkVBFBg66pHTsp3+SeOZ1XmPngRf5j/JXERbM29N5zxUMuQXJxyE+T7KlDiBkHF
A/+8IDjm9PrFin0eSZ8WJP0+VKnCIZpptpGZGO3cFqkkOFzJ/NbUd6UEpE70o92mYyieO0qlRpFV
BZr4rcVHGO7A7iXSrvotwZv02PW7zTXZgsUzeofDyDAZbfEEEj93BlITG+MHCZDFGcTZh0g98P4s
z+yIut2KXG7V7sFECJF4je0Iro/tivpT2oXU79iL+D1F6bm7Ysf7te4XWtFbkqaXlmA8KvX2lYyg
jJ/S6OIfCTewDa6Ev3z3M+PYnwXyOZDcQ3WRbLR4hf1akKmkC/W/rv1TFi/lBTvUWZ2cnW6+cwCq
MdlTe8xiMeenC8w7fc8jjdv0MWORWYQSbjrR//9eJVJw6xXhj5JNXcxGjJQcLH5E1M5x3p8DKZUI
sSuzL8OOb5jJc97DrtaSd+Td/Z/InTEHUUyuwTTjrJlUMUrqF7QWJhzJOHhmErJs9RKDmhsghfpp
vKm83DFnFCMYpzW+O5oErShJPmxOIAcnHe09Uzso6egAjNSQC9fBAKNnb3me9SU+2ELrpe7EFamD
TA2awCmRGVB299K68KC45FRI5FOWCvJvPlqtNnANPfMLVIsZre49txsp70By02jKicNFkyr4lshG
E8+rlyDDdGAa+CVbBtc0fcbHimWt+nRp+4mkvb3SX8xy2arLHCJd1WZ9NN9gUoqVMRUqCuwriGSw
kLfLPmoYnR0nlHoknIl+ylzfMW6NP8n7fL/u/onN9uCQP5kAvCGENVZ7+cORClgvzj/HIaqtMpXX
rjBwQi1m2m9a1rDJBhNrfMTrgqoL7DSwwjkYCh1XbhA7QlwtZdkne+H0B+xXxz94gpAuykqSgrmv
MagLlraXgYZzKpYPKbUQVWFOiBIw3TyMnGTKstCm2NuM8ieco7VHys52Cm6GWWFcKrdwVFk3DUM7
dAbtAvAjhYE3U5s/ZIuLy6nitCrhILjgHccRjm/qJzLSk40HnbiDkZeiPy9wZwbmUT7OSnZZxoPw
QgaQr8OTdNSh/IKh0hjtjSGDRZC4Q7ryAMtPCsBPB2ipXW7mynrHexZYJ5sARFG5Ht+zBB3F8Zgj
HAbdQzapBi6uWghBbuf1/jNXHHIKDHOpZglcjVCU9gvVkepuhgCcXhhs452RYtbdjJD1rXb+hf0u
CkBZzV/M6qPdTqOv5RTnT8/DbToS+Ryt3TfzsOW/gvDuU7h8HJRgPepaonhiI7RoY8/J+hmSZbCd
C/sQ+lYpEOtFkga0rYVMdelvGf4qXN7QnS9Ht+/gOowjcCLa289caTNIe3DmH5+CGjup/82RQrAk
pnkwkTi0q1OWt9+HN/+UQl8MLLkJcOjRimUBIoNaXZJ7bkxC8fvfl6zoQkptuJOMWd5+h97vhXM7
iuho7nk6J1jkmiwDGvOkRDpe3txlN9ylGCgkGHLuUuMdakOtrDQfhw851GrLmOLJqV4eeX7yw9RV
TOH5xJss/75nORphwMprCJV3PV+AbJ1FBBVdkMcVmpYYpiGQ3mAL62PTyUw0vbph87BzgasnAl1I
PGGOvnVeFypK26zXzVaUpGrHdCd7vIZzF5fvqBn/yWJX89/7YZOlJZJ2U9AI8nAtYbF2kmYcLwDp
6oz0Myk4GVuNIUh5YDGqq90mZv7/PEuK+VZBhBRAhDjcKNIbR788t8+b/2RysUZuIGFP2BWyatK1
NRil8fDZaEWzEEvyhQd7gi9zlWV49NkUZPo4v4IvmS6eenAbjHM/fRTMWAq25MFKqrSQS0ZnKcO/
g5lp+h1DAXfv1kGk6edXwpUEiEKvxdPFZmGqPThFZISc5LMnAbCVB+lAtMuNtsg/obXJcTPqxIxd
jpu0mWxn5Id458PowZIkPKbl/K5epvnhzta8kINtM+GQ5APEWT1eHqkMf/SkMz4KTj5CFuxnFgfr
VVI9Fzhz7k9BlLuggAIsRt80AsDzAyANQ10hB59COdTvPzKXP6r63ysXprb687orKZ/DA0cpySVq
6VOJpxNSOb7Kfk6YrpcJ91Jnbxk8sMdGSSBY0mkxj1Nmx+TUZtY+JWpvMddhc0hX71GK0gshpUTX
gTuvepDnqbS0w3Tl2H3S1v4wz3Lm7Iv6vbEOXyRy9tMMvYFQ+cJrXu66J2H2WNgZRcWenTQgFTFq
fHjbnA4V0GiFMUZRn1iJRqiHGhi5mHB/z9xmv9v60XfaCkM44Vn/iJ68a074niFrgFH4QdKaSviK
WG+qbbcRljWveafSZze+b33hHl8DQ67+uATYRtBk4GOapVntG9hWo5Vd7v7TsrsAm1x/jwZTdB+0
IWljByQNXHpzbFqeXAHb8LFPNyLB6dFMoBSLJ+5p62UNknrAYHgRZBl2PK4GBMdAXLGzO0uan05q
Lvp0h9TvOVoezeL2XBDuMqN7KEJrSGLgYIzNfuX8ZKFpN/ZnNT8pnTIZcD9vFXFZHUiCN6Tb4tFt
j5fJ0ATvj4Mo7jsdFEej9XSATu00MzK8oaROk+UTP6XP/UrbmjWsojllDDhWiNaz4KO53IRVivhX
c14M0wzFnIaqf0fggfPdtIGpZ/yxnGFOA0aaGbh2LGc4T31vQy1tWcOnKRKLOcURwI7BE0ykqOtJ
YIK9RkGqMcnsycdndSGn5r/hQuEC8CAxfnkYdLm/Hmo3P/QWjuwjyp0JZuX7UTe/B7Ie9W4VOIPZ
2BKgUcHlOG5oSyss4kzpYf1SykZf7mISTNt+pMawV/zE4EVNm/TUeGYkm8rwGSTLpeFI0gNDvyDa
KveGg8WXwUbmNHfBJ+tPsD1CA4wTN7aQNcty95b5ejBArTcj7O6VjXTwqVHG9PTJrACQXo29OWTb
YoA2Y4w5iBgmaG6mi5yOzKsudkUNUcMjK6Jefz2gyxKmzl2Lsw/uYv6vbDYdksfFoceQyk7/jce/
kN3YN3Q9So0W0Kz2T7QOhFoep6Z08clCKZp7mf9pP3wZhUqi5Pdm0daFB8w0Q3LvnQKx/g+9a+dF
IUr9OQPovA4l+/NAbCCOPbeMn5NX4IDhNytgl322V4Xltm5cvoJG+hWxAsJh6YE3erAhyCLRUYiV
48KGU35tChTXbzVRKRucy05nbQpURow/4hw/VLDL3SZM8cIyp5tTeYYEOq+ZNjaK1FsawiKf/R44
2YN5r/Ky16JCYV0sx6wwASjddBCyGAt2yKwtj6Lf6XjSq0nxXqYlEAf4Cd+UH2cvhj3dc7Dkj7qw
neTHf3u7d9NQLG4FHHFn7E6JbPGDndza18+FpKLPlxnEcD3elXtvI18Kpw/CnB7iGUiZw8MFCy/E
hbGQwGmQEhEETY0ChF/tKwtfyp3/sVLnjUb4L9uqSGaVqINsuBeLwp1L9YqhvwJgABjt0zE8qP2k
PyrZHZTVb0tXQgY5Hk72wh1PqJC7gzrvIXE0ENHf7DhEeyZxDpxCHL9lPtzpShDFgSzfMI8iwXLQ
31o64iFrIDrUAezpecRws68baI+LT8QDmfNKUNBFFFK2DwriqkeCPJ33FxovmKOliV1EFVZs8jsr
bzld3lRoy5R83D0zYEzei8DhHJ9mLKapDtA5fs3M9zw1hWVv5kH8E0OyUxt9M/JHn6V0GYTTMgJa
zj+Z6QroSBpd+qWwiedqR+l3w1w4Sfo2uQ0qDN+BYetlvID255hT/I2LWlN8LHpqLDf9xAJS9KyM
/te3nncel4QAdNLCkWqL7Tv1sRKIjDm5S2zDAGWI0zU6T6HKOxTbE6wmCbJc5kqhGFdiDALyLSg3
DrzZN376WTzK9dQbWwXv4bz1EARLXTryxKnThHxnETOcU+pF7p0Hwtva1RP2BM/BfwbmiqyLT9iX
9yWBrEQErbj1zSHilChhefZMXe+pPe3tjuv4zqEDeMKnesukIym4jgxH7WfvOw4xAG8yX4y8qrD1
tzWJWp+ahqHS/aHqmvNu3DwaUF1RS7MDgN0VgE2hWezKsfuHM/Y/2LWp4ckwnXbxiq4T626JenIP
AO3SuU4LdXBc9eecM6RQcrrXM1xUmTUjJvgfbSikUP5Hm+K9ilniVDfwJqbSNQ53D401KEO5gWWp
fk8BSK8Ei4+cP7CKB+HtLiibJcC+0AU+KS+dAR9fknZKwz+XT+EwAuf8m1FY67jn+NKUt/vqjDQV
Bl3nRHs547qqzpqMcqqeOayyZelRyINJcinlHo34G0YA4DxTZyTIGWwH6ApsMBfEjcH5LcmZ5V6P
mN97T4bJhWdRwM67+qIIfpIJiBN+16OGm4nn9l/VBKIZlmF32IPBdsHM9qoAjair+z/2pN1ZSskh
hQv37qLUZ/n0oAwZC3NbRFpQrDJjOs9jQTCp8B0T+Qcz+XYc0uSHl+LosK7B+Bhd4/AUd3PHovRn
BYvmX53emTHbEs8l4pe55WibJ+liFArg7eZh8finnGVo4zzZSRpzoO0DD5GmvOVS+/aX7OhYcPPl
asBrpuQuBa/x+tgls8rld5CIJrmYkN2F5Yvb2VT5Db0VI14B5hY5e/FHPOtCqy/tmslodNXvKcVw
DnyCf48i1t95O642w7vmOmSWgNt1FrD2lkCQBA2otvnOCmH8x7kEDYddgYwp2NvH9m0AZ2EvTygO
psstk0WDZ1IK8dKOKyPfdp0BOT/8qyAIG6ZiTbrpm5dxRoFi2yRUv1Lkkm90qeMI/fwiz1KKv5GF
7hM6idGDtKAARCowhv6tCkdVA8oSTyDKo2f9ajJuI2vg72JxD+Vn2AR9fFntIXwjDNAStxPr56qt
QBY57lqjaDwe1Pdej0kcIRgoBrjd8zMN953/UAd3g5PxzSpAQr/1TJLgpmALMJLvjTYsXESbVgUb
GznYsXOLgacn1H+mxCxudKTTmqfhROFIyA7zGFaWdgrroEVziJSH3HMs7kXj7WzhiLrMI9BvG5/G
pp2jvl3xHDn2/ZWkuNGwXj5aiGKc6WfPO2IEUfuwFmaTuqfGzzcUFubgNu/0K3LgKPNjmZhJyt/Q
4ZTdr4X15m1vQ/QBDSzqLTEMfpqybVkkKkPBYceQJ6Bgy+Qda3OWh9I/ATOcgNSp8kzcRJk8nOND
rGuTBnjPtb9Cm/r6cIuOADjMWuocb6t6+pMsGuWoyEMBvISHMnj1d8i97axUJjYBY+/MDjW72MhW
iAivMaaeVkIhGLmOjJl6PFCmqGbpE2O0kZf2qrtqETufg4zXpT7mOjGe2ypV8FFgXY4OsZOiR0oL
rDGh+9/l7v3vRRakhWxIcIOPHu4HCnD46RnbutVUVJQPwUQMYPjSFc2uM6m82/xKnjOQ9lqStG2/
IrFP1HP7UawmXbL6OZMq0CxmSK9bGa7q6m5Ke+ocMS9Kz2dhHksEIzYI7FhU5vaJ0H0wD9XMMG73
7xg3NNemhwZG9VpuNWDZurFNJ+s/E4gDtNoZTPoKddLHD3TRBjNS1Ysl0nI+bgrab8MlyMgu8nSG
fzGnJmyQmvfNkzNQ7UVKpCB6pBAw3EFx6OO/yUSK8OdxkUYAvhdwMVT4P6060ZCH64dEdNbPjb9a
ioTpSUzkVOKRPA3R4JBqIUvVpc7urvCXyq9iaVIVJ3V4Obj4ig91cXCIl78Y1+sQq1ZcDKDnkgyA
SN/4mW4Lowpw37yfIX7GVSvZPutCNYrGfjtLNocwH2cHTjjBd4iY0bT1CfLpmQ/m9q0aOOx3aZgE
8pxQgylCHnQCYidLQ+UWUfxx32v75wdNQctQitKjyHbhqIfY3LY+UD1H5Y/RZbWsC0C3Lq/wYseS
v72AVgfrsZMxeaQ7QcKhkqCfIKoo956F9iIS6O4OmBmzeyrxJqTBnT4FOUpff7hagblsneI9E2ec
rA20WipZ6nhrSmjGnC2DhewV2F0M7mslIXleIXLWEQ6vuUlf+HL6izGWNQlpys51Bn9FBGm9OqjS
1Sq4Hedd2B6JVzBHk5Wn7ENH5vzxh3fuv8yMCGcrK8CDDYm+UzOahI4XfSYq1knwGbtkD11LpGFP
gy6LkJYg6EM3e7lMyKGvqI7uEOrhq5hk4Scf917roj80WJkS37yrJ9qk26wEXjS1NFKQC9sZKpek
5Sb+87G+qhow4qtcEgVI8HhXLimLim9gboPSWLIxZ1RE5cHn1aEyvs2DeBtWZNlwZXytnoq2xcV2
7UvqWTDH7PImyhHHjIl6I7GJXBvYe1+ynXMLl3yOtawo1/4KTCqoY3wH7FoK2c0uJCX2kTPlDRor
CoGensK95REeBuZLKHse2a9h/suPL7JXl2WURuBGC+mAsehNIL4T4BTLg+7QE8Di89zCBEhQylzy
t54XHsOwgDiBLUhvvXIdJeycdjC55QscOVdLt24yOinlg4mjLnW+ufOgL2H/6Nn41x2o3y9XDr8w
2z6EVurtJUZtme/V5cVlGWf6i5nXhzOB2A7jOUt4LJ0AjhtRer9vihoeQAZYByaqZK6z/D+I4cOB
9MaPnIVxo+J0uNE5kYVDqFw+XMQzcKKSIWy8jPHBBC7vQcs3+3smDshp5gaLgs6nNIp1Nked8Ubb
+BCFLLhyC7m9qAsHvEdP0hXzY9ePVKhSCy2tuHKo/mdQl4fhQaaXOigqUrEvyVXT5A1fGNfMN5vZ
peFtFRoNjzAEHyvAXI4tx4WJVZXtOMGoWU0thCpo7Drqk3u/NN0E578iLH2/SG9NvAB/bkxqLuVo
58R/i3hE0v5RcIlpRtQpaVuWD1BRCrioXJcKsdy9sE6idJBelHIi86i4xQEmJdd72JHSXTADN2o8
P3RsqYf8JvVM2m71jyID9KRydCOIu5oCIfAfhI8ecVipiXZx2TNCXqa1W/Kudk30yIGQKO4oEdN/
xIDrWRf91bKxqVG+j1QBsyMaiP85obS1VUNlJGkimenC0Y01r1RTfIXK2GgV+CMew6B7CwSuzu9v
NakArpuvWBHDKKCajXFVwhF7wEaG3g0IB98wTEpC7ZoM2GIIO53B1YAnzWZZBPJtPr82OwVdCxAj
cpYo7gQP5HK6jVYvzA0M0ehHdlSExPzbG0OQmDgbjIH8AG4Zn57b+Egfwb+MzLUjIwcDcWR1YaYY
99L+WN2Fxe1mAv3TJa2/pCxdk0a7rOkFWJ2oejafZHn8WQkHS4Fq9l98n46JGCEIYA0LH3/fwUW1
fe0C3GIp1KiCvpJLlH7n5k6bbKvuhFYWOuLRjHXHL7V+Ex4oLuuj7WCbBmQUOXMrQ21bFJPLHIli
t1ZCZO2/BGjdosCBUVSZQyK3cGKAZ+WdTCGwR34PKroM7t4c9OJRfkeQwK+ZDfWfVnm3hWZkASKk
Sb3iZLn0KDy9kYZl4Dkud0Ys8632IOtFvhTtT0hrqpwQBAy/cxX4MCF9KABka6fh4En8uKAGG0D/
//mUjdq/prEPDYzt4f4GCHwI0RfHphMgattMevPR0Hwae1V3p9Hb6eMxG9GvRmkzGb/Xv/pCwu5z
jIU+EZyslmvovw9FONU6qiMKcC1aW96l+HKhhAui6ceXHp+vTVUO0PzPQ6mQ/lotJWZhnt4ZgK0O
Ub4weqDpIhQR7zuaxvmVxjW9M7fgLpPWauANzV/R0WF8+m5OOacwjR5KsaAeCBXBD4RG9LMShQ1x
ITRg4iXv3Q0oVb8iTIlcY1+dSMGWf7u2+OldCl5MqixoYbzCng1QB0vmB+hM/nkyKRI9Gb59O1K3
3nzClek4s2waasTIGBC7ym+awJxxdC/MC+qikMRLkiQsQlyiukAcXqpi1Ak+pFn44V49g7DREn/B
4wAF1D9OOBs43rn8+Bn04QovTwizQe4OZyj6AcdXm0ldJf0AY+lD+TRwWE5PzPrBE5XOpC/eOrVQ
uq8IjMlmC8F9TvvReLFgclPcdVLLNwV/w23HPT4A/A0IeiC+c0lXNxzce8/Hr+lasZOB+CmX+EB8
L13jzs6aOAG01cL7LxAkZyQSRUCs1uPN0qdFelIom1JOU+kyxVNGVslQeq54utf6sFRk794ZEhPn
/nMXffw5u7BRoJF5cXCg9GMtCyZ7a1i5/6jVePVVrAKPECM4I9Y1edBfkbgHa99jGVCdo6w/xK0n
NfqqYLAMyn8hqIa65pi2YhFhSpMpBWmLAHrPgSdumk8sf+piU3rLNSiHdq24XlCSUcNoAhvcSwFl
Jg4FQsnf9h2twEGKdnF+pUdgn3nTfFGu1gWoRDGyTDx4KhWexATF4EsSENdrC6hhSS4D0RLYxDai
n3jKOmwmBBcWhIk9x2bS/lmHt7Ks5Cztqf4WKE9uLtdz2mi/Q78/tQiBJAEFze2ZilbOLowYFwn4
hefgaN8YrcyZ1uES1rAT/33YLs9/9UkHFmK2m+9axzZ4l3hhgLLLkmneqyRf3sg3Rn7fFs8GqTG5
30ssGwkL3xV7bt/hxw2IxTXJegSn7vS2U/s7HWit6fxwdSiXpDVYWRLcC4IDn6AZdWCVvoq/6NfU
2zF8WaZqZLlk+XZp03HWtIg+wYGGWUXkA9w8JcAS0WitB1h/AwdvEGVGcIOxXy9khjkN0bBHcRzZ
Jn6tztnUaXjzPUa1FYVkYd6KNJE3aUjpJqJLtHFvFbedsgaaX8sp5LXuLCH/B0x7/qorHYZ+sqMQ
at1CIqzttyfUUvrdi5462OvUIU6aTUdCgzUckig1nxzC0Ny52yfXcwhI5uy9SMdL1ggdtPuV11IP
kipxYE2UmGaea0NSzbR51UhOPRqMNIJGp9sFAYWTuIxg8Ennh/tJLfbbD0101nFB/alDQNPc2cRa
zdXoAt1K8fBtu6+tXoqgLpPWeUMZ0GlIeAKK/jwrrWxp96+ByZoikj2LEsXylhhRnmVgiOTuxInv
PErvyMex4H1dMYROuzfPmg9MQdmZU3GyURTWO0XLoOfMA2xcNBN9pv8LuAoLwGe9iAUMnuTy0Q8u
kOTUgqXaeN985kxnxnTALtR17XZgHUgUBrJTLhsbRfcMCUxEfgCtE+F0iUUI6sPU4YODG2hig7Gb
t8q5XsV72EcVsKoSY79BuasdTadaICWwvtlBTTnIUlWPVG24rVuj7y2DhlKzAe+4iolV11XdoYCw
HLFOvucLUwqvvwf2wUq6jpt7Az3SEk25qd3vN1BqYui0dBhC7SDnGR7uBUafErawa1jRixL5bbW5
XlSugbuvcqyCkwftwQnI+/PzZ7YTcd/M4vPfPPvJXi/4qrD9lC/wxQZiFET9W19MxLWvIT9Gk29+
HP4oy/LKnFbjtIHhpU++bDp1fwXdZ5//X3uSSuIlzQgufgZpaed5fS11jTdNP3NY6Es35e3wePZC
XpFsxhcOHuqd8THeduDSp1RBDnV7qIhjsIqjczAz4K1Yf+psvDNxoR2T3j9EiahMzY8/uxlogyCH
5VD2AJ4FySfYgxdg4DcjDjA5DMulHnV+9UJmwpdJ91G35wZyOHBdx/sZq17pJtcksUihdn9MfK+g
jObDNFrA6ocEoZEH7CMLhg+60uYsvUjXGiLOgWrN+/+fTqmjpoc6BAmqD2zUrtEX2Xo/keWM6rvN
h2IlSocRHJSAeI3kaVAF6gPtodYtQ/jiilakTtBHAfkaafjeK1uSBjXodplTUvAxD2B+QOPsXFgS
aHrdHJkbx7nqLotDnJMKVnSP1AXowN4iEXE3QVeN7RIoabVVub6A1dbORLb2Nlf8XXhQc7Luy6HO
vHMn+IUKG+nZFdseiTPnwG2YbFR2VVTqIb0x7WwmcQaELNfMNd2wfIbDhxqwqXNqjC03nSNVlsfZ
dU0uUw+mpmdQiHHlJKCp9tTwI7F5NpS5uW7u3RTs1ddvRXKGAoPhcptxwISnEDDcI/o7+xHZTP68
uPLHFAHC5WOCfD1WEszP9DKWXcFVed/82etHIJYoFZoKwaMdxE3jNAKA349H+LaxvcFPqVaGYYV4
QsbGyR2e2R0xfgC/Q3P3R6kxO3y4N2OgNSeYJWktLP6/0VH+wQSFBnJ2DJR9+tv2IcJRG4+wTnls
qG/xRNbVbT/PkKX7fhctr1gRlfRyQMeBVd/piNraQFIenkuIbXoEbOXWdYU7zRCarHp1QNj6GM1p
t01u4Xv8U2HwydpqcBV997IGW2yWBIBar/X5avuKK+a6+niSNMCm0YVBWIix7PFmhet5Ye6JCcOP
I2oIe2WMWYICq8/JU70trPOVWBYVbIavq9cQ51HT4tth+qM8LS4RpXKCTLJwT5MRt+F1TRmOD+B1
gSSOcZEn1BaVdSK3vPIbMm/n1Zoo2tv5AlfVz3hzwH5Yeu5o136eOZFgAh/bzydYd+eUcHtPWRFK
wq5g5Luih7jxR3IVUoIpGYnVkjxkwg2KAU0ldlQ9tiPhba6DR+11pBaNnEBW08XpY8YN2OnQkUOi
6ezl8YQgJsV++X6EPEz844ns8Q37wVOc0QOB/TAy6s/6vSmccnad884l09bQOplK+WHZUgkDzyuI
6570Bw+yT6x80R15frZX9Am8CBZUt8nWB4yURvW/BidSdcghmEXCChJoGz16xzlulozMKyzjj3mj
VUXiHiwOvce0sOcVOVsOcbgw3Ntc0HqFusJIkdj34MM2Z9bXx57CPZxFZHk8ovhGsTW/28B45gmc
283Vp1noSt8zMzninhYxUrl92peBf8LT+OXHlZ3nR7JHi8mmHTu9LcEEleRmloFBFDEvDiwV2Ech
ZJuQYLkPFZ2y1TPFLMsRd3K7uPz9BCXxVw4BcqCX75K+VlHCYaG8UBzHBSM6f1sS12X+ZbPkUCEP
BB1pL8qbQE8tIgRmXAp8WxJRgpZgl30loHQQiyWb6SFcdGBoHxTjARCuwJNMVauYdICE6gi6FGJT
bP/qPlWwavLhNnFGrxGtVG33XwYiJKjqm3PZZtvvj2nJt4usSz7wixq3sZCtksByLB+oGFhxyTJI
zozHNj+wMAZ1bd40xCL95z8FiDen1LFAvzVtRdmyvjHN6b3tGWH/Fjv3sGPjzMeZX0g5HO1xo2IR
BehBRVh/qkxDnWFia4fN/c7CK111sgW02SXL566YVycvJNcWnNi4MQkWIp2h6M3YiGQBrdKy1pue
IV1J7fjDOPhtHqAHaoPRuXiSSanyWgSYZb4kun2+V+eiZreunrM98G4vVKjNDX0MhYML7vkGmEPO
BVj5D07CCxexTzU7EsAafIFoQEHLJHmvomx5tXYosY/MuaXvOFVTYyj4BnnYeLX5V6LRrIOE3MX+
ln1iuuhVxu78covaC6xvUDagSjMb/2zvqhkBSAenw3NPqjq5ZCNZjPo9j0ijchpovVVPcJPap53j
84OGToGmYjG2QFhHEvXOUkt+MQTfwV/BNSqgndytT1s8kLe5HM7+MU2E3L4pdPxzicTvBXkcK16p
8w1l3/eB2UMwbOPAj2WU1ugcf8YereI3YkaPwFlkxhRUAoAdLdkQNHilHCc2U7gPjDfPtdSfHk7p
CYaEqUPG+sLE4MQJ4biyp4cTDk2gfdCwB73pAJfuEd7mKGGapGJoB0EStSLbxSGn0oZvY7fsQjNd
1OHTrZu6dU+zQYblnqco9dFAgnC7WmUhH+eEXu3bHRAe+d7hguI+43pvhz7XjLy6Xz+NtPQhuCAH
yI62dyQTwPtuvYL9bQJZr4Tbe506mxslRSDK5hcyVlToCvS1rBJKYdmWj5AgQAA+jtj8UQljJH4c
Lmkktxbeizssb/XjooCi3S3m3xb5r5eXBOXaHN6fBI91+U4WcAlE9F4qJyVXE1tPy8AL6MGq9fHE
J6k9xZAspJ1cVCjP7j3q+AVf2s2VxaING9eD6yH84B3/Xai2O4c341J8KQBOv4i92JRcI/V1zih7
D9yEx83vXa4k9PQSCI7iIIXXkTkvO9R/CNcYQ+TkrOsKejxrXaGwuVlwshVdM/uVwdSAgxeJLd8j
Gsy/Iz8ATkWdZ3K9pn0nLWNX3qyWKejhRFMzRl8q7NGMVzza1BZC/qtNEWJKoMxczGz30YyE1cdM
gdDIrDFwK0AI+73sv0L1A7Th6lYFuBUAwxf0OL8xSbcO/109K1QIzH8ZCQQvsyERmAZwqAz64vQu
prZiOgXRGsNOAkn1nJGwYu7AXImG/Eypg3jp8n/F24T+eMzOeu4f1JDomY2ngiglGRz7lz2FEq/v
WGdM0q4Y+JzPr/UpP4HpiQuKiFhdLD6q+m1EG30qzQaLmmOafmdahJCnoIvQJB3KAC/3ezSAHMnR
aTwnk7DcIGFNQV61P2DKdKT0ZDYrlJ2LF7M2cIpLGjM00f2QRr8NYrfWck/c0eejPXyv5JjOeJ1X
LzUzTtj357FcAT+HpN1amziBlHUKdZrw4pVTTqcHCIWNslf2zRK0HMjKuXXWtp8hIOM9Z042WIId
44L1QcAIDoU4CrTZbQADGXppsNfAupQJUH6JR99IWOmxfMOKU9IMK2er4G05l5jYWTJnrH2rUcHn
WNIMU95cylCrhJXgBL+dt82FOvKDz9QzkWAS6Gpg5l7ysrmhxkfd+ZNx8zhXOZ/jnLSk4G15Zd0F
IdQDLOxvxoUzVcoWZFN62i854dxqEjaPu6T4+lv6U8NAQO6TEpIvj4RngeNBtcqF3lEXglzIAK0k
c6IWogSzPPIuA6CaNMuJPJk0pPA32oqxVGL0oA92YqwC1kYy8wdUdFCOb7jg2BG6fcgS5NMBXtp2
RIl0W/hBKaAdVxJzFA4tKbMe6gFxEBDyj0VKDFPOmRJ0MdlMs32P8vXEmEJjR6t4iidN7f1lYqOI
nDLIv/HDDlfLXJEJcrbDWgzTpRbyTjlUQyAQvkq+QNpDHB8UDUA28EGZfWeP/5mC5f6OwnAQSoAm
oEUwl2xgYKSu6GfnvpeqWPlHqtS8B4MKsHsJYr9YDhKiEVyQlAeyWzuGOdq//uPS4WvD05Dk69O/
ZcgarCgPnyeEcuCICHnJyi4S2fPPlCbw+nwpbLiTTU+0vlezcouLgtT+d7/0mD/GzRzTUx9KAAkW
CN6BNOZycwws25Z99LRk7Nf1SRN8WpXnRDdnp45E9JeCj6YU/rGqsZ/VpqOgNGQ8FJxA1Sj0sqk5
hZ8BXMkhn6DCaGqfX40OAWNmAksc7cPQ/DUn6ucai5+1bEoZJ0zeynG0dkCgE7/8ZEgMdIH1Pv8t
pSFEjGB93aARYXz0gA5VOfzT3K9vrB6Jmst13l2dAZaDZ8kguD+dBQdDRa7OTFcPWQU0rDxfR8/C
U3aiM9QxFBniOwVHi/EWtLBd7BlLBFd+jDYT/E10Inp1c9657/J+RnxHKzRwF3dMmBTV38xdfWlQ
LSWwQ5usEO/f4uk2bLGvD96zYGn81VIy8OaaLRGvB5GOZHrM4GnD1PDAse4IpabXwO34+Wnl2VXm
UGKxFGTV0tS81HJ0pttekA0eaILu16eTy/MWDnbpfUnpZ1DjV2LpzPow04ekuunk5DpqkNE1AOjy
nDcDBEGTpruCZ+aJK9+saNiib3lDKoQhutaQlWMsNgqTjWGbMWbWQJwZD/I8GjOZ7l/k0+V4SOAb
LTjrG1ygFr/ztyM9jL9iHfdjD45iE/X2uwSk+cRs6/qHO50Rr3Ss/hcug/YsN9QqKpxESslO7auQ
54XGP28KCR+ZKHYK+dde0O5D6IAfchrD4F8kBCAOPJTtgKyrcLfAUekJGpyLCZ9iNtQvmAqh2z84
71/uW1C+EmUd4b/LTb9fp2IhDSXjg5viF4qxJQJyxtQCHSZrGQP+YR8X9ZjxGAVWx0n/DkD4D46Z
Y3NKED7bRbL9k7U+IOG73S/WjZsz8If8XhFl1A71BKckQQx9D/s/hlYvnW9sBkeF/BrBdD6zgKOB
taQdu4Q0AyHiBWW46iQ8jGeMlLo5+grdrhGQW3llbQb2yCWkR2dvGW1WlBT8E9U105wvMhH+0G0K
KFZVqsXN/rTi0Au6Fc4vEeTOk5g5ppJaBiG8RJrD/FxSKiC8+WrOyz8VRAh9ZHluNDPs32dbIkiJ
pfThJNyS+Hc4tteR3mEcP0ZkJK3bkHwzg/nR4/7qkJkruBLzwfs1N16nhHzDcWYbDefhkfJeT347
Ngdcj2dfoSKafBCzgBmrkznieXOmSDwQp5gNV88REswkJySuHsW8qPNKr5Cmb/MFiV3VSoQ7SNEF
ORfd5mZ+L8/kCsphNTZptgdD/4vEzxSRX/AIRRohRiaXAh6NBPykToWcGpFPv61GiaBeENfF1LCr
vcB2dGbZ/YXNn9eDoOkXziBcqNF23AVe5LkKbcG+xRG1NpWXML/f+C4Dt5A8B2i6L76ejZVObYh0
mut4hM/R1smBVgZnslsHxlOAIYyBo9H7CFV9Bv1swcYeXkHsbvIQT0LW5wq4B94oR9GZLYj64JSb
5JbACzCYQ/l+qtGw+oOTLfkFrrJ+zJ7kya2Hi7YuoRoaSE1q/B2Lhj8VZb4K4F5WSJxZS5eaQcRE
t06SwDYAWzcTwK+mf6FD1+Gv0c91lA7vib0EGr1qx8xKGzF2Zi8xRFzq5TkWuLwB5kwt2PGbx0n9
r8T+GuhLk9BqCqb4CCzRPC0Na6ykLzwQtf56sTFOO5GMI0TW5I+nktdL02elw1Z/EHZlMj065K1D
QHxlTloKCjSqXoKceNkZwEn6nXDr8/zxzpWDaiAUwrWoD3PPVAcDNv/p5JFngy+4dbkHZSBUIu9O
DkEjLjpiIluMqIpdCO7VEmMMjdTe+r53bbTMvKvHRX8CCfuJqpJ9SHHbbd8uVj4948CQURfUJBoF
QAnYR93WVgiTPQX1N+kOruve4y8S4K5Xp1qZfgUSfYFJwq7hE5Sewva1x0GKrQffR/OkYHYipzyK
17Sn5RCqhl/3ia2V1/JWaMhL+OBmi14gfYGckC3bouQI5/NE7CoEjNwPgv1WSEIDSuWJxjyJ+Dqy
MxQezuXNrUhaCcDVXi57xLEMvL72KncBr89TpLmnb8/6c17AXqmsTtkx14Jjh3TO24PYYVaNBi/j
4dukCGlbmQouoJkJSETxopPY7GkMh3OutvPYNcwbplrHt2lGDvTyqNkjRjf3R1Gqv3iz0iP4XwBi
KrdwFMkHnv5zyk/rC/WnUD6ZwnMtVMTzM+LmFfNV2DOhtbCz6Jx8LqWvV2vRDV8IdHg33XlfKAsU
nbHbJ90PDa6x1pQue9ufmmI/1l6kK8BVhkdr+5V1KJ/qqWQPQeOcdbbF6ybnJVOnQ9XRWR/7zcLm
S2cUEaeTJKFlYzBKCcJfQAd7TUxK7IUsim0egolrxzrX2H4tM+iOyMnmVou2JrG1dQufEneK7iCN
jHh8VXYl4S7HmFdiyA7XN4W0D6UCxWmVKsWwwUlk/W/vhtvbXdV3RjSWti98p0Ir//cfNzsrF3YV
HVDWh0p3tWOk15IvmF+lOYM+5LLFO906o3qkjKAca9eaAkfoRsIrZgpoU7ObUp83rE+G0k9uvf4R
gRiX+RQTucOV7XPUDf0oatYQ/4KNO6lzZYTzT4gGd7D0m/LUuw1gwDfBilkQmdV+4UAXcH3im0mn
6ZClYdoU4NS5hPc+5xxDdMOgdDzenjSp5AhvfnNhtN8eRQxiUUP6NWcD6fIVW1aKLIuzT1ERGK9X
Vx6Y48+GjRtjSqdwZtoCzeJTkwEqdqNRcjOf5fsJSAlti3oCMAewbnIXXaHx1vsVGAy65P2MD1Si
vMYQDKMT++s42CWfZ0le2Me0G3l71igHeYXlW1TopM8qA449q2/nrY6WTUupA6ua6U33F0dDOFAN
bC5CB9yxjZ+/VZAIMbDX+aILqEG5Xd7gVqxeU2Wa2w/6eikmF+B1RIoPe54WSq7/d5KXiLa5VtAs
5e7d+ukVAF0PZ9RIYYxnVCvyvZ4IQQDlfsHcleRTH8nTgdEbhbi1eKS8mMyPk9YR9TP8nE9CSRIp
syKeNGZdVGq02TylLGTm6fMtsdxE1wtbL1dMggHK3PSlSfhrOSSbH/e74s8t+ebDavDmSmhTiPUb
X5pVZSAcMEUgVFRmOnCIb5mvbZXiNZ2uB4AxrDmhkUvI9FrnRpbp/fL8fIOd4W1fnT3bxRLGHDW/
xWcVY81tGIv6/dlvQkXfGD0JC/D/5rMmrrxlwghAmrOUNLWuH9BcpJPPFiRyTmBeYluSFEzGOK52
GlSkDh0mGm38r+3CZq5QH8uIm0XRQZx70ZNrHtlG7MqGiVr+h98iOvrvYls70Tj0TD2924wiuRlB
vhiwjAn4xTnqVGKZlBAzEnajdWKVcErcFClUuKyXlN8SMvTd35+Wht4cEXarsXffjGfxN0XBPFwF
nQkiwHOxxlQfucy5Y1Imxx81Yzvk+uwhstJ8kT/qBZ2ePtl6lVasvasI+V072wjtEhrnrB/A+hhj
IkLmOCZwOaEWE7zZ/rb31271wbukcVdjk3wlY+SFd9aLZkjRBWtNJzRAc/SwFZfzW0qrLmkqGVzR
fWOPMoZZn9rFUzCNDsNeIrtAZtQFtvWePlqH3e0HDg9A7uMJFyFsUsS4K6wKgqEneVgQC3DEti/c
k/5XtWc43guJimKMCVLrf1uAlUaMfa9JFW+9g3vs2ojergyVBXutNjqO4usHUiFkyORlyAwGVM1T
DGPlYamFF5ZtCcqOcCIaiGkHyEnJ1H9g8GtwSZ9zVATRHaYkV69inAsoA+kl06f9NV/KjGkx+Ky6
K6QOmrLIUvyu4MK4z++MDVX6/N6+HK31KJjZtabS3cz/1KcsXlYVP9yYvEWR/776N77+GQbL0JxY
d4oUt20I6Hm81X1lHfslvBrMMjT+eky8IoOAV1iJKkREgMdUT7a8JjOliKq3yjZL9blxMEXp0YXY
NtTzc1LxeXN9YsA5vnfVOkn3q9hmU2ez7h3mfL5sEZF32JVdczKQAPX6GT3gMtVxyFG2C0OSzzJ6
VdUwRGc2DN049Uac+p8Znq2Glnp57/m5ODFjFyhoEqVqqRzuhuUnBjhNUCaVjVlCmsZpBlQ7HKua
9qU+O1ZlH0F9IquSYtyuw/ctY4upSlkC8tdWD2ZRcj83Yz0mY0oaOzcCs5FRiEqzY+z3nM80v1nT
RsRdPBRcYGWcuTDVs2ElYj5Qs2wbSqREAiuaC39JTSkD+ard84if2MXSR1BBSH8euLMQzGp9VeTe
gT7KJ2Bwd42DZlT7EhyDu3rcNSUrDUaL1Kk56V6n/pn6tES57JQjxqgO91xqKeh/khexUz+G6B6Z
ZtzYLU3xnus9hCEOJrZ0NkteTBf/E71bQtZsFnrgTS/jQ2MgSYZhWzh2kbWnb5FTpN8xMqUmzrYE
TKq9FrkiLvxmimDQyJ4+W7GYtgQDKRjSFiVitWNinpo/PeD20C4vsW0jH0gKh84I6zK4nY1A/jvZ
pEIH93VJlQyl7FP1Ev3ylykVJL6Y5XdtZuinvtQp4ZRpfxTEbSddjzVD6HArFEO65ZP8crqioh4J
bvVTVx1tKznm82bwH+xIgOtgnad052gni1Cnj/+GDonDWdNWbXrX7jx2e3EJGKu19NE6uDCIGiIQ
xR1lRLaLiYNh9ToeKLRa931TV7gHPEZfsp7PNETIDRYEzkrHkC0rLP3MnQmol4DPls9YxZJxZn8q
Kl5MpOPNlvC5LTqeR0g7rniBv0e8zcZVichsciN8X9j0YhzZx3Aop8IH5dvBgKm07bmPrWpxpXBP
dX4pPeGKWW68yxwmd1xlHdAxjhKCP1JEbFW2528+kVBMKMHIGr376sHyd1qpRBHotlPqvr7WaLL1
qV5o+jgwUqALDmKIXjE76qfAXJTMKu6XepFlDRi1A4+YkswRQC1ysxPCcXVVHdg46yj5WWHejP3b
ZE9nmBi3tccSL/B4eVtUVUnNtwD3F/hNRWn0+OH1l48Ujf/7t+hr4iIpWlJ9VYj40/V16MyZjZHo
0Xwm53sCjac9e5qeQt7Ym/1CVlb2Y8KLgdZ80japwcZjp0HyTIjkiJjdPN6Zonq8MfJsgm0Gp+P5
SP46j2NjSTMcJedJW6+NaArpogonFNRQzK1rzefi/Og6FNS2VAXoFRft5bFJL6uSu0iyvs6Yvaln
f0OOR2hHF2XEVps4XPo8XvUYKO7UMZZj8eC51OxSSVsTfjbQj7uCNva6GF3za7UszmSQ2P4elVlP
3Giy3hLs3PMRKepJ+nNByERcNlMThwMXCa53vWra6+8hR4zrBU+ww4GMjMY+kXIpeYY7dFk8g8Iw
SJ2E5rFEZ3X7hszYnofm56yhR3Bxd0UPBW3EhQJDusiSHhJb+NfJ6PRhSXOZlsex+thTnE7tPfV9
G++HovIR7VcjgOvXtC0h7GqoI8OvzFg4RqKPL+2E94uDbz1GZY3xtIgbOhgrnsgrGKYcRJFzHLvz
MzhD5Q6Qh6gA8rcp/9ESEevbV5yOF4DISnuGBn6rQ9rB0ZQ30B9ONvA4S4tBu9DzQUCtxCuOXLvi
m+rjx/r02+eHPLx7wN3y84IBSgQRnmPBrT/RPkAt7gUm7+A5XwB+LHPKFbYwZNpppeNHOUuOSZCL
AiZilqosyAU9irNP1MfHfi06TI5DkTyu+QeV//gZrCVZeW5dThNx6hmQ6q93vnWsQS3FP9x3fyw0
CWqFg+KY2Ox3GXayIuhbaI/aQim98Zl1/MggPiOYhPvUp+67jTOmESVZpQyBtCduX9oyQTV4KG8B
T2C+3oXtBrwR5gOxruwbnx7GlVFmh/h2U29mUPUBhAZmG7kBLj521mTcV8pYWRnePCbpwgjD49y8
ICIyWz7uhFemGdDx3RQNth6DgM9IXZdo5W3eXP4jGrpMbVL3a4svLLR0gcG1KFYlC1xYZIDw0vTJ
6rgMHXQPU0GCEgnIJNBnq5p0BWI2x+swN6ZbKnBRboe4/XdPGFVZ/r4ccEmE+XCGFo1Y8Sxc9R0q
oxW2RsJziX8MdAqs2x8495Vn8IdxWvG9m8WG8JonMH93G9UWHSYb/DEgdnb2VNJpZYxAQk9w9aNb
WhZcxmF2OlfKW12mB7dNLDoN35UJxf5Jt4+M+yGA6CRh+s7IRzjDj94MgzsuTOJPrdCQYKlI3OW1
6tqln4WU+i+iVVUONU02S6l3oq6KNiYEWryRh23E8jlmDURd0CRJ1OlwSN7AXQ9HSrgT+zGNGM2G
Plbb6NtSuscaFjfncGdW7flcD6VZ97GLOne8a/H9J1VfuQrBQR1YoAEEun1EIB0TS8/RogVdIarC
XSc8ZFTV68WUB1oZRxfI4PlI4ETgPd1XHjLSA7JsU9yIPd/0P0qG6TKLQuPnb70SeyBmJV8sgSYM
2rkPXqRE4Uodbv9VVtTe8w6K741575qW2CR9Cfp65y37Ms5GthME2sYYW62FREygJjCki+7iexkv
ZcL28eAu/yeaUdi+CmkWgqEhLZK+AUC+5qCNqD9pyUTMWPnCaRXkoPfTZWhK+Wq3xLpCA85Sa+aU
XCSfju6SlGoet0l/R4DmmCavIs42/ktmF9ufKatV4IqmVmxvfswhFPMeYO0CpMDYoDfvgp1uFBQj
8G9d4BY7P7h0t6OJfHEBoShHIE2UIR22mpmI+WohDCv1za0DZwfp4vYZwTGNdxuHMweC/ardXUTq
mufcLSjJL7Qvq3o9Cmq33lQW9TYdKugL9m+86x9o+hUIAdUT/PmlTzg/Csixg9KCh6n3bomCpSk8
TADH9UitQM3oFlR219+0P8FiX2+JDg1WtW4FRzlgKqEiAwA9mJ57k1My9zPxo0vGcuDjJnI0T6EH
oMYK4lRBnbIl9hzaj4jFwTO9Qe+bHhU9A8A1z+fdvAHRc1FaQT3htnouhzEmhy9NgdZmOwxEo5Yz
qwKgQZcU/IgtGBxlGDusFDOosytqISGhdVENbGhUWIDx5Nt5Q5T8gIamXtyPdZXSgvA/yKDuJS7m
Ox+rInTv4CX/4JpQQbUeGzmNXwRj/Mv2OkRTZqwpogugzn/R48d+nHCLeLKgkzcnvGhM5C8g6j6o
nuJ+j05GeCNJ/2DPybFtQ2epUttRUpOAvzPXgxPDd8qHNs7nE//Es49wOUp6b9Lu0MEiGe3GIEJ6
fWF3RmMlB8t8udbl0RVe7lktwYnJ8MMBEPn3N/IC0WkEJ8jSGHHCACTqUGw+/LOJP6Wr+2rJ+yLN
rV2HjawidqOsEKx6mr9k8BPze10wuoBC66d2FFlY99cwAv2G+YFMJ0H01UTHu5wynDGg3SLKz0Sw
ODlcngrxSlPnM+t+bHkTc00rG913g9pyrmDFTyspDKJ0JOVvZU0qoKoeCCkK0bkMIX/D1RpA54Uc
FXmQmhaIMoAvTAgqe2kjYboiYQT5jM4PJ3M34oc9NSXj8Wpeu3khkAHhM7JiJp5pCna6aOCfoHkC
l+AErSdtaGxez4UcHNZOybj8IhZM2XapptgI/qYzrsT8XVKWTiN2fQeBZ7x1xm36OQfjGAfoQQKZ
m26HyiWMvRV9q23KhD9RxB8Pb4MLOtCBX1xhOd0WS7g/e3a+V6xa1NLjvb/6GMR1InRq81zZ7DL/
Z1SBp/jcbyESa/PQ4CRZKZwdUunxME6xS85y9XyLplVIizm1O9kcSsHdnvZWngjPgsMUvzS0YXB1
C7QPHzrv1/HwDZbPdvQGbBAkWAIvUA4zmBJoIh/WVwYi8k1jbXsyqCjCgHn8CyFMk4bOtM+TNwHU
pUgmBLNBoYYudPmIE3CqZ/QjIfbPbhJPZEWihJlwF4g5csUgPPY5fpG9a/p1kRV7supzCJcsxHEt
xk3fFxGg2j9wFydqs2i/8VmNxJqXF9eIM2TkoLpVHSo7ac0BXSQAIuHvDchhgCfhRedzNoxH84pL
cTrXS2dmuPXpvUvO8IYdguMO+flXUOGSmM5ugI7Y8fUeepYUlFwrMORvm8AuGTSP3/fKP/j/VK+S
cnXlsnuytw7CeDoZruVwXODT4kifW1Mzo/D6eswxWIgX0iAbQQiwgInfAnFfo6t9OS4J9pgBcfQJ
eVYVnyXjgzodm73lt7iMasARVjV59trlgaSUXHRQAEjRJFf0whpVZlyZ8clapNcTCrjo0P+wlsN5
Bmw3FWVg8hx9frB7haXfhzwlBWCbwJcdwygTO4EXFUnFN9U0yIKBKLr3bFbN+gFDNK5hK+MZypVh
msiGnN7MxV+98ZvuawWj0PagN+NIkCKGzMXuhM82XqEw32p7fW580Gc3+LhaOuy6ACiUmdjRqDPX
DQn0BJlYTH2DSwAKi2nrs+Xt6QqUX1pOEWczJ5mtw8pbYbKD/yImfiHODJaS45ndEGu393XGwGRZ
DrVJusbyRsP1ZOnLQ/HHAfjymepD6wO/ZKuaLo3cS6tPiEvgfCpCaATbZ3+6cL8fT4NA9YyNXQ+3
a3mE+XP7BE5XEf5aZiR9LSeeqdveErtJgK/qF1ClbBnWknn9LDfprg4Xd5WLyi52U/rwg6vpwE0d
RZX6PrVWJv77r4R2gz5rSWLv/upQZu6BCNQV5XF849RH+DLiV5Ko1TvkyRVN2ScFRgc09b2iRXRn
YmivSU1cNbWLOdAjzHPQPYaRz6d0GJSfd0XiOoZkv1ELI3prrxPieIg/DyRW3z+BmHe8nZYBx4yy
vR67uTvooUFXh2WD1TH6tKFeEhmND2Gi264gzQqkcRHkxiRvOlPkxJ8stth4Qr9gIfMv+q2mJw1w
fhw5jNF+F8cmcKFMd1dE9AcKEXAduIqz/DDaNjSDaYzG45SEwJ6NN9yY5suIsXdlmz8Q/4JoQTIJ
Xk0MI6FT7FbBBtY1KylpCjdN6tNf3IxSoObwFw6TcWu9G6s9+GoBW9Dk7t0gXwF/SMLMZOJiq3qW
L7KKH8pus77KOAOrIrAd8+rV/jme7onm7X4Tib9/lpOsNKZ/YbnMSGO1QoreAdbesA/o6v75gUCp
bMsUAfn0KlDObWUSgNW2YU8mLb+wrA3LUVs9sfscN94ux6ChHTgN8+X9fNijlCwhNpFnnYQWu2zI
PoJGZZ+hsBjPomjBUYRBf5XP6kBqg/gvk0nxFPyW5H8uGHNsCjqmwpEPAY+btlh58hcoTbvbiynm
zwIr8XUZlvv3ebPypCBYbanctv5y2GQn/JC6e+w+mL58wERyz4OqWQeIYn3ViEHF2sI1OJ7Q3xRD
uDjUmS5mNkUVCuZnLmeIaohvAYXBm2ahOpOgAdY3lcEsk1wad4PZvSGAJW4iweZhM7FWKIWcuYmq
Mt5khmqXo5yrCONp+H1N1+Jcn6vp2cS1quCtLMPmSKgPX0iD5Hht4FYoFoxAr7nohKn935jkres4
4SIV9p4ktLUyyea4A9d743oKHV7eqhnxMVP3JUm85wWTyp/BpuIj4SvPbPiPT/zscaFubiLLq/yY
sFTFSyo2zmA/pZNaM6X70kmYQBhp7uxP25XOJegBGYUWEB6gG7oaScnEIGFWq5DvW3eaFxpkn+rZ
HbbchGGFS9X+xke2TdfJKphQrXcSpAXjFxUnjMcqa4d4u285IUL9KY5yqZkryYMPWhxubaFDZ5v5
18Cb3xU1wAFHxwOMmntBYz+whAnGiLVlhJwof97gk/pmJhD7ZwygFVaZB1oxDoGcttx98SyaF7Ek
EiJ1c33lvnmwvbwU4rJbfpiB0QcWOAGzRuhPPuPA5BW2lkWDGz0O461YezRi67T4h3Gwc89CjIL9
GeRM1MbpuQfkeLzeD7wAxLcdeQgtQ9YSBfIP5skUcYUM2N80Tv9ulrCVGcqeeH6qLpjZ3NDKwEfp
wcZaOKOxDybf9eaXN+97amRgSp5nDJjBCg7dA9oGPLRL2OcL3bS+4Z5rwMbydn85ezZImrjpYUPr
JF5f+4J/nNCexmEQYD9MABTN+nAVw2IRsIwnJguq0lNNAJDExJGDAKF2U39Cig5N0o3rRqP23p3+
qbKKZxRzHAp1pHsWpvbP/B12d1/GqJkwzxEe6NbstvS20VQlX4vd3RXRriTYVhSh7yLETXDpf/tl
sGb7m2y1eKqNfVWsX1Qf1FmiJGpHWBMQmTbJQ1FU3r7O8ZQzmaw1vxGV7vlW0uDSHsoliLSUAmLm
ZQ7893K5wqdic3HC5iVEBXoYmzQVn5la1vppyPpBfAWeZogTYHjzjmnMN/sN/OxdqlKAcXWXFf8i
0k7dVBwAapjJ+eLoxALbZT7K2442mrxKetmKSilqIId/OvER7neswAYoSTE4bFQViGcWy2o2EV8x
J1AopfEFkotItF61GbXoK9f875qpEqxj2WwAwKYIGz5pj8OmCqeEETb1sJMEQ5UkSOWc1lalNCBS
Wl0IOL0KphZt57H4LSt2FzagogzcWIV+csqTb05kW4q/yKGTjntmeVf4mcF9dg0yARwhkYnnUvNs
VulXRcvz/RZZAJ3EXWvSAa1Og2tDawMi5SoX4Zq2ygyiYRLm6FB9h6VlO5VQF3v5xY8muIFNH23g
dIqm0WYCA7TGnU3jEpX/YikNhBd7c0khZTUEhnLuD2xzb85VU0vQ+ynSIEKPwyj6nX/LxDntxVb/
lOzdEYJEnCa88hX4FzU1gAwq5baUyi89/DypEJBlQdmglSooskTxCO6l7K6At90GzKcXSI5E4Ivk
TY9kNo8k7DNFzcPUkVnex3cwc4E46WefCGHga+bPzVBjRGvB4E/WGO6oZ4uKdAb2ENFGFodzAtVl
neg1Kd+g0tQAMH5nZYTaFE+VqZE+mXm1V3rspUvZ7R0CYFAEqL38CJ8twjnHlc1KCMgRYFDqoRpz
DOZtEVaG9Ss8EoKZbj5Z8PCJhkUfCFkuQ7Ot/J3/tlO/WfxdEBBot6z99ss5vs2J3Kfmi9M90d4y
gA8DDcDNHcvjayl7kcvFUScqa5ZFLU2N1DdC/Aker4tseSzTt8nHxwG7eskPcKOg63XmV4m+yPc/
sWwW/jh0lS7SGYFmNM8CHvZSQeAVTAnO/K3g0c4AnUIhU3PjQfecwZW3G0co0pu2mY6INdbf4ukp
6edtHYaEpGri0tNH9QxsgtP095NUOUs5LzQxFyFdl+/RenPYm98qVmMsPslCgrFXRS6R0tDihzVm
WkXrsPjyzphZ7sM8vfShuq9v9v5umpzxrUWjqWx1S7dXDqSqCjV8zeZysil2AWBdPZfVNHCYtn+o
M50cr5G/84Mp8ieaFPZfVYg3TrRJZ1DcVQXzz4YisjlXZzkPsqO13dgydhRoDSAnBRuMa/u7g+R4
keIaD8r0cJJbdeuEYfsqdWMVpU59rT3HygrXEqqrzZAWiacpXeYJc59WOa8wuXcScxL12PvVb0MP
w2noBIVv05opSoE50NnQXgUPgdvjt7IeQK8leqs0zA0cevmFR6IsQKXV3OIoxuynupzsBVIL4g0X
Ea2HcUjOEO49/sqd7+auwLx1yEAu89QVFwGjkeCduWObuD2thVbYtwtBtOzDEPWEBTPQftU0jTtK
Bn8IHkTZt/OVaRMks/JpR8NM5TU2u9hJrY9Z3RsSdowjxJxznzzGfrC1rwhnwgh7/iA4xkSlHsxa
u+pq3olWBlOrZgZZEHwxWIVg/5diGFoXTuvcu9KuWtZhtOjGoXbxfMvzN3yyxKKV++GpUFIgjKE/
qaMQ9XAgstOxIJBKgq6TUgZD/qzn+dp3maUcolO0E+DAnNnAxSEjNryxP+sk3yW1o3gt8QeDOkfz
84Cv0ZUocWhgPqQYyShN4zz4suqIZhEs4O8Ry1Ok+bIo1cfbV8+5xHuVpYaiqKBQ/Sp90xW59spP
MX6hf4/tTs8qTgDzrfEilYFiep7pB/uRewxPeBzG7Q1urW3hebDHmAplae9FpIoOfEN71gNfHAIS
pF2XM5Ayg3oMeQq99F+7DXwMw1z5xjn0IQIbrixlkdrEWyj8Lz2OVTPPGKREsWKBJCsby12cY17G
c33WTlE6G5828W/Be7GOLE40cd3URAdVx4Yu+5Q2M7/ZXJiuwFaC0ujZtWX3XMJ3l+N6Xgo3cbik
DZqXoL6f4VMABFjkGTQiJW73gJkxUrtVAMV64yV04o7VYFueAKYTTjhO4+t2HF8ZwWE8SI3Qfwro
sU9qg6Qiy/R6owKGj60L8FZK0xIIUtAHyoVKDofZkzwYi6yDbxpaVtueZZ600OLFR45KflTASqV5
ayL0/hpSNNJTGmuvQeXnhK8TeoMEwhZBgD7UZLyrOmCa1i8d9adWnEX4dh9QHGNnef6cuC4gQRJM
mJ626wR4njXr72Szb/jP2ftIThMARtZvdWY/WSvTmwQsqKbkwBJLaRWtdzsO3uIE1aCD8yE+RJF8
2m8J6v/AJpAXN5ivoryZezETbb0IyYXekMs5ZBTFQw7qTVcKTMijdLi7pNcZxj+nFS5j2UXFwZ5x
RMl9EtHmhDZWck82M4kkzb03gvd05Uxqi/9lNJjtr4YLr0WC4vuLTnZiIOyyZm5bRMTp8cYOuE1Y
B4gsItQrV519/zBAO8XCERyMexjzLm1zqRX5y2cGwfKjx9pRUdtPfvXHz3AvRypRAMG40A5PBEWf
CJNCKf4W/uRHyduaXvw6Nx+Oqe/UWEOkEXSghFqEUAqGyPTplPHOa7zCbkUqDBh4JsdjldRUbvWF
rayq78ZvNKZqv3EwI6YRk21beJCnjmxQGyitTkJGB6509CRTJO92ScgfJa+UTKmWgPEJCzoyB2+9
vgw3DMDyeH65lOgNnPhzGPtxun4Y3ZsduTP5TDWuJVvDrhbqLY5+n2lhY8DhwjXHxOzzeDNAQ8lN
t2v1r2axeFuzCqQJ7YaLUOEz8/B8QmsbhqvikDj0r8EPj6FNpDVdDXJ+kWGiHAHpmZ6iU5FxfNvN
zS0MCrRBZ+f1fhgMl0bscW/lE16qYyJuJ+AQwojdjRmdEw/bAtjTkEpTHsgYvhirM3OG72DJNAom
KE38gmm0HMSUpMq2TmYU/mvgswWC5rT552WsqbkbxL9XsFLBA5A04oRnZD/86sUxl+BXD0jE0AMJ
YalZrv1uh2/oWb/2OO1NOk+A48RUAODfkJlPCevbFxdMCmamHRsfLv1JUojbCDjPD2aI+WqGs1GT
dwbuk44iDUxUOVthcSlR7eABmjGK/CnLKObqMj51wZw1p0V2JRZBuidc0nSH1CdrVkA6tH36ffq1
KrjWUE4OYV11HXTYelu8w7Dg0TvDNGFQNqx7DCgteheABjZb690xiWPNNHYE9zyEMFuiLe/gsoFE
Y9jSJLIB8c5ZI7GnxlIq6i7leUGJeBWXdNhcFja80uUcJrLc7Ksn+laAIMiE2S+PZQwZ3iDKkJsW
Cojpyof/Z/d3h0/9IJNAtS5PX52ho8tXuH5YPsNurKsfUEX/l/5Ky1zX+nxEDqU1mqmtFEipvOuv
PwqlXuRUOM7gwh0RilQeitkXAtp/0n6vEnu6iaRAu9YkBb9DrpxO3dPrJyCELNZnEqwfYuccmPTp
SZFkxvSRye+V3C+LisWLshISNoiT2lWW6P86dRD23L6qym1fvvBoa/PKYaicSez6QhtFSPGXPe7T
VdS2U/TJC08ngF0N6aiMAyD7oJ3AKdWOdFTRLxDSCXhUS5ZD0iyNPhKDzRUtf2k11VotY5jDwLLX
ltGrlr+T7p1yRrzGxLPRSZei9E7+FYPwS3FCLfdB5+mlVEUQqmkXRqMbneM9SICZ1NnvSMuGh0C+
EHjkWxQajk8N6g8CXKRS1rFItOwuJk1HURstBhpK9Lv2ahtQWsVAyVgkxzajDukdHP1dwvVhFg+2
BRhzgUpMQ+skn8xdWKBOmh/kNkTucCww2NLIqJQk/BrzuUm5uqfjey7PB/YKkTHFR3GJ6JpufRIk
g0WKftuBt0XnmmhPKfXmG7ll0JQDfGXYztPiKzMA2bzo9mQIoyJKvtL3gCgO//5c63++ODQoHzwG
i8ex5NOeA2ttqsYvaEK7lhMoNAsoPKQ86Hwz432i5Jaq56+lOXWWYnUT/7Aprb/jhGG1ZNfMhj/B
MMz+LRIEj4f8YewUp7kT5XbNYAUK5XIuFYiTsrMj3edK/eeaAnIALNWlSmlyRdij6HdQYIt4957Z
tZSs1qU4tcJ3r7zvRcnz2pI1mYlvqrApKZPjMvZrCE7KATohbxtqCAIip35QZsHNkqTKkIWpizDN
44gPV7bZeNMM8iRc0rfe9Agvs9qYxFgsNSDUqN0SCWpfduVegEN/T3nUG8YtShT/TAgVi5DSlEZS
kp+U4x8E+pGMj8Z/B/w5GywUod1O+2dP6WRROznGQP1Jdch3OvOirFBqh4QW4zITLYlVcRsn5rl0
IbwaEYLsAcA3euBkAQo06YjjyTn/xPMVWh2WqBGuR8vr6I+25rTFGBoq6pTh1fZt+iWVc0GKBWbY
n3+RQPuS3LrgWkviDFxL7SLfCAyTFYFw3TPPy+QNvPIOqOyJA2jJ/rgWCmp6Ted2PRAP4ULR3leW
Zynm/oQwda8cbgnLZeTwno9ZtjZV/9Sj04cIz7z+GitqDb7tIv3LeVPCTVKhbMtZCbJyhKE1dgYM
VLTPVnHmXueZb+ZkcMmsPhvbV6tZI3FvW8pMOS5DCSag5hC39pvppWzOAOSOkVHca01gQcFxUTAB
nOx6jWKfDzPH0qPQrE3VA/38uCsIZWiFxacTU6szUpmvpr9vPdfsXr5n9NCc5IBIROwmrkkD4dlk
E7fEJyrBVb3Hmt7Mq15s3KXc89tCstArlMKRCHOMloH3qhjBmJDElE4eErEBE2kpLiynGBFhS9OW
D1GBe391X5GYUFMXWVd5CN/snXXnrw8Zho0Xvrh932H6VQ+HlrMmKc+I8YUWPoLB2Z0/OZrdxrd5
SosRvJiFvRyfjZIYFcD0npjygyn3YSwQXaHoiIGq5/Q5umXb+F98AgFuXfV8TbEKZRpBe/+ZXJtM
txq9vh+n0O3Dv/dVqODIga4b6fYmIc84aA5FaiCmaDeWLpn7vb79aqBT0dN6sKfkpD0iQEW+xeeB
1WFGA5hY15Zn4YCH39br6tmqVaNnPbj0MtvuGkxUG14m3HoORofyIBE1htqRo8KnGjsGEl8q3vTj
uTv7yfaT8ZrZ+oiCLMgwW7zyAe7EIMxWK1YaFGLbWpWsXpETWq0nAdRNE1lWip9+7brJI85XjZb/
PtzQ9iPitzj2ygpHGQGPys9d+/+3x4FyEiJPDNhE97Wc9WLlp6JUQ3cx6TnxjC1isbzyrsCLLuOb
glhNupxct0kblTJXpgWsO4d6ISfE2BlPgAqlE5iV7IDFFDcu9ig+4k5w6Qqa9niHKcSNEs8BHVVv
PYzKHa2MpHHhO/sITcDqI9ehurpEbogRuaaN3+2DyqSj8WvB1t5OFNm/JDvqPwhzFtz1Yb3oJvuQ
AfrUuJ9yJOgIL0Yxc4lZRrtgS+4egWK7N6oKnbGhc/SZ3rQhb07H+Pku5EN9X1NJaNcTh5ReL2g0
mA/kRrdIJfv1z3/n2nBjE780eWAZdByQPje/6cYIRTyRFh8PzkfHkHoqQmGPFQco7hRCeNO/rZNS
+3XsuYi+9/QVUMmfXCMrebe4zKMMVxcNF2+0w35cHaK9gArq+43P0reB1zt/3ekkZNabYOV2KauH
qwIQy9FoaddsvVAe+kv/XT+rxOVN1LVDQY4NEst2nnITMWKSh2uo8UKVE7UM4wIhEALI4QJFu3v7
KVUUhZoUrtz8I5gUU/LXzlxxsfShBuVv8puikyvx6+CZBFV60UGzNVVYOOWeThuUKLkaP171G0zG
w3licgW8CmFyt5G2rUMxP4i+qPYiECb7br14T6K4UeQPr5x3ruWlv6SNoDFUZ6TNUakbxntY/yqm
eaSPbI/rCxFhBrJEeM84lU1Fp78V70OM9e6phebkkqr33UEAJ4XGzx+gihJpefrlcKkbAR12RM2Z
dFDvDzwetQsbbmsMLcpKO6Dhih1g4NLlXsmD0JAyhzJNnfRdlyP5OxwODls3qMOjuxVhGL6+03Ts
UxCqksqRtSGNLoWY6w8CyeQ5uc0kxFbvTwYFZwMJcv/XLqNGA3Ch1jT8wrjwqAFkM9umaoIuzmVw
2kCJbs6enqthfG8HFs4yZ2otrk5V3E4ohRzlBoKwrw2cjQNszve9BtjpQx7IpK9g1n9LCX8dHiDA
PCHR6wspgr3sQ2mrbNsg/xcDzSitOzVw4Sa5NstkpA5JSyVO29mm2dFZ8wzFBB+M/ZB/NhhMJmA+
ieWBTGw9h7L/2hRNCXc/EA8iyPG+rJSjaHgSr8VIo90/T6AqAtXDdV9nvh9UigkOjxLPS05SJlmj
IAWfxX1JZz2JZuKNU6zLiGeDGxcPBDQStd3tm07K777pkwEfe03IAF0arsxjxiSzS+WFdQaoV/Jg
v3XFdo/H+IgEkhSheVYkM9CXKAlYAYl04oPSjKef/MEieeriVJPKmkF1/xn9iL/sXQ6bAu8mLmE0
8QHxPlM16+Xsw29zLHiK+Sa0kNpCTDsqN7w8p0sCkyNFYiPmzhdJuMNVou6bCF0a0jt1k4ALCmsp
qzdZ5mON4N2LTnksSGb4O07jWFLaiMcoJ0INHyKiyBKNrKDd3nGar1We/KD3fmdepd2y1Xy+2pbS
t6B5cghGNds8AmMKpWnIg0TF4ivuP+oukmy0sJnxxLxWljOTKx6LatXhgaV/OAYPmFz2ovzlhaoz
w/iKoNxSrFQW5tlzUmp9NmPNaw30ggrNnl0atFahjChYzKZcGPOnlBt8xYf461TzMxAPDTfHS4Wf
2AGIxCHod9DIVDdo5Dk1bQEXx5Q9PatNAMUtDy+RJsVJx6X5nQwT/A/KIx6ZPGQIZ9Kgde3uDFIz
ArgX7uP8P2+Kwb1UD1aCZNyxryi4e+OQzTgUrDV0MWD5nbPRUgjGEd73lwH44bEM9Exi/7gDJl4S
C4Vk0JU+0KvBeVidNT6GNIhVAvUiIPJ2OYzUAbkRZRlT8waP5SBSOVYK3pcMCo2uHdx11+eQ60Ue
/UZew0/tVh3IQuIjLy+G3oYURYEDfM32oPP76iSkyRkSIcii0Jqt3L2ndqXwKPNpQbcOtnk31BUx
vosFmp0/Pq5F0sxERbIg0VEA1KO+UViE30KBYu6iL1rkIwX2j+eh9+5zdQRpKhaHdGaNaPk4vtS6
0+/lb5mi/0KqltiaGdeZBBuXAck6KRdw30/MOOFz37ucTStUaFkxyEOYyIuQZdFjzh6HHeq+h7tQ
PC0mi45GzMKdvCCS3qdxVYKllgNM9bZrLUncmOdab+y8nJABywHXUxF+Dc/9+8Xsa5LubkOXcquZ
kxNRRwMd9MJmetJSVSAvVFmAcTrGQdiUjwzPAR7c7FNrSacnoHcDg2IdiqXyLGst3SMiGU27FYD3
4Jnjej1yplXzWXXZbde0DSCBJU5GUyNedVLrV7q9d0A62zR1CYNqkk73bCileuhVyUz/m7wrXSu7
NVw03QqyMR3HM8a2CDvmDxrsir9hwFnaZLs1HWrOpL/ON1TB7N+fZzrV7U9WaXRmEY24B4KdzLLN
lspsWncON/L0qlfFMQ/ODmO2HiU6L6S9p2ibBW0NIc9d1p6TIEjgznJIqKp4VT7l+PcQWX5mQULj
UZ794jhXdtXAY+lNOx68QcluRBlUsxe1cq+dTCAn7lVxOCDb3dMM8eaaCjMm0tkyLyxhmmMkWyY2
oh0fIfWiuKLvuh3kTpK7dMN5v1jAtMxgzvNjYUQHNFESaYuoWtwczjhlP4lA/eFDfh0cdKB4xY4A
NgddFkVhAgBtuWTNVBXpRhaDzSjvVNfpSDXKPX97gNb/QxiGwXbfw4CFeO78hjiJzV6kNwT9rm7J
2ZxTzDk491b1QQbqqtwa6GfKa4QK7mjtMelBE2192++k2WNbRvZ2H2xwkt2/kUhYVbgkJGTPGUjP
5QJbRkI5Ov3OIkn7dKm0Q71zAR3RjAMLi3ysglR12Opbn2Fj4sQFdqSzylPqFglaOcFnrM8OFrP1
TXe1ptqbO5XaIS2Op7lqw4dA6fh4EQqyJZMNyKjqPojCqGdmlLBWD0yiZl565jh5rKZULz+Tr6yf
4JnueE4XI9L2MKZxWpzzhg9CaMfP6eib/fEjYUoERfw0+TJ5pqbfj4qR7TEeYyxWhyLO9Ra+cbOh
zwSJlBGq3+s96Lvm7KIjC4FTMeaNHZ9+VxLBi1qVLUiAGDWt104bjKT9vvRyFus2wS0qPPc1O8P0
uE41vlD6762ofsxNlEgKRiWwL1zMMXn1RUCsMCxyO4Nv5u2K9OeicylQedQXsPSPOx3SwEJiSeYp
3Cg6EgjxBZ+LiBYhPN2l2arDz2KAoY/CpByEf74bmSRD9w4o1q/VTfFlLxkhBFoz2wZ1sUoX34yP
LNqALdz+VBYHakRrenqlOP/0sb/ngbTfcMi8HnVpxQo3P4gNtInrw/8ewbFr5YdwIyuNEISqQac3
XCawrNLW88dgf3b5hqMzgXzqavJZTvbKMqOXCASLk4JwHMcrDPMCNZ8D/t1ootcn6fM37p6Fm5Mf
sCm7fQwlaLRGnK9YJG/FAryLa1nKcV5yyBL5YKyA/jDOYMWM3dq/fJ2vShEMYRCnoRooGgDlqMf6
VJt4OQw+c85d9hXQyZA0EJrGGBq1Foy8pwQKTaZxovkxyp0Iach6Y1S7vRLKX2ilE+ZD8DIr4iOY
O8wJ4FhWeXkMoDn52j0HqmtFoH7EXrqYYnJTzDmvHNpqQXyy8Suozbn0Yh/wwarF8Z5yImNJLC7J
PotQbV6sw1LOfDyljFi8SuttKyjilpdlHy2XHkhM5zUg3FSIkDYrSzAl+HxJWdWj2hDNgk58rXrI
NOoTtSzMw5c2z/5RBvn6Nf/moclhnLT2WdYtS2a4IITgLuE9UFslc7/aj6KZ1FBBBxk7tHnDt2Aj
+9bsMDrtuBQFDLPwaUNIOV+u6dDXQz/pQhGvAA7KHQPiE1em4ULmeNEEzZGW9tloKlEzoqzd7CsL
p2ltEijlnDQ4QXxgY+silo1u1h0qnBZBjpSMVmki0aV1XI6RY/tljAeww2SeJkxPZoAHAID5KffJ
dEksL9hG0kOuQpPZZRKMsGYkY03s+UiEga4pkA9BQvEmHadHHX5oL8v6nb6z29NNvu0qPpE4fRD4
OQl/7/7H+BdG0hgxY+/iElfpOabpmX2LUGN0sSD0AgUXHvuDrsJUK2akmb6BR3PHuV02gV2/+Zje
H6Ck1NJWV+Ld4l04Tyi1tvtGlm9i0b1Gbt92dIXFoZr0s6hQvuCEzoNgrQdjSiNil9mzriQb6P2D
o2hyc4H24MNq+v95/jLqGrz948+uCQrDHw24jhE2y7rrDfnvuK2slqJcd4fprQ5tI5dvNa93rZKS
ejblv8LvcPG0CQgfbag//ig4h6NE0aHGJ6rvQrmoKqBeOer1SUjnPc7ZcXtcacVPpz2d2tLSzjSR
eQDvPhuf/jC8/DMrNRgpbTeHf3Vh8vk7v0G2qOVHEhVVQLdZnKbK0ZgXyVXQdl+wNGhUgHUTsgbF
o+zUfRzB9zxJalaTQnJD8026fOaQC2LgBPcMFn5GZaqg7tUNrFF2Y6KnF2cLfvPOt63zY7XadW8D
ErWdSVgqISKhVe4Rc4oyV56MHzPheojDSSqu/CkMMYK4UM0ZAtNUrBkyJt3c4aBQqathCzjFfXAD
SrzYV5iWoJBqDpMCmxfWFF/3BsJCZgt47uOoW0/26boak5wl+wwi72FdFqSKL/hi38LkO+rZKKmO
+9VZkXFzb1QXHU7As7vyNq552VVnNKuVNvOibGp/QAb9buklijzxOYe7Fw+4xalZFOSRumBoBjRm
URA2O3Usr2kEqGd3qZzqQjeRA+rfBVckIPE9a88hYSPx5403fQfvqoHK8DXXDH78PcjbhxdBOsXE
XHxswQGUh1WLmPh8GsUO/AXVHyp6V0Wq+dHNucGjGzupKrgdVDi7B3NPGHHdDOxiBRxeXyfIgLit
qxuOjJz1JX/mHDT0Zr2Vkn5/V8H4zZYLflAUfYtSs33poqppKH25IWQ9C9ZYyaecoRSErXQ8F0Dn
zSHQwctl6bMxkifbt49iYfCdMxEntU8W1iuvEi+Pmx6UaO8ok1zgAfjKq/zUdRWnG/D/u2cRXH3w
RRMoN1zEDOHI704ePHdU+sNx3fz2zf8J977A4s0AX0xN2KsGo6PBl5Ezi2LkfOLV2RMK150CWFxX
KKfq/CDcTddlM/hzyhxjVIIKREvSRYdPnYSIkfzS88QFjZ+dT8fv/7QcB3AxKqfj7mIHJulM983/
+H94zWIvqfUNMJLHBQhREdawre1M0RWMyjTq1TMZ3GxDv/NRyDNOyxs2x2B2w9YVlK/wPU85097n
r7czhpb0TxSdmrdKTGxQA70IfiTEROtVAgz+9/pFul2YG9r+FDZBHHFugj42CyI/8g3JxJlpUt/3
BVuDOw/NHNjSMbnfJZYTMEMV1sXxzD9Xz8SvZ4dI6W1ZsAEdUTj/sC0gEoLKew0OHDIF6IB5UNFy
wRJEMi5xm03LuM+y4GtWgJg5OsFBgU5TumOT3Qp4P+TPA00Lc2yXgf3n9IumPH7lhyam7c/a7iHc
WAY9tIXQHvsj7fwpEsi6q1ZYM+XuqY9xJz/v4VROGpinLRlHSst1uMggIUv/CP1aztRNrK+R6ReV
BOhjwa3r+faEti7PN0cUpxGhEOQODdeZS1wGSmMQzp0K/u7LZo93PGBgPdC06Ht+CCUz2Kehc3e2
GlppXCIU0/ZvMNvNHfJq4HxInVQRLCWE7N/x8DXgPlKQyxiuiUmu2uo+NxWRfzhGaNpQDBqci9Op
SVT+lRFl1hrpjwXGBRD36iPUv+I7MzD7Kq5QoxL3XJQdcAOLV5n4tB7QWSxCd89cGrEXqgTPGPlZ
fPGoWr7KwN8w9Rc5H6rZfnUA991C4VYrd+d6FDn4hTk5+WD1bj0Rpdc1A9SrhELdQrd2hGQ/1a3P
kU2JTyZLh/iDTF61DFjkK/akN2FugFSdc01fH+Razd4xbUsS35dBBelhDlTZBp94Q6agcLppk4cP
WrtoobiXL/Sq/He2kQzErLeqv6mPNsrwC+YmeUZBj3EMUvo3WOpZb95XpVYq7+qJvx+nPQTiHqZN
Az7E8A1DGMLjzYby4I0sVh1q33QwiLKeVzHWYWe54uxnonzAhPcPNNe0lUY67Rq0h0J07EV7LWgN
jIu1hV+9nUHQkvuMmxDPyoJzXV7UC7L8AK4Bm4q8VHYAi/MAw/DphS8EiIoz3j9WeXvSPh8nbL38
I4BDvL+jJdGWJ7RUJWcix2tBgL281z/IaiYjvTOabRz6g7VFCBO3b4sOIGxKXM4WqZ6jkcbdB5dP
nU3Zvvcqp/KrGlB2Ah2hisqPYhwo31XnaW91fCsXW6IRIW1DpJ6g1NBAUXu4cZvFwMITIFcw28Lj
xKlkMzD1Z9+92RLEfwRxFVFoTP9YCgkbQQJAmgD0zeToHk9YSNoxfIfJU9dQrcaQBIqATpZQTqgu
CTwFlLPBRf4bh9NZDE3LQ6JEeUWNlWPUF/xtdVdy6jpx1QC5BfswSr0FZ73MjfPvcNbfZfU3JlnU
XBfNQucdpse8oO9EL4ytr5f9y8VV+FSblzGKFIunLVPKjgfZV9tHyXuH1MkZbCLr/vLH01IowyV5
GZ0CRXr/iScYdIVGFtjW2K7/l6wUE70P1VsMBXPGTIP6i7rCNiDNGoOyN9h2Ap3UlEe/SuSusTQG
3SOLxK/moDdYV01ucb09uGWCrUTxzPLvEcN983Wri0Ns8B/iv2QYiM5IuktvoNkuiM/IiLNkk57Y
B81TUwdYSf4RLtvuiFUlKmOyRVZwV3RtJRGrCWDjhQULOlQcPywgb71ciYqrDOjc5w/ZCvM0PsL4
VfRFp3rMjDnsG1RhGRGMO2tR/nYe9rSW2gnULzlDOmoXVdBJ7FSFOLyOZ/Y5p8i0jMpSEpqtGIbF
c3MPzfF9LZ3zT0AIiCag2O/DIC0I5ZnkipNDToJvANa1PB1T92Rg+aCpkD8DG7r1awFMNM3ghrTq
qJBubWJVToAA1miZpbQlCVpMtK1b0UFjeimSjT/yioLhB4qsaAmE7RrCOaTEF6plAe/1kOst/sr7
3XkPi5AFeI+5CLBglYIvXW62sFt6S6YAU9NxLq9I3Cp+ZaVC/VOeSr21x33gOSDfh2RbMDPY+kjC
WqjPOpItX4zQfPePnYQKesgaeN7U1b3CrYZfXre85R/iTXPnU1n6cBzMizWCl35c6IyUMVRXcsGh
Zbq42kKNh+pQ50kzxfVEqjQnjM0K+xydVJzoPGTd497TldwW7ofxxG0Q3FMpOOexPGqVnAsxc4yu
kZyI7W9s4Ej1vZA/L0Cf5APoCjVkuaSShkX01kgt3xg2aV8e+3oAWKFu1ryflytoAifes7gfqT5d
/uF9FE1cfoCCLoNB0YHl3IMHJgr1p2TWJtgAO0uTR4ZbQvClDF36S2h8qPKcko5I9ekc4fOGBKEK
Cnof39Ri140CXD6jpuWWmBX8GRAqgfV085zJ6QXcQHjoSmD/Go3pbSH7PzLXrquh2ut/eWZHnfJ9
1GC75hy6ymA04kagROcxxKG6+/Zev9ycS82AFcEB6Awf8xZ4d/fDZj6Ch52nwrXCsENk6QturHYz
YMyBoZuNm20cp2oCDk/I2PP+6LWRMHB3DxZNeoHJmUybls8Z9iBiEuSvpZi9J3k54O2GNsNVumO3
CVqv5pErzmdEUF+xIeBm+mAOYqQwpTkPsUqEjMWHH/NJdSPU36qY0iaLBc0UUUMba55gyfZOZGti
Pm7oBJCHeMl7QoqcRaV0L3kUz2Ai3cmgxROFqKKlPOUUTOoKuDHCFyQRgndXk23KQiXQ2WKfk0xt
MbLHgCMmU7TgTkBAxyQWyWFvsjW2HjXDN1KgCZ9lPkANNVkT18Ky8kxAe9vPlrIg4+N4lYR+laKI
vjDMgr7pVunfnuCS+VwZJCwqk2A4qgEniobPsCv3tzeyrn/ecSd63xw9C0xgLzQW8f4Yz7+dsuvc
zgjvHbwHwSSto44KzdlhLZ1x0hpp7rAUXAzMrIYh5JPf7ND+hpkE9xACl/SQyRQoBjV1cTtbqMd8
6JKqL6QZlJeWiHOGlWNKXcpKasiWsOqDR++xf0pvbP+WQwQA0SudmA5PV4lJIf4jjelR0fhR0OTy
Gg18GPnjbytX9Svnm3/Z5uxvC6eKLfzlXJFD/5bhw6s+q+3AsH7YJuqfV6QT2HNVHFWpZpDkWAEz
ZYTQdgTeHFIt+9wAJecgA1kidzeHzia1X0cXo7G5mzMRQySwiNyacJorrh8FXwGI0Hu7gptlp5xA
fzaWRsxh3/oJEGnpJQxDuIxN8FX0nZRckvRsFdoEZQOXG01YDnflF5h9tsWTslL7luR5Mtv8Rc7w
ETkmftdHylZgIjqZkZ1QJuMbuK8KWFCMipKVSMR2FNEItLDX64yN5hsPZeYhLnMLk4nSM+1TNatn
qitxAH/g7GTFy6G1qB3efuUyKJFhXPcoxFf1+SzSf9WWh1BtrbttktKB+V42lPGHkZqZ3KDAN/7q
fdNiZ0mrxYyCUJ97GsuF5I/XXwQNFi1uG4Zb9OccWjazxJAA6NXFX4qavomcyjHU71O0tMFfNY0K
iaYvGJBMKbXYMf/05zzGdeloOz/3KIzIc/GA1OqRx1n8bK4OC9JAXmSOUwBEGODtULtlZTi+11ap
D0XSQ+48lRzQYijvIiKUgplRBz5/hCHpfOHut8xyvnZrohStfjmuw7EXD+wkz4w8GQlRxIXx2N39
emkusa9uCP6Kw3T4EjsblpzKtybtc+5W8WBEImEu5nXc+/hos8NEU50hwtzTparvBlnoQfbygGt+
o/nBCr90k5J0ddSb1TruYs2GOZsA89Kysb0QKPXg/URvspXIkax/lmXKUWCO8s09RQ/TLTvESANa
Q3q6RH0aBWT2ZJLy10gyYq6X4KgweSrI7iV/vbhMVg6er00/YXnB6dhqAXvs7vOMT7uJ6XiihrvG
8VEOZfF4bPXaT2dtIk/0oO3UCUNNX5XkG6xTv62OmzH+SzvSsvMZAOiQNZJWOXOg6XhKy1AmlnnT
dRirvxCiGl0WIXiHSQrS7GmN5OSaSKRZap559K1JJPaZmcLrpQJtj5qPmZQvyQwyyWTdxHj3b52+
oKfEVfV6lAjdUYDhIZ67uH4JhlwHl9rVrmRy05Nmq4lYOpGtPJLq1SuQbQAbrqEkHLBm3U/HkbQ6
bXkhbFoKwG8VpQbqHcPYVnlgaRbIfUPCzNf87ND3lSn5fuyxSIWuHRKHTEiLDfFWWMoYDabuJAyp
X83tLi+SNzUs/iFN8LJWsSGtGqaIACalEZgGN+rEJw/G9RorzbRU55nCrsMs1Bh1Iok0fPAT0yLb
ZeJmr9MtsYiu6Ttsxa/2REsbtCGDWg+SuAYzQBwlAydU9KZsxFM6adUq56uSGZ6tV1131A6i+MlQ
0RND1D404dF4EyxueGNOoq/6j+ki8z4GU8KLxSVa6m9tyJDwTD06Sk5BLvUsF1vTLF7GbPiob8iK
+c359nVP9MIkEo3xx4szvMkbxigovBdPIsiGvh2xQRw0v7ONY3trq1o9QI1B/yPXSF4f6bQVCRaJ
TMnljzVIeZFFODz32qY4CsZh9LpcJtKVnWCmi1cLL6rmORWgIbCqT5xlB1Kb9vTj2sUcvRkA/KWj
SRnAH69X2S300MWO2WuemOxSBQtT9QTsv/A79jSYqbMmy+YVzrpns99gSEeo6qY2Zo7IbEnA6hxN
SNfU3YnFG8mIYkGYydJaRThxg2UuFBI6GQ30ybzZAlMJX8Ab6pwuudeGNi3rfG2Q5UZYIU/Swp4K
z6r9cfNX5EYUYlMzfQ8XFOoE7WsJPJ0cRQjU3ZmPHFhcMYx95N80CyOyfhgazwPKjC086+eNYkEg
DZ14QJkppabieYq3vG8TfmPZk+zt6AiOGbjIuH98a2r6oWjW5wI9Og9cvzF4Z3dIvYTE0FWU662m
HOctNrCn7Tds/1NV5KKmoVm/rRQKcycmvdWT6NMtXmDjwFZSExc9H54pWA+/ShjKJ8/hOpA/77Bx
QPiyXpoakb5ROzL2V+pxOVBCjEwk0DwZ7l6txD0WKCHgYs/4YHhmpSYj1+SMYzXH8ZL8QsSejsGN
ZTeKe/Ez+ncixXLfBzLw8Ajzv25eDPW4SBdwvD+GPmhpagOJkvSnCAafgUOUjUbYpAK4MlBZHw6a
FSxGnHGWSJO1IBR4STHrn6NardPmUnDwVEUaectNI6N1NNHzZT8HmuQX+IZ1E0l7Hcq/TI/omMba
39Rn4c5p/fSqNXOxFrQrJ/Qo974XZdZYbVO05spl2rwGZX+mFBxlKO8bH9O7DoWip1ndXjY0neQ2
H/iyIKWZKCdwTfXEvx+/NjGmmc/d+4d5HxV5O6GxOg1gGmBx0aX4YVTYKxiEB111+pg1Pa5JlaZF
J1FJz/Nv5zNjuNVQcQ2BhxrwZ+GgttHqJHY2I7UCg2xArax46nyhBxiGWGrDG1IwQ9ppoZNjWWl+
aIeXoYb1tZrlG1M3sYMqYTbR+wKeUYMyDWvV6rvZNgz5jsvZekgDmuY9lbBxwy31p1+6iGlCq2nc
IlO3y630+2YPi7LK+669iCIrrObVb23klU2PRuIyFa5/EmDrBSMyrx3j9C17Hml0/hPmmswUHZCd
ZisoTZb2PlFD2Mv0CNK5ynn1uMG1+DQw/onQVyGGxVAH+4Flp5pGUQdxEqKNYBtL86aqCSbXLpbQ
bMM5TM2Dx8HQ+6hdCftKZpOLXhzZmndPdEtbPgjhAW13T3sQx9HORybPkF837ZFPcro2oW4M/UXB
1Lw6hc04JQ8CKgll9h25NupPzJMnIBAH5vN3y9WcoRm296nm/2JBED6HABqf29bGQ3GIQu9CKrZJ
Wncqwm6e21aFRoz0bv5ySuQhKlGPH63jdVMRYTNPtu8iIXGV57VxRN/5tWBuR2jHOShd/GY4By2Y
QWndR6QDH6o/Cup0/rVYWApomy71s/cGxitVLdHYfWTlnXCnX4aGZHWTnV8U1J2aE6l+XmchueLp
gNiF3TbDXAOySYg3o1HEXs3LhYrm1j+0dWarMMq16kQ6F8EvflcdoyLFFgzpgKgLM+nNY/S6jJbQ
dxlU2/ECbJEhRvg3nevA7l1F0eF3g7JqoS0FYUtBRmOIqNyMccl+d+KtqwoXQMy9CVGaRt4GWJTH
v2WX6PyzFotyfuqEC3zpnjJwDrmulkJE3fdYlBmzbJCRHSOEdoHPw3PflK6DSLC1fmson53xOHoy
PbhfaEClYdEH4oV4116SsUoc6rnL2VRpp2ByMn8rah4xlSF30YoUcXuDyxDS/RGhG1mM38JQ+b6P
u0No0TTD3pEVaI5807VPowTy9jDqy4m7j/i5PMfX0ZCvLhzDqX6Z/68lTpjPxc6b42BeLa9+Iah4
jkDhxRtFhJIre5Rna+1a7bhsmkHojfrHNxR/mlWa9h63UJoOPmwEStJ3wWMxU7zqpJjLmwpyxBiK
5q5+h3MLpZSw2YmdnmXuuIZ2Ru/oRBVxfa0YVyS7RUrmArFQEyzRBz5jbwa7wG/uzFWVi5X8Mlj6
eL5IH9qjMbEw7rhaB4i5nmB0zPXMmxqgXSNpHIyVfmoBa6OrwntkVmT8exHeFnE81xcdmZuVLPF4
mONv5N5QlUOaNg+dAif9o7Iieu26I3/ReVFPiNhPaqfUvuhXieNmpDjv44CXkUCRuFUekjZKFMFA
kSLK2x83p97U7ffrqSusXpbfDVwzrN0vf9fDDw1O9Pu8pxyWebLNtTwav9+RKCf7WvzJL7GdYFxh
O5Qs9WS8td5QphzCbqDRBS9DVpS0KPCQPn4YEGOvo0brs3xP+liufkAaMmsaREYHgEDS0NM4cR7O
X2nvY0LidxVkRCFlK0KA5GxzdlAeXHhi/T9IySu/HBpy87Z0IaYLem/U/kUCr4fYpmOxfbbnUFup
kV8PAL5ENV21izCgCr/PKyJJ/c9eZvRGkILP9Xqhh/yg4QO7z0HSE72wgMX2OtxGf62/zjiU9HbG
Ot+M8158EJy5UtczuAZatld3aOGjBR0OR3hj0G7fB9p2LaKDTIIqUQhwj5oPZ8IRqIQ5JZA8YBAM
GdRjeaQj+FFPLHFPqu5FPsbtBCKhUYE+HsJx3UW7QFqVOm93zhp4HES9DWa8hQeH6dS7863icHdN
t5z4WAjbdhtXZzZSBT8y9Kc1FgxNPPCdY3zOWuHIyAkd2JWIGPLHHUFn2Bu2om8f6xLKDKlaGqnG
faC1VptTac3WgM7f5iaPHP8ybkZPMfFWvYeUcOaZN8zlRCpzdGQV/+z4yErjGqyp+PWXso6wrLO/
KDYfeXcyVnlB9Q303lezsv2XemZLax6lErogrIS7Vd3l0TXsuAgd3zt2qzPbcdlW80ipYeQQ+VPF
WqUT1PyrN7aLAGokoB6X00nI+tPA98P0AoBbpZV25DUFCltArSyY0Pnha3vgROGqlm4mBXA5Xtvy
vghHVLUM15+pBblVDieHsQnjbSOOchwEitaFBWZ/DC7jBKI5uNO1gjO30chde11euEZRXRGOocGn
hIDtPSjw1RzGqH7DHYACZIHyTiiQQkuJNahKk4PtLK+UUFVhICMFS4oT+A4wWVti351JSos1hxdD
iJ+pRtcEJvdAHFOki5+LljTT8qZeXfAkO4FDHKbTgp10Sp6kEf3o176ydso5mCmqWjHRk6iqMRi/
2uJwBgJuQHqlvI9ao4rIgdwSi0Gdcmq66j0yEPTZe7vuwQlP0JWOsynfu7MniRr0QXoD1O4dIFTn
VzivoTQppn3pBJfTJ50So5D/PWq3dixN5SZZkWHMGjz3/kkpWdC4VJ53gaO4fq5wfF+rJc9X+28G
Vnqvmk9p/1XsbVRO+kTKDz7mHcJ7mi3jjZj53nKoLO3SCm2qgYbo073Zm0R8CzVjNMWYkwkd0HZm
1vMlDUlS3PA/UkmZU1KrxsKpzDFo9sWcRoqs8D8nEK90Mqe9ON7k7kpRGjUtUgrPa7N1AzCqhApl
H/FcSDPvkX1HAxKsQ9wvhzJzdMU0b+4fPFrvkAP20oJ3rJM6eE53Fc5292u0Kizm7VeHTjxrYCAG
22gsD5dBhhTkDnjTeaG+0PRT5ugehW5CbRXHgZmYEjCR+zroRQCK349z5DbM0s4Y3iRQzcQU27kb
hGMufoyRSVXb4b/qvpDJsr3Z1CCKYhQ98M/pM8wcS8Gn+aPHEgqcMNeOuY080g7CQP1UWwmtp6Ew
Eo81zkv8EdDZfuwZ/YSt3AB4IdGish0zILOLUa4bg4+eRQQlQRzjIQjVMmG99ZXZY/QgVzp7KFYI
PwWCKLIaqUfdFkSPkWIck2DPu8nelF6lKjc4qAIOz4IxQSpxpFQU4kzn8LtNzNo5K++lUdh/rKaY
ZT7pBMBLMspUWx+/8ouW/65AmvhuIQkgWq+zlKB8mheWVA4s06KB6OBPCXEvyjhZZ0STolZJ+pVX
7gJvYbzocMWVA7pHEbfyulX5iR+JUXBicl/iIe5/WNd1utA3DQCkrF2K2pR2p3g8sR1HlYPWFzZw
+B4xSSg01qGhOruGIKFE6HUTB8UgPWDj965rh6pyoVcfxoojfg3XLAc4XsTfA8LawR15fK+ti4JC
Bp9tV2ZupI6Zx0YJeDKy5DvMa8qQ0m+8btEzCmc05slLJ6lwqSTOTrETaNgsqOYGwnfZEUFNY2JP
XSl2P9w4UehyZBrouhPRbTUOXYhl8EVpl/lZqV6mBVKjXYjxBS8g0uJtA/oetCRoBWsAapXKmW+h
Q7RChZsD26us/LWS1PzUhLbCnhbseLRlslkFuNTksePP5Nvp7syP7HLIg51YetUcoLIikGN3GFIk
o7dKK5JS0SORVy+OTdj8UTXNQCT03FhLWxw7ccJBb1GhOxM3aBuw1SCM5n/NT13xGHIPQaHf/QyV
A+gNFPD2QvmXyXPWMb2w9iUEAzUi4HX9Nf7IgrMvxqwGcIBXoZSzjCPcTFLAGVbnB+8vNmldBpvw
9SLlNeQkmmig50QsLz5IVPM1t/+/XTB4rf1B2fHGXjGn1hTQ8cBVPzFbqfZPUM3D+J7hetb5vOTq
BOcCc8Y3cxDbSUMsMal+26RsHDEj3zgEEQdSdM6i7fA2CmVRyjx6lbeSEkWU2yVjfvpaZk2DPP7n
/05HoIZAj2NdD0H6lEqdhIZ39iQ3Vy69f7N+n/ZdVbcdcJ7pZkDPgrEwR1Phjy/d1hbjrDS2BBkp
/7783hZ3MDIqzpBXKIyduDnr+UxConW3fhpJCo8kPXBEYATLo/lH/CVqS7Xdbf1Wkf70wPIxQ18U
bEPP4A2+RBeX9pdxDN52uQGMUkzi3XRM3DryqhaHGTHP6qJNyUy/GTuv38ss8gCj/a26/1CHNrIO
rN7KdtmYQwzFZ5suyxEVb4LMIMX6y6E/F2vFdSt9WV7qJl1s6T2nVlAVma1JKriQ8Qw/mpbr3fGE
dHgr6yNeHOJUcx2q4IxJnrc5lpzokVts+wp60pmgFQma7VL4IToncTQOmneEC7jnzysl3L7jFFjB
tDSz/h77KvZu/7ZFqeyW2/nj193rPT6upNfCf98UUcHZlq0CbOYbqJgPg5xpal7WpRvgrO88r//X
O8xuHDl9joHh9uEHr7I73L6Lod5z/v4agS3hDuxy30h6f/eCQ4UjlZSaw6LDsZ7pNaIfrMfI8xmR
6cO8ni88xBAN+xvZyfAPIY41sS/3Y76DUH4xwezcrbWLs1WypQptZy7NziSSl09KJrmbAtbsCyqD
cJx/B6mkNF03FuNh1aDOU8tKRcm5KqE6Gn32uydq2qg7BeuW+xY3UajcvF5pT4RetnyS/iroK7oS
j96pZPQrkq/F8OW8AZ6FJusUDSwkgvFzeu9jSNoZskvE4okDwlg6M6VjI0QBcskVPdJluV36M+UU
Rhxlwy9ZKCaT/rvVlJPEq/lrL88w7jpx/XehU2YNmveQVLP67Dx0OK3Dsq6vlIBL09SISh2CBrnm
Pba8JrbMT/q2t2LutRFI/OKdLzgtOFeAX6dU6BWjfI9gPLfPTeWjIKDcLruGiFXdYIuByFjQN21c
es5sA+P/VzIq8e5jb5TqdCmmbwaFogDfjuX+fWFjmJZdObmQGuuaT9souceqHPNdlBpKMFgj6xeP
mwMzTHYG/p9dNYk31B9oWgEI5YbHPPJBEVYLXiTsNl6Fl2plwfiu97DOjXIXqSt9JSQEauALAzVh
V8GQVkKcapghDcUED97g2J9t60K77EjNO9KqkThHGpXpCWjNAm7ooN/7c03U9Epu4AvNGeyWay+y
QOLtObP24f+eZVwGkEriAk4AYq0xkiSHF7W5P+ikbsXS8dDwdky6Eb56uIQcRu9aPy11m/p8FKj+
tyrv9ZU2D03p4+JZJwyaPzFvgsCci8X8pMRErbruOzBS15jm/J1IcWCLgReG8Vrk2dCem5J6yqdc
NFXMDAuY6eEvOM81Yf6z4xMtIAPQRG5o+MHnrhFuJhJEOClcg2Tu6+QSYkRAsb7qfYnWmixgtWzo
eNSXCl6meuPSyUiKetTKe2px4BFX8RYdUN+lacvv3ie73+tG0tfliI4Ml74XHAPpycQwo5rFPoST
kOwBAK8Fpdwp/B8Qoo+MJ+Q67bkiygPlwyqSRc0II+9r7e7VGgHG9XUC5r5ktdEU6UDJEeQxm6ex
41cFKdrt3O0UH0YG6g+ZASVQNzWv9lDqRm5LcwnQNESTN15zDiSIFGIVmlDpPdFC8C2eyeMRfKtd
bnWqFce4FkS9vpICly4E/sq8IQ1fwl+7V/YZTjVbGFZYqLsnsKXJnK8phRaRaEd3Ao+7V9WkPeWS
EiflW7OImCyB/Z91OdoO12/dqlM59/ksCblnZzvZ7lFCtuOF3Ai4o1QlfuATB+Fx/fm2x3m8xkbf
O+twdl68TFOU+Wb0lfEyCoJ4lqhRIEl94vEtU9q2dJO2fRDPokgcBFM9jYn1z9MVCzUbwo7FmziT
QmFZn2gtz8zXg57/VHnQZtO49n2W+BOW3umQZaR8CkvoMatV4wPOhGaGi124CNM4ELlN9KN7Zf/+
eIypIUmuQ5gi+RPuz2tUW+lHIctYiJr8JupC1ZC9c2h1Q29cKz+QF5WJ4lmoQZcpZ2JKdaeowQrJ
sAPTXtmumnNWrXm2yKDxPYNLMj6du9gVxnpBp70jzfHt97eyQHbF625lHJXJFj99PQ6csoQCIZFg
PQHOoYIME8wyjfYWKvi7tNEKdPmH48relapp78dM+TIvSTGKVbJWLlvWnvY73ZPrgT5mJ8orDcDg
2WZGyM9Cc8vRgvxibvymjM8o9BEZebibR0vxuVS9s2a/wQHMT/hPG7Y32af4gzS5vEUmS9Pr3Pdk
ren8Yui2AXKjHdwnnGeH2XJjKAvIwjTrpkcNtZy2L0xrxhoZrcC5M5hny8ubXz8EgC3KKqdPzgKC
JZxYlzpRdUXaIZq2lKwS/oQ8fhBUrd5Ycb4PYyTm+73RaIatE0eLl5WPC7HUJVdtrsnLMalgH0b1
Xb88SJvcTMqrzN1Ciu9K+YhM/pz1ldojAf5JJbXaZt/HWMoF1f2iXNRKrLZuQgb2ioQR6j7qjucL
l4jYh+xFkO7khLUewZGumXXrsw8OJU+XJE2LnDS0jfLVFtvM4xzk6ZN9NuEGw7OcfQTf1Bt5piaM
jvcGYMnWby/wMFHKyBa8fGnS35dI+E2J5/tPL16Rs+fEzG83TBpHRcAaavcgTO3qgMryT7c5PSFh
8BKzFZumvN7/CKCRYefUY+nlEqSm6ssfJNHZbW+d7A2G9bgwJZZSbP7UIaYByWuQW/892/i9Ng/e
NRfx4rEjdTRlcsGFObeG/MeoM1mCdRd3JD0nLd2b3ZhYUOO0yD7SZd3J4WdPw/2gPWw1PdSDVj2P
1Fje0TT4nP7gvcbDufjYUQbH4/qGJYDn9acjEutXX2M4cuitPDeXSUpO+bjfE5XQdu+Uy0voNZCu
4f/T3EaBx73jhH5HOxhQwU8pSiC5hCxkie7RGODivTIjAU1CRzH/fmrU/6Ezb+ESrT/W7fbN1MP9
SzVwRBNn7dx2CQ/Q+hscsg/VjZFhG8zqK9I5LTeuUbextQ3X8yE0EQlFPk6SSt9nQiQk9EDznYdh
jAUe09JWTr40f4smB8zdZYSKpsKF8mpZbSjJUyR3WIiiex3JbkQUUBS7c+OTiQfF+rx+O5HsGqSr
hhjFRmha4Hi3jU3dneFcOY7Oo336WcSugrbVKbRJrqTgzNTUQDm5WWxNq1MCXcteQqoNF4iYROIm
P9WdHrH3qDuPVriRtxjrOC2yys04Yr/gLOi7pLJ3+0cCNvKxYnzTVogaiRUV1p93HuH2KVHRh9fq
3VWWXK+5tFPqtPf+3UlmvAc1q8+T/6hzwMcRsW5VE+V95VA5L7RzTFh4z/pf7DHUzAEEskb/CTH0
YZ0hyiYwKcKAzRciRer0BnsYX9oWnC1SGf4ExHRJW+67I18+aeGzrHWL0p72gej97YW3uHL1+hbR
BrsHneprB1uy0rLAbmbQMposynE0vg3DkxbTpE1ZRd2Ed7kZtBfjQ0ymXzXw7P6s/cd/XEGz7Ejt
tGI4TZQfy/CW7uQTi6g35xknVli/75ffZItmrlKP4Nsy+T90nS3XmYieDoHEx9vF6ieVxuoO7h4g
ZO/ZqIVkj9p/O8f+PfKVM+VB1QLHxC4gW+XMfM5i3O9Kb5Wf05Dh+s2POFt5tNeUI5/kOKGf76XP
RuPwniMPrZ7OmKTkOTuBoyDKMHYBpJo3veL1NYxuWngcBBVXx0S2f8hO3UzpGK3CY6A0yetLZ89y
he3qj4XAOfgpxRl7ffC/ejjsWaBDQMESRbdQfynrh6WY4jaTwmwwrAd78oayYonKUDPhtg+a/zjE
UcReD8V64/ofxDe0uJUkRAhAfsqo2BjFLSo/64nI3PCmUPOKw2pB2C/y/IujvGrniqEtw1uaKjPA
K8nZCaBTcaCBJe4v5nXTAd/C2psRRSpsa8BXzqOjx9rjn8A/lC4B9A1F7GjiW7nnu8xDP8hBQQha
WTjrAuiCesRslW/4EEOPH1l4xzSap5BwIzX1W4jDM0D/bOdZUYDevuc82cP9WiZkrIeukXCDfkog
Wvt0AOl3f7V063hwgm61slL0CPZ6jgUGOUEcdztIkYjVV3m7rXp2+/mSWCYI+DDbTgc76E6XlVvk
RS8zNY2PhQLmn8MnVtZaMpZuuXEahhq/s5DRAIozSsRzttau/HxMKlenam0rKNvk6sqZ2yR/K939
3BHx09f2R5FJ9StwFtmTCLz4nnAyf5YN/PqWNd8Dn/HhNVnsSDjCma6HgovSxTd3f/ug6HKxvFV2
JbKbuk6rGc0RSDCNztmRocFP+3GSX6bNEmMbQCs8e0Q9JJDUdPKO7FA3nNnEexCV2L/WWbyif/N6
atEqqiepnH7ipDvu0+4Zns+1Elo/AQJ9yXT6dHH8GKDCup//pkf4TEs6COfghfJTXZxcNod/9YBf
+GdTcqF65LxiJbBlN4sVmQtEtXupZI9IAqFFjP+tD7/S4lTWdiJNi6Qv8GNcAV3clkjKiMmSvKBU
Iq3Q91ZemTZNV8w0dCVtW0DyAiKGMvpuE5xXZNYoHlbPSClH7RK+4kmCNn9wORvbH3Rsg9f/5KGK
3foySxuJvfCLAjfIGHFnx3TLM0jIGFhy5rgWJw4dq/z2v4zGeiZq3DRNN8dzDaoctnZ2QHWbFb0r
XNHAqHLZWzkLouSA9kx82yH+aHFjj108gBuNHBeXnfWjpF+9nvYlhJ9hZl/LuA+STRL4teDSBUKm
Bnd+mo30sseBA9d0lgrqRi+5zw+UbIBS8ob3zHFURam0o10tVABM9T2ezvviLpAQLSbsbC4vmHvl
mJPa1FVMHybrrXAsgF9nMhoe5V05ePUi44KBj6cEQ8hJN49YzJwZa3Zp1349eqp+r8q3xMq7QR3A
gCbMXPCWJuKfo/Sgj9erCnIGclu4fGWqYUFmEDG8B2TWn0uYakK1hm/WYj1lAxEvGjGpo068m9z+
beZd1jprcyGSGToUvE3SQaRCdp7TSAYqmnLsz7grq3vaEiqLuNXIS+JrHoPnzTPkuvJtLdO3CxO4
dZ/AuQknnFW6bMTPkkvgQPYRKimQsB7YFgIOOUn2Wz+MvTdPqit4bMwWkqpKm/7IT0AJv/VVwSmR
tv88miXTRCJbukyEan4iW46+5i5w0ivxH79J0syW/uia2t5O/wkPGrA7PYl1V/dE8HMHrmhmvam7
7KBSDZgoXi/4VqkHHZgphmBLiAOY9YgCRRz994sx05eZDULw/LSIh9ApoFJrffBw/J8Kyg1hAf2f
HlzLuc03BzsNIBjoHFP7V5uvYsVYdVeNwqRPfJYNCJa/Ore46NgPepTWYeqzIUJxhsQv9N+XxFEa
6aVXiHYgtfL9k1xZS7/A408DBgHQ6+TTUIhQDqXlBjrAg3BvkqlerXzn++Fm0/kl3bvG873liVve
mCxmbucOW+MNPiEYH4k7GJ24uiGigPtjnyU9TEDIjzJ9LAsZbv39ctvMODbmumjfJxEbQv07Hk0E
BeIAsvP1qNIKJG7s8joWeo4HTHbYm+mQfenaLWPZCszImeaL3gQwOghYwEmNIqVXLr/wTwUQPu9p
ITK9w/TBPmF4KEsAltfL4qGqyhIgFJVkgunzGzV3rgckEugMZUi77R3qqV/mnDcy6s+H8gUFbxjT
dWs32yVPcJnhEJE9I5zkXWM6MvT5VxPZvbRY1syJKGtmFnszyMNOAjg0mfIRfXqttXTcBBq03KAH
xOwRwznJ1mlLM2whxz3UjsxF2WGzqbYINaokQFbLszAyEp8TvPN0VdU1FKtZRfYOR6OoZX8noIqA
108xTkOi1W+YivW0Nba8o+d/ZmmNTsgdupTsaA8511NZUu5GXVovUQAHhbrNKMMfXgl29OaXPup4
7hT/ff1fYmNsYdBHniyPQl8sg4JcZn6ftxcIKhes9ElAeYfpqUC5gPitJy0nvEOg+w+QoJ3W/EA1
aqPTXEqLGoPp1q9hYG7/BOJt/KqQvJyeREykxK/ZkjwYi85Uj34povo0NMu02QChNBRAKVB+tvCQ
NcZ5kQdeOHcCTtmPK8WUCWhdJuWaTAkRHdJjMct6j0jhOiSvXKlHx4hM3+PNFDKmrjolEcYAi07P
19SyvCjx0d0/RefMQ+k2HESF5Rsy+rHWTFvOghJugdHEz5XQLW36/5EJtO74ssYUgiHIGp04yf1l
2b/DZnN6ZDkTOz38tDR1JMa6PrK+fOQhLSk3DqtM9vLTb3eWu2uWJ8QvgxfllNOCq2MebOPf57zr
974Iuxj/UBTEun7iinTDAn/q6InYkCGHEhh2xOa94UuQAMVS/1kN3z88zbjTQueaQ2J+FZ5FTbAQ
O+vKlwDqAz5g6p2PuQwWvJ+RAs7C6KHxYDMb9JpVTqh5niRaZ8C5+ptvu8OXjJL7Go6VMXvDISEc
LGcBc05xpaP05FWL7TtChG+rzjLsTLNxwDcCrI5s3QoCnqIE9224eI74SYG4kUyEHzcXOXNeC1nL
OIHZHY3MZIrmpRVAiK7KUsPg/5Q85nGS/fg2sNvOtWv4Rhqv6nDRyNnZQOu4LoL4aYQKviv12no8
PMFtLKdOUjeJQs8Ur0fzZUGqLiYINKhtK68+ZzpPCrahEkVqMN4CyBWoZDFEmj6ABIZdBFIkTq+x
0Se3hrb13FrOYXKM4H3ahKqY4YscUtLHaKzXpDkbpDrYU7TEvHRAGsmGblg2Q12HO1axCdei1juF
OXB2v+6GNmdARSNfJC6cKCdAsegzhWdKguL1G65DSsDV6IWgrf2hlGEjGhfyWoKZZpZeWizLS6dx
ZeJw97VcWBO9U7fWfLxLcFcqWPs/T+7mW8DvvvPD6w2TgAt7BSxQHg/Mjtpk9UD9jZ5SezN275xI
0aMQh5J4h+/SYKi+zb0SVI89M/WbqDzBTl7txMobW94fMNmCZVDyVaQBQUbrKLILfH0vU++jKl/4
VVi2TgB05zBFbn3+UgXtR1aODJtP8UPf2LP0udugmDZlPqEYjSwtgjcNOTUml9+tVXcKnFmsJJFO
GUpCJRRO4oEZqyd99fPSCW6EZzJAvIPwpPYevvOB97jd0/i/DY+6MpNQPCEQ1PQt46g6FMIFr0WE
L2LzYUdqtagAXpBrD78zuKo5vRgSNORn+p653180k0I3JEMRjI+E9FIUZTtlYFjkdPaLprOUiVxH
mymV5NLcDV8HOKeWX/YHas+crH5UPhYiIEexj23CaImlozUZNagHVSSrEbOzYPgAH7Wru09KleVu
+ajW3CvGBIANmqOzurjzZlj19xsIbJDhzXHdSf2cMyEEiTmxakUnnZ46mIhvEiP4+gsk7HjZH6g9
4m0N8OjvM1UPG/65TqE6Nhrsc+j5a1x1jCweA+dNdxznd21lbUWK9Gas0OKI/UTiuVdAPTGkQq/Z
bDnmrKcxPcmjM8mWjV4Cb923e98adwQ8qsjC/rn874/C68On10DDLt2Qh4n9JVi/iZ0jvipc7/Pk
ywnHKIPO5GSll3Bjnsk4t3ci18U7ArEjjF6XMqzdVGPy/NcGdTcazYFtZLJ+AY2G4rw1Kg4/3rp9
iyFW1eUbTNvry2Gds5hRF2uWaa/JDw0v0cUCf+oY52ebDpltTeZgYhR/0dGlcjsLRekmEiprClI3
5Plz3thPExE1FFz0KfX1+uXItVaFFEgVODZzpDgjjYfyHVggUTp+oMWKwcLoDxkPWmNOt5Bpnpxd
9EUHUC19MBQDHWMYtXqU1IEXELc/UmspeLNECVZeTy0D9nygl6RZvEpoKy2tVJjfVAj91csMF2Uw
cbJAWQZBmLWVPBrF0U9gk1ly0vUnarBfrCUoxt3yM3Z+8QJIlyVrb/sXQKjDI+FN2tsGkp84lwby
SRPcWD9RlXpPEAZRd+i0hxk+eaC5ZvgQEjI3xDOdkJOqIqYtiuB4xm+rTjlBhQOoQU/hlW4n5AQp
WXs/cYq9iIQpq1a7bW17ASfVdRjVfHh/6yy0JSEiQQ3lzBWKJyzif/IF/p/ARaExuadDbfYa9JyK
lMFITLAxs5dw6H3Ru2/YpIkTMSmkTizamp8b9b7dQ6Fwu7AAQ/QRs8g0O2G/Xh1yxIvoK99HPf+P
pEb4j1MwMDlARvRo6MDCy17J0cT7ckHyKBcSgtO4102oWcHVFYnAd/odaCCUvaeEWtOCLRJGaYjo
DQOb8S0IwF8fFejMdt6YEXaBBwnAgPkFXlJ+jnbgYfVoFJJvBZWJ9eb1Zz4KfnIl98MkqBx9JGzB
5HmmpOKnx+p/YYQASzNmjZpP5b0K5pREnlPOTKKx0AAqdPuNBanfHTgfUEapt/3ItGF3EdW29Gtx
uXtumr+WsBOFJzs1CX2z+RS/NKdfeYf9f9oqC1YpgNK1cCRuEt7ReDxsDAozBujpBKZ7GjLBhrlO
HkKR+hQ5bC+CSFOAVbUpcmBjZKPrDxtFjAsf3RFRJ50C7mo43yEdMy+YvmbhmmKnkzCg2z4NK5bx
4Z3VP07S4h3+q1DaqSV6Il6zocB+U3CXiak9iGW8uuNT8YIvMdQF5RxuMENrMzIiZBLQ64j/57CD
Er3ekONKSyVZSFbJJpBPGj04SrsNIXt0xjIU/MKhXPElMZbDFLUv3m8qjmsT4rxo9cTXRfiKd4r4
1AUdZdcIpvOoUaxz7NE1plcLHH8YEyYLtItnO47lZsxF060ONz62X1yCom+mhlXOihFzCVm1uMR2
jrPWnKDnq9w8hxnBNf4P6XuVb907hmSteDS2w+LjSF7bk+3V82xpw0PX6TibLRwE8YdtCGn33inb
TFHDTWrFvqWDt8CdpUf0UGAIksMzefQCLpCilEslIEyWsUgk4XdA9WDY3LiJyuXUa45kpkyWv1Ih
c8BwoWJrFUxgzo72A2dpGKjO8xV2tqiUEbAbD80NbQ86CpGBn1ZPTDBDUxqFaVD51LrsckADmyBN
D/sUiNWC1qjT4h3owwgjJz40V7hT3LYsyIUGXEzAu90I2PZl1F9wyWVU1J4O7GiIcYsyLtsxA+WK
2FyP3sI8XnM3FkEpeom7d9CwmmKxaSDjIvtF6cY9a9HveljC2aqp3vJ8IxowMbIcWI3LRMDp3Qdk
jRJXCxW4XvKeaDEHwSMtS1eEYZewOWRZyXTfBQI8hv12t33D+38pKEW60pOGcmz2lzCoJnt8gPtp
o0lTa/MZAuL646cD1P0/BcSNQBjx2KuFTSGKZxE//ZjSRmrZJllEqH5RsnD5KveaCuWubORkuamP
t/oUrAzvNHDzBBVbgcPqZbTGgDs/b7TPk6d3gx0k2O9a22T1u/OJDsw2NVsjik/vRrf9mnbwyDQN
asMabDRmBKwMgAb4E0siRZGZ4j7FxDEiN0ND+0vMLxwqX2E2IimZR9dCf5zEtUdBaph8vRUA+q4f
nxAnl6sGPGdxUyzDcx9tCXhSrihHDD1ZmuYmESaO7l9Vd7IsYzs9K5j0QhbZxJLjT8u7lXVKwDX5
0WNPn5r2pTl5+hsgw37OxboOlnvsFg//ek68E4kYXpiuDg1tOVyuHs+Gpm7LG1FYknY2cPbUzL+U
Y6fktYiDrHv0KecHMi3LahChZjOMpE9OnnycfFNquLWGAH8e82wBscykpxIsBALeVIzG696Uhlta
0DPxL14pVgEViGbGOWKI00GuNJrcsFnWB8eJUVV2op+OQg1gL40a0IIWfDPcYFgfcdCjuVBAm+x8
b6t10ruE3EsOP168GwhU1FWpQ4qZjZxYNRproW0PY6+kSs2CHz27pHBAWVtOC8OtcRp/DhH0KYI6
fw66mbf1WRiPwUFm1WAKFknbI1ki4abxSV93c4A0TipWn3wu32x4YLuBCV8SFwW/Uv1yH42mpqrV
oIcJgI3M74w1NRHFY/5M6LSTqV3g9kaL2CT/PU5IHV5Gabzj8z+6fUvV3eFXDWvVXeUteVgDNYUD
Y2aYfx2V90SC1zHvX9WmFaJInousoSY79Snh3UZFGhd3dOCFm9WOZR9LtSEIv7vbMTsC/QcRfanv
cYszjGBsgVlmr/MC75eZ8AjWr0XQ3Dy5MEx+V/yWBdhA7wfosLmo6tXNs1OtnrN5JDAsqpotm/ET
hPhxSlUm/f5lGfDXUcXKjC1aQ3Op/+ntgDYyB33OR/tRn3LMGrWzycObgXDIH4YL6F2163D+2IC/
/uV7bjeeLVJR5W6ApM0BYuKpEhxAG7+oGrcH5jrSFlGX//27uaXbaHBvznKt6JsUbEsODu3imZX5
qgZP8EBdWyrJPVGDcAf0ucuPmEuKfDXbHelMMMfTY+TNcRoDxB8N+3Htd0j8ekKhHLCZuvc1FAJz
8M2sl8qFxtSXXv+uQSwqxfFEsSYEsZ7d++cjyp8n9RD7uL/3HSWOQumMCEqXPwCYXjq38ceScUp2
eA6A0z9iT52ZO234PWrPgrtaRkRj1eYVE29z4uXr7QsWflVNQKClDyAKn8KY5gh8Mut/Tm78NLmy
naAjqtY0fCPXb4Hg3XZ7LLJ7tP4kv66nOYbkTfjlY4OEDb00003nbubP7h3n703IlcGOJlvzN3Pq
fZvo6U6DMr4+J5W3WgmhkYtMFy+pg0Bou8e17BTdNajBoevVFMB9Qt2qqtSj12JhbCuvUAMf4tqX
LG1pk68StzgZdlpM7K0/XKC5+XOtCtV7xzP7VrfbZ1TokDwmvqLwlxAE/ywEcJu2y2qz+4/4iU50
j8aj7hJrU+KyAKwKHgV8qL0ZW2iTQGlNL6skKwEY94uMhqnmSIcsCG4Pwt8bKGprLE/TD1z8jlwD
+ySgQmjRh+W8SF0nfC+T2Rk0sDwmgLgTgq2TqTSJCTxpcuQVJRQXYtwmnzAhLFgVydByTRXwzSaB
bmuKs1z898ocBS+qfrSUWWZW3n1XnRSblUPBxqvII47POYS9wthc7A1l8lZPHSKNC15nofcsHFhW
+Exw1UPeFSfAoK63/KEy8LG0bO7AptS9pIdYtOUffFUfl8vdomVABL0ZqoE6Ob5/22Zzi8sU4cLj
Ew3Sc79l0tS4/M8/DsHBMNsP4irtzuAMsH3zcJXJMYNA5ZZLiSjSVd9zpIC5nFq24OfWa47ZKD5u
4JncHyfwJj4F+z2ENy1bvEnCJEJD+U//vHovmVm8piGSDRprbO0qiBmn72kREL95Aa5xbVWdAroh
J0B5wmVbRzJK+NZOMx4WduxVzr0qrootZWGEre1jit6qIFt+9gdYrz3kWcLMLrCHuU6XAqp63ijC
q6OxzBMdamQnSPx7SMaNsyOdJ3SNuJtGWxmRNK/+fVTRDJIw335k5OLgl9pyqkbWkwhXPLQ0kKSi
iA+4mk8Rb3ZUHHiM3EGEBCs4doWkCkJIPG++U4eil471GVJHMOkb2dQWvhuFuvq6XfZKuYXR6HW2
KWA8fBSwwpvaOvbgC8l23X7D4iD6D2OcBNjBq6TGk9NaClW9GEjZloiGwZsZ/H1ZxUG8Zjndb7Ng
JhQ82JEslk3LyF5gBZ0EH1rwdgzoKS+8yB9aIGCmO6/Po+ra5/d92aLjsQJdwSQdrG0XATEAhMoS
hIUmKz5kmjQX9QmPREEflJbFe03Du+oUSWbKXg1JRHReAhw2kDw+c/FEDB/S8G7qUWNoY9QKzx01
bfrnTO0Da1+dWg7D/fWchdyrpL0P0deLMqFo/ZZ3e4i48INcnRq43r6GRTgdErqzTl59o0x6b9Rm
DaAUB/W57qiwjnOOQazgwZemi5Bu5bxDFwDvQXpoqcnnpwVvdbc1Amy4lea0oNd4vTO7DoSBFZ87
qbJWv9/CcCFIbNcPqlUDROGr5kMA2aCzwqZu0PpONYJ8puk/MEroSUTC9bJuvs5/wxrm0JkaSkzq
Z65YsFB0HAtBHavOubC6Ui2rtP6NceeqnJH60JCKNbP0S+WbmjKnHcYMCgbs7dt4CzChNMd09qns
oFo0I8WaSeNdRjHih9yt9mUmMu0twjCehEC3k0RuCOehH1yphc5VmiAhdQxS+0GP67xdnId/YdOc
RduYlGEM099K0t2Nqt0rPolv3ByS2xEqlhSZOrThTvcC+Ct07v81ADkI5UCGAwQfwrYgji2aMH0n
ZDW4rmoh+TM4YnZ72RvELAEVqzUWZFC0QjNKScfbA/7Gx7uhxQaGHlVeYUPu2h0bFu9JyUu9i8Ax
2OpQY6RS649gG9XuM6l6Da4g0IP3XceHWZDp7zISb96TAtKjKi3pRrgr+ZLbOn47b6jRKqPkmshi
Di5RDHD0RVsONJlGf5EWv5F+7Sgk2NDNj2UJuGwPYouJHOKUoM8f5NfbkDPle68kdZ/oma2WMjkH
mGQYTbMm+hbwT3RgmKtp1Ge/TfgiqRldyYvShKg0DWkWmsv+yM48S826HQpmHEoWimO6/V20nLjj
oBPIdLt5PstJAiBqp615DLSpVgcD/V1qv1NINn8niKyQ8KJLZpnGw6bsNzzwWF86uhxNDBnRANKr
b9bOV7v+zBBV9Kvjp1JLQEdxEToxya3cPbwpV91MzhwRE+aYRI8gRvpqR53MQQHL5SasutLX/R4X
jtG3zKTcco0GBYoqfM+rkSkL5ANHgymSOzKszbBRnMkyLuzQAfgpnZujeA9DcT1zkv/XtN1VqB5r
rFMl7I3WeiUBoKsPuoTjbzUdeEKHMzcVsY37F+jrzAKr+e39EcbsJpIejH9FtIZXSueeiPHYEOcn
dSywFfblgdR7gJ6cAAckXsvdFW0BrmiSHiuWkyE1h0TfAsds2+40v6Wpea47QJBrH9Z8i3iJG5MO
hqb/+347bxpiqn4RrQZumqB04P8H0IgKlQxKEP3W0jQkPyELCfuLCoaLgbUldoh04qD9zinq3Pvm
sWHnHWhV8jX53JhNyD/hfr952YWnNxLEjHqCgG8txyn9BAMK9ydsm+3TVaAYG6czxe3KsSrtiJNi
+SXUzfVmjYT1Cj/8G8bBKNN8dpgD+Tj8v1lvQfCi/qhz0lxFHUPlAKt7G3VQFcYJx0WMLJRnuduJ
ZClLJI1V83udMVV5ef5d0RKBzJRtjZZrOYhAjw/iqnvSTr9iPS2YKDcLV1t1bmP5HNwh/S+T1W2C
ybQ/QKh8Nkifr4KyEc3SVeDTAvsxNOxS3oUq9QzI3XPFZ0ABM/uFX7hm114ocEWlIpugE2LSW5fc
vtcwH0cJvNmVyQzGtxrox2nqxGLIJnbx4VpNNCFyyh9O7f2rtGFcpz6lUE0yX6uLG4LW3BOStAo6
W9D1Do1GFw5g1BBrbwkiz9M1msRMmmVv6UZO6BPMTiaKwiywYZGZSvIXkzVHHqvoppT+3WAYYjmu
+FNzz7gLse1E8TQ5d+1CBXglbKxfOxa5PobEtyt75wYnhy+RoV4sY2+LS4DKIPZS3/pJn1dRdPVP
0tY9m9V8MCTgk/WNmsADXp1PDnxoqDVZPLwfLmt3OtRYLtSzkea3yy8mPy+s1ukka351XokPgQgU
tpLQ02sewjrIHn3GFSiO0wJ6V+755OcCkQN2jHqfxbzFH9dQdcQ2ufslgz9EXD/o92kSxlLaSmup
P81LbiCtGXFxrwMYhrlvx8Nxv6y9gUNV5u+Lo/U6mrQTd77LYXNLZFi4MRFFaizJV6KQyVNcPi7g
RhgrpItbo+yOpKmmRmWZ7fuLJeLxHl92lC0KX1/BugVzaG0qcKMZXKaOcwEXev7bkH86zFfyJ9Ub
UcQcuhkkXvifX+WFoQQJqViq9rC8LIHboL/Lb2U0TE6JQgUaTO0YlNq+Pa/N4Wy/SJHaogdhWm4p
ueORxv+JPH0kzBrwJ8JYEKmogFnWluNj9OqJ2tpWYIVRByWnHvdLNPmjmKhTiOUEbOwBlzblv4g5
Lybi5naitLfzlhBbO0inhLySwHy+vvB85JEZbnAyJnOb52cENyKoZZVEYixqgkkXEc8cfvdPPSga
BoiMide7pBHHQDhpkGEm9Acbh3bgVV/9ro7kHQjVWxyRKCR3tDwp9ok0VV4mCeSKLurjJZS31zHR
3Ie/guIbT08/SoCDx7cKL1kgbWyGGlM7j+FHhAlb7I9FkNNREA4SIsS4mUt8QrgPQGR6LeldVhGX
hvFEb+XNQMWjGBbmIWQhZyD96dFQkvXWgBAv71O6Azm7/cmKetp+g6JGdp8jzqK/tDQsTDUmTaAT
HBysphxO5uuLtODl0+LCYEll+boNFCNi7lu6s+sqyl5eTsQjxNHqCzjIR8r94x+Q/SS0Hy4Viunt
7vG4SrW+MIt8I3KaZXAU9QUEQEGlyNVlcY6hKzSH3pkrV11o7Sa6QmqUAbJ+cojQbnqPkf9xdgEQ
y2oSeVzeEBJlp0YnUumkf/uiVf7TTgrE6bVHLckLG3ITJpgk8e4PQENw/8kKJ0BXGs1y+88dWMOW
7YHX6tiEQ7JXYYCsskByxWTR4pxGqQd5VMs9JmcN41s9NlDo7QgchfCTR9Hse/jnJJGPIiVbQG0j
O9kalRmn30OpeMEwcALvn4WdCU1AfnQ7VXG+LKatEWCZW4I5+ZErVQi2A0j2ore0So76P5CCR6iI
by3wlj03cEjYGa2i8jrjnCcgV1fqupAHpL/WLdisDLwhUpZ7pQ+pVM5WP68EPV9p/NbELfeJSw9W
Amr7cTaXDu8MTVrHYPwshG6XnzieICj3zquoaz4xeuhX1gT/wa9uzFFYxRi/EQ1NLROI0JLaH0s0
P6rWtoVxF0Z3IcBPCG6ZriVZIjyp1U/XlPu26475rG1LXGSPL7Rr2IYt+qjA0yBhfQbR15oVaP/l
e20b6anjDnn+L4m/A3rdCHj7KPirc2jJM6+J32AS1f+fhHtm25UL1tdTMDXLPodU0eWWkDtfGToH
HF7fW9tArijhM+04vcwUCSu/P+/gODMXi7FCuK5UjALyVFvCwRxiapgn1aCA8w+aYwTWSUGAvkjC
gc+zptnZjwSZ4hMSRqp4GfjBv/hTrKkal/91Bgx1kyr1su25b9HlGlpTSyIO8cNsNBJGngqII3JR
miKr6Al+VV9fQ3NK7IkfVigW5jeDSNNRUZq9sTxKrBii2TEebqnSYYnYUc+xzIjEE4kHaWgv82pR
UNa/N6xzzrG58VYiQviWTamWfshkLfK2EEJrK8+IbXGTde9BmaBVDD8P9EO0kX8k26ysEAxyWf0e
o8lvuLTaFAP9jfgLUpx1Ez4zTtYpy09j/0aNf0THsmHzGecZFDm/1X4hSNDKA0JKKfwdHrSwRLQm
4mU2rjxB54k/9l2bitJrBjQH+HCY+xyAdHSs9j0y58A7Ou21bXyTGF08I+VznezzyUgurtz7/q7s
wmNGSkTjSPjqiv05MeEybNu/qGe2qGnCnlVJfH3rvkUOsxNsG3wYvfLhaXMaIUzE/iV2aJt8nRqw
NlJ5OIyMoQzfCMVPUJUQx5Ruky9wj0kbZXnY7QTVyH/cuJDHCLQH0LpypYaKizLwQThX/s4XPMJm
tAt62dktyo2HDSDmsL/qx6nLgEO0ONGYulaBdplT3fs+GF7ZxZuEt16+xgFXRYjaPM0mkuA1aBSD
FaeToPW/87zfRKZV9xznLFBlTXUS9IgmHrQo0Qp/AJS6o25DIjgeL+jgiTUiomnxRtjk4MztqeUN
K4hZzS0yynIaundis583fdumdupnm2ynaOQfe9KRFbAEaW+/8BccNFKOXp5FWlns70KTC+bYZyC4
0eU40H0rtKtJ6phb//E9tjlBczyoizD+5eG5QOrE5ZYSYaYyowNdurpd/YZ4WgSp2yRb6s4u84SA
6z7+tWrWORltrWIyEcQHKWN11ObmNIKmF4ZLyWDeXH6xMUJrmvZzsv3HyRsXHuxXtEKLmbA3Xk4f
EUvI79Aw6h4KHKLBVK8sqScI4UbedeJ1xu6xT7T+wcVYXNV+IWKmni8RAwWyDfkOoKAgcLZVyqnA
zVZGYnfqS1XNW//VQujnRdjKLuJyFaB4yLTXTTt4/eUF8pz58TG0zBS/IG2xfOd8o9JQRkhM/C+R
iXLocv3amcHl5I5y2wbnCJJLmhWfZAGyPFiUz45ele3+2qSE0mFLQc/XFLdjc0+Fm4i5Vwopf+F3
31Q/TC/4f43YKbxup8r3E2iuxArhaLIz2upLwI0tWOhXV3JkZZyl7Qb4d1SAusvfHrC4Dps+/vDd
XLDWhTa7+3Nx44XjIA+enJxkoFRihE0sDAbjL9pLcp0wNyg8ghlMH1xBi9Kxo0RTFfN0S2aRv1+c
ZWAOfbUvm+jNv+7M+d0N2uOD5jN/1hlcdbfnlK/EEyVjo432Ogi5jC7RCapiEHjRgl65uD4M3kRZ
BOvPnWu6EilRbaPhK5POqo3DdEjMLZxBdVr/qXXgDA06UXl+NQ97hwAJCe0ePrAJmefbMaTnq4/n
NzFY+4+Pom6RDJQHbMbCH6RpGgTd1DE3PKO1uDMrsNJs+Y2w9k6wANpYmTPIqOZvgJX1yNi3Goew
F2zoVdOc0B9a3vYuL4lAFXiI7GKH7do3CaQ1US5w0zxtKUhh7O86WlVXI5mwIzr5G+BGtnMvw4WZ
Gv9dCXFyB6h6z2eLp1YSdbLMBhNPWK0UUzJp1vkktG0cW4oiRJdQHa4xo4xqF5HjoTbTAyIgQ8iu
qX4j6Bh6yUsYZSicujRnP3158avV9J2nKbaw0hjDwV1LdcT3pBu6ArJg3SOkkpqC0W0O5CpgeEzP
wYjOfLnKpMg2U2TLPII+hF3vHYUE5Np/FfIsxBricDO3XK+N05gN3O++2pIyLdOyCT6K80aN42Pm
slyq6yJE/qM5ZIt6zhn+XkdhexYNtRFItp5icui+0MmCA2LeAh+vmmuy3xXD/KPKvS2WuZdsalQJ
vgoODUskuDRIAPSvRuReWMtNrkM3qqRJUG+MD1PO8UHr3KmR8IxkFdZtAhl6VUhLrEjI0p1T8G5i
I272kxKBruJBeKz36IkQl2OomD1SvX1rGsx+coDx3aT5bckWR516pcOlknvrxyD9DbCpGqlrukHj
PJNlPDvjyZAeJ0uh+ykEF5dS9GGRsimBCCGPnV+UR+3jiro/wYioA24X223exp0Oq34jM4FILa5/
pKmJFGIQJmX6pXQayqqVx5Nw3tdcb9p5PGFPtOV1DoqmyKlgyJ2pYii8fUI4xk+kC2LJfDmVnV+M
UjCNcNQmLR5551kEIO7a+0hKK7li0HtH4FjAri2Dw4U23Gi371avW5M+SehcecHnTGnI3febG9O4
SZGiZUWgi6XHe1hcHEbyiMBRVsD4QXmQ2ecOMQ8QRdMN9o93IyPTmz3u2kuRIZhSgtrm+m8cJ9XM
YHvcaioaHVlz+fq8HEvP1o+dKTSCuds1g+C+rHWIka1sP6PNrry7VX5v0PclQAaOjSPCDpiZOKZv
kbY6eQBSgJU6ECU38+XUUz+UijBKGWWZsbwjOCa8rzyuuxBBjAoRRd2sRz3rOYYChwpDB/H3dNW8
GTm2YbL31Ovr5QZPEsZWBZ3lkFsP9HcyULvx0Gkwzolw3ksWDCha7LIOkI/H3WQXiFcltIMkz/1m
Ddytd0GjQT2IrBkr75lWd0HxMkQXWAAhUmn5cH2zPYBJrT6zIkqbKTzC4rbQAZBo9ebKsLZyi/aQ
yFLPiIot1/eF0FdTNTSSQ2M5PPo7/uEcz2+svLHhUrb7aB8LppnSYcpzGsiCN3Xt8sA2bDfpRXL/
LJ941dYlWxJIIwIzpw5haiVdP57woq3IKVv7H4XE/MXuW2fMCfa626viaEf34k6AOj+zAWvpR3iC
EDrfngdGPUjokvvoDRf1jrdLhlSwPjk/XQVWIuZgk9Ygmq5wrb7xF682OhD+DGHd4+t9Gae5Mhix
x323hDxvP+zrXZixcy8WVPv5dlQ8miE8tepEUvzP8tPmPgiZMCzP9W60ZSw1lr8JhQnE6PSGrjGI
WS1mnvMh644nHhCor7/PfI/AaIfavBJ3U8q913QK5SD4IVK5HlLl1gH1fA/Fc+2/3/xjMBOEvp5s
KE/JR24kZ4tV7aNHt4u3VEAPXSi2mAqsnTZmTIndpGo6UaLizKwXwpuurmSeEErVyaI9uS7yE0fD
ttlaXCUwfZVvKpbqoX+W7sD0wn3frpjSpxPd/nGyxKE8aUdZmetxSQrr9lIJPegolZF4gzouX8e1
ZB78OzoLtwTX7PlcUVd9e3JSeilmwG+v6eAlYhVReFzjBucK+RUPJfR+RwULFuQdeKbPT5t1FlQB
9OGvmrNOAOld7b8cf68GhUXwDydb1v9YrVskm8iZ4BS6f5jZ3zWL0Zlh9BzCs12JQFrEgn8TMDIV
ZKJ2DkCVutQgZgY8OK6U2QJYm4DPlvwociAbmWNYUNbpuwIXthWLVSgvq4WSs0IT2mCGEH8wtdLO
i3D6k5J7YR00Uvws9IfpckZ4YX2YpCvgsaEYdFy9gvIDUwR9cwwnHA5a3U7Jia8SdZCUuZIGjI0Q
Ls4zJ22cHen4X8fCAJTJrhXHsKIvfWpwTb4Ig2UH2kIxU4EOvCXG3qwQmxr9fKVCvez3H1mgeMR1
xYlB2iAyR5+Z9hBwNHbUps12oBnRCxf3KjPLs/4SCEuiSxyuEcGoyA4WTveqfeQhJfJZBNnzPEDO
Unf27g2Cu6sj5thQiCjJFujW80CBYMf5xH6+sdzD1TOPCM1ZDEQ6o6gV+5zMdJAWZoqav0YNBAj2
XNN5duAPqhdR/rPhzMXCJwoan19q6oYeTq9iNdRUuGi/hz7ZSHAlJvk3zaLyKWydQ074VavkW31g
YIZ3XbUBh6xF5QqjICAEsJr2RhBNaluOoMoQsFXL3PrPLCcBs0crlAIArqS6aKYTUhazbcmjOQh4
WmwoCu0t4STmmIXIkIQd60SqOFa8Jjr2+cHIpn2uNR0BSPilncUZaYDRgmMMsiurRF7Dvd2ERQ2M
LH+fH6Qt5yRPuFizogSSQhhxkosEGV8PFSUXBBmAsbsKsQTWTv1tv/bTy5RTeXK+XwMIC6pefzcQ
MLo4onOWbLxHLTqRFFqMR8kM3LOtLlsR/Gxa67baG5Q8KatqzDwa4tuRvmflTAkSRL0ojlsn+JQ0
IU65DXguHMH6SDsVN4p52HpDfcMHUQoK4/u4B3E8NKuZ3Tg7DGEtTxxfLu9SXXf9V38PZlnD/m2R
X1xBU0F2Epf+6Qk7pREH717gbf47I0GAcqNyPezvXlrSCXub3f8uss6oMeOT78KHjfbNHpgcv8Ky
hXTZqluih7X12wDVcJeb+zo4jdsxDNArPrx1jQqiciOXSzci50Uj0SNcPenyu20Rcsv2XmOPYDWc
qj1H+tuIrz/nVmJj0IfmaVbAj3E1M8ZpmaYwtJNlPDetl09IEcOLz+CiAOp/dQvHGjEXaIXFGK2Q
B3qHwZVEtBJGEt4xsnF/MGaY64vfr1DKVaNLfyOlH7R3OnvOdzl4nvv+CjYJP+piphZ8wyLsu3oS
gMw0fFoJhl0JYhFncPxFZAJnBZMCkTwsA9jpIvDuOCyIANImTCgKnLdYpW2mndd5TDXAlD0BQAoI
xv2mQUFK8XRXmv9c90vYThVv60Lux3NwDetM+CLV5KyF3u+Mg4JBbnWTICIZl9Sz54ArpM1EyPOQ
TgfY/yEvFRgOU8XhqgCIJZYeopysvjy8Wi0onqiW4563pD9nnPiJzCPbgNoM4ZXebw3vgm/0Vf0g
1ZfLG+eWHOvmmbCwA0J/jZfcm1k6kRnMJGcG3mA8J9msf7trILHag6fFCVi1YlNDPhhfYmPaHDL0
5gXWKCp6UNx8+r0B0EjVsqxdlOE4no8HIBYdfX53sb/n5jb9My2mYVzlRBUtfU9dCeQq8YSe3FfY
gMIPxSakXJtLeOKOfE6szrRw2l6n3pxouD1LPAhdy5bgBd4mNI9I+8uNeY4kPPgi1FGhTaP0w3Yk
uZ2SRotr9roua0U8CCsC/dTZM027cndt1uFU/3cvWn3GD/mFtcunnhFhBy6R/9ls53wsU/0ybagN
kt3U4FMuM3rk/jaBt/UGIT2RMZn7RfutFafT/miBmq+heyk13u0Kfg/JgQNDAXfHQsQXz698ik5J
wsBmNuAW1Vq4eCt+eoO7mnUjKW3XMVZvKmBVw2P7l+6AHvMuuXmbbeIu0Cqv649rZSliPBrS5QWO
dxyHeeOl41ymD3XE5xirGAgU08eUPjmByXJDrn/dz2emZB2FE3HJdKF0v2X0kKnSJN/GJRNYm9eO
a0q8kSHMRp1dODbnBE7mVP1ZZqyV+Tc6iQ1KgJNexQqWBoqN/VR0FOoexWKfJC3XQbcBpFCpKWxM
1iEgtsXxuSvuxDYbEtOnfdzhI9SIqN8MUyWEpDSU6P5UiC1d/lhqEpMR6Hkl31wkQrt1lgxa1X2R
Uno4o3VuAlT/aR7dc5swVUhG2qyVNrCQaryWe0Us52Rf5TovXt3M+3wRrEvOtHKuSh4GLFATv2gv
/7Nrf0CRJPg7BYtp+G24HK8lnsrTZxcx8p5CnQ9fjxZ80EgqURh7Q5yLINznSLYn8IDbGcRJ2ACw
ThvIFwWgcPAzm7gf3SL1Q7CGOxJrtV5LzI2dyFdRMenG6gxk61BTYwVWIr/QoEXsVuVfISpe2ZCO
N886gZEjMAKf3Z+oIy9Jk1Iihps0Mp12KysdELYTtGqzzpQzjddgsvnb1qYju0JW+jp95kKXqTYk
1tkgYTr78ScE9RprVenY6DmPP7lI5+IhGI+6OAyoBc0+ShndsXwAdT4MN98EUKEsP5oeC7HBCRvH
8FU0wpg4WcdtNI8jisbgKnDjRzGcv6UU7PTnBM4gRu36HV7mFgOjIr1AKFARZ+MRfdeTIreKnoaX
iLaHaVW2oWQc1G+0QFViFEs+rGNqGE1FwgjMtGyGQyrkDf1/qYE+89OodTHVu2OHxtaMq68OT436
K7x7cqINHWQD+JdLQVSHcT4ioijG3CwMrdiYAH0zRU3UeJPeVHJJzux7s6ksy5RBGWQ7oC5cJ3Tl
k0t+f93o6ZTcMt1EeCG1ja7K/Kvf6Kn9t17hhRoBV7vqR1duMCr7iUMjPlVGfQrv+TtLgFTABEr6
xtbNSMVCEo09IH53glvYscFWbXOCV9NNLFb2mxeDAlIlWECyiFEgJRN3oAyMIBoJcEIeCP4Gu+v0
7aF9GdQJ39BnBOjPJIRvu8MDKvOxL7WVh4h6vr/kuBWyHeL4TwczbMhe3STkdwk/vlSIcLgXJKas
IFZCUxiQkzd5lMCTZiIPBD/Mhl3qcpXqb0OyxCuN/0qx/p8XZsPEdgUczOMZ2GWDTZpf99InYgrh
VsHP+Nugi60S1UnTdJ7DOnVDDO/BMTsXdhNg4oUtIutojwiOk37CPTPkcWJdcf43eNZFBm3TwfSj
f/XSE9XBnIoCKPavRpMFivnZZZLwAJ4kl1sW/pkfsbnRzsCUUXVfhYlBS/YqwVn6pK1fKA/LJyG9
UUCJ/fuzcEPlPagQrIzyLVbQ1JKiGyeiTP44HjzWbcp611sRYxGQhN2YgE0yXj5Mc+DVx/nJyfs+
RyvPXu/2uQ6VJz0ieWlNDIig0ZUY/ucvT5b+/rx56BNY9tvewyDga7TZfXhISPleKOJ9iD05ixvQ
nMnpLnzadYci6VDB8ylaRJ3UBYLyhsMl5LIyO64H/iLC5E9Owt1vPhdZPdd6GVpRlOylYeaIYGqX
YnUpC9/Oon5hGGZsScyivgjujCYbbHFTcEnA0hm9qlZIogFSNhkHMB9MMkzoX6zsp1pg3nv/WU20
cXFsk/k027N0XRl5t1cURuZFFG7BDXTWeEyfKHle4dxUyDn2FdMiUqP2m3p5f1uCAJ3w6+w6DY6s
0pN+Y4kb6/8eNRF8ooaooOpQ9yteDxxSuctJsPGw9s71iTMQz8RarkshXFNiRrRZpnIqJ15qjQnx
6cJhz55VR1Vy+uSi4dr8BcLUV1WbmfyIkwgI5d/UO/kuWyIt49QDt/Kd29ZVgZIxpXtTAdV+dPJ6
q/YWxqC9BRtI0SZnui+MQEtPkgUk0Lqapl3gwjyb34IIlIwx6hA907YqQnQ6RAObVnhTkMGAbzhl
m4c2EuLq5RT2wfkSLDBGn4Qhdz6JnxoPzFW0rXeRaxMgnJaZbbH8QSvDQ1RUY+NtjeCeCFeOGwvq
R1itJwlpz8RnX8hCG6y4fxbaA+tb87l6MeqGnKZFwym4ikaQArLtsPpmqNZ6xLfKqeZJJfS5ho0O
ZDwDKTkh7OXrEagFuZakDaIMXSI+QR+eqDL9bI8e1+gFGPz4m355aKZ1VhVfXh05NTpklU4bxk3P
Rc9dsawXPZGrYzp8KxwkZ63w2gTxv2GWJSIrBOFdPO1g/4+vVO3ZS0G6Du1cbfwuH924ZSRrz/bc
910mC4vYn0Hq2neUaJv9cuQWP3+gj2LdfCnQJPhC9XgGfGvPKKQPsIsg4On6fhqLsJc+C0ecwzSj
mGVLSZIu9OliNXco3FGTkPiS39OgH0mb8QvOKGLaVnoHZWJivzZDqYPWmjV8jn+/5e7zXGfNNqI9
aVjFSq0OVNNHsO6KKulg6ZDmUWD59xozuNeo4chWyEhV/YCiiyZiQvoglsH32jrZnd5OtjrgM2jD
MlCdYLLoRWl7HFKFC+5UtJPwL+B6R9380S7/+9vBlUGzbohl8i6P24NgxhQ3htmWaLcrWZ1nvwmp
312IhWQ/Nvd4d4eLLvCyTGYQV2SjduvIlI+SlTn0fANE4f+fVD/cUm7kK0RSgr2HzYKc2U+jQ0uK
iKchOHPsGPyHNm00qf9dSZhOyYiXVo2dCOhoHKAL5a0cNd/ELV4tlKOmxDD4Owtq4u3KmiYpGEh8
4DftEWEjzIHiA5UDMPVsCw5hyI9oQiIvo6RDB01rwD/nuSX/gOGNCKX+pXcJGWOVEudpw1gDSLeZ
Upk+xjijqcpBaB6BYpGuHWxzkUX+owu3jKKxmsAAmg9bvNNQRqdcI7z5r/+CykozpWywYwmlWszQ
rKMVGtxMUxldcyD/PFd3FPocHooBYIvijeT0kKPEaqOoZTIaw066HsqMl6ks1AR3p1WKhFMjjsMg
Yp8cIJdWdQcs2kZDg2L65dRz46O68wUQ3xhmWnILdIgWGvv10YKcVUIIcPjBHv424Di9Mhy3r3Pa
xEEyefzVp7SDzmCBGXfcXjf4DXqFBPsZHbDSX3LMxbpVs9Lst7j4k1AsBY9Rx72RZmD+/bIVyZ4a
i7EJN97jUvSA3IDaTT83oIZp84i7ixCUsKilKTZN+XR3KdCl7G5PusxvbDvwxSkCc6V12T72PlJ/
1N6mL0Wk5suAf5j3ZzP+S1IKlsG8rlSpDsGjc0wZev7wND6m2kfu5fw2bBtjJPJcThFJCYLg7evv
PTv/xE2u5Oh51WeLrVG+/H2kg9SUvnGZ6aGKAteUtQpnuUNFast0WT/tin9/VHOVOYNbNQPrIoX4
Xccoz7Z/S1LHa5Op7cQuWcGQtdbrBH5y5csRUN/HJC914CmVl7I4xVemHdwraWKx139eSV2PgN+2
UpV7e+y5B4z9C1bkL++bnZlzSnIANiu3tGZHynQpoKj3bxwoyhyaVIoexvZ823y5Jd/sEVPwkV9Y
ege27Bd76MBsEhdYFFk/SsPyRRgk+qMu5GEcyFK54zx7fzR6V6/g4+cSx67nMEMKbw6RtiDS2hGJ
ZbiPL6B2xvbI4UxEGa6qT6uxvxedpteKO8LA0Ey1XUZjS8FdFCYBjs5Wm7pgFlC6jmCGAEO+3K+6
cOmeNqTqFlH8/mxbxsVhTOSbGqWfJHhIgBfZ+vfw654KwZiUM8zaKVk/Zh88sraE0VD4t2/jH6ek
hj39Am6+U+UnT1cjvOxQQJ+vbdqUPx8znVVW82gPeCq/5q+0dRp09bOwJvuBiKkWjpOYiYCXIpM4
cq4SxSQIe1xqNtbTFDFA+G4rUaDYlNQTl1Bgxj7HfRpWJACSEq6/A9inEIXck/r8bJ6R9hviCDRU
zP5paPNLMupVr8MQnaRWR7F875LhHxG878jnqreUnDbagq0eTUXI6ZxZ1wO+odxqcqIh0IRzxF4N
OzDL6n151FYXabzLaBZhDRKBwaQ9eruWOBsGfp3idladCAflElCqUmfH66W6IueFw+VHC5X2DPx7
T8+/eM/33mZ2L9Na1HyzyLYd1vzorS7zA1erCdF9HxLK62ry2uCTcH6wGyZvzmNe2eFAlsGYeIil
+FA98x/GJoszCIaKKAqpUEf8la6FMQGhFUXlh79RmwMawAp+6kNRuXe3PtHsfT4i1ag+xewobLtc
8mOk2l/jNPJBlq7+dd8TllMwuxemdIEChtno22CSFEo+bGpeBSw5Cxv2ZoRkD/aRcnKDzMz0YO0g
JYRI/VWQ7iMH9FjZsep3TFwSJxgOgvq3lk5rsHG2n1mzackNKfeAmLdy1118W0pIfvca1a2n7/oj
O9tznOdsXN6FCbLRWAgmvX+uJWwHUwW2dO4jNaaiX/lnWTxjUKuT8f5Q/VxDs64GBzrWwddRl/t0
SAByAVw3Fk2y0u5p6RRWLaelg4geydq/NmJaOFfJfgNO6RzL7mJBA9FnI6xdNVdki6o3gcLGIwta
p2cN1JZ7wbGHh1vEaWleHzEraqRPgC7aIiIDzlVlXdtRwToevrjni/qCQFPqFFlXvGru3mJWnjRe
JmujYHO2Pu8S/oNeX3bAD6SL9hMjTFuF4rM7eFJiMX9G+yAQXFLSLGnQQbY8LZnMkeMLwowS7ABO
FWPaqk5iFptWe9OOeS1PWI0SEemf4Fk/2vruXT4pJQBZCTKCL2MAlPHMnQK6Cz1694w+ZDD+RAVk
fowSdP5t7SAMNdDyoQkZvES+gzY8tbsauD81buV0SFtURHHLTOxUvtk5YiwC4a+YXnmQ2b9k8GvT
x8CcQs3vQPveWG0FWpEeVzxPdMBvYm6KquTyuTdhF25TmVsd7+YAWvy833y+CVBC5kYwUT4ktXqv
wMUys0BJbPyTfnqp9w1B03hsWRMKXot1Otv6ZgSB/ybeglr9YIEhlzB7T8zByrAR03UTwLGIO9vc
0SN3+XFgsVepkGp18NPmgMfEHzIjLZua6vaxZLqWkU1z9mKcOERpdPwBsGXhD6f/Ue3MXrmjNL3j
UoaqSc78E63CTQDxYJIAVlGU1vl4D+LjpSn0iMN4H+DNXdQZe5F/murfKtYXKZ0xT/ulOzCP44ep
iU5bT0Rp3aVlNB/Tod1eBDI7Gev7aILYJsPiND9D03ejpsaLf3GHol0J80oUNbJp1kYUGcw0kPGO
de7ZGMDn0lTYZbk5DmDmvrvOyIfbBt6CKI7PQqKsIX1ynZcbw+V1ErDfJIcmafZUvN0zbAPFFEzx
ASIZAUfNMh7cCC21UhFScZSKJh0rINk5Qok9nu3Ex16ADek4z9cg9cf2ao0J+LzfsrV1kwnGFY1M
LddVHsHu013bRiZ6W5azggnPV8vlxTLLhlX2WAuSACXNceWxxBuWWo0vi5v+IlAkodOawRScRsuZ
HdBoxU8u1ncqPcE6vOnarwPxCS2rweBfdOtSn2GsuI/wyLRlR+Qawdb6EECc7ZhcEvX5uf2yXgFt
PjDRPn0FOX/aCM4dTroj/arhGx1B9kih4XfnpA/lyRUpJ6AnHK2FrlHM80Dj4xeHYjw1mWsTPsDP
uEInw8MPfHCiFUNWrRqTDgkqMcnpFHkWBW5vOiB0GW/lltmIxOmGZIzw7YXAyI1C4GJ3HJyR1nFP
3ZuBtKnfJC2/A5HRSPZgvQnQqxZLrYgKzauDfqJrX4smzyJjnjuAde95YPS/Q8xno1qSQsew1gri
/JqTGceqWFh6k6mea73sLT1I0TdroCylgpVqTqDdHGw/JU38UNetrYR9QayKbk89VlwRS8VGtOzr
3Ahb7i9RTQFgBMlSZUrdTEWTZaaPX1aISoN8g/PYF44R5eFK2MxEt81MZlTpiitzJnS02hyKSdq1
FcjdpfnJlRXkBLvgzpSpHIDi03UVgcJUCB1/WIvwsXu4B/81Wgbj7ibN/qYx+3FgcgS6HZHcPMcF
B/+I/DPj/W+Y+LQoMh7od+wSmX3tYYO0tFEBcBkVyn2ritCUmgyBSUqTvnWAPJsmYafjWmtnY2YV
5JKYHUuPaxCseqcTkN2tUOaM56/voMFLcQSNxbw7AN+nWJg3EySd6BAAthAUhSY0cVTZERXKPiR4
9OPDGIzS4UFdGO6dphp9SxoDQEKwW3n9lrgcMdlEAqms2I2PbjQK5eF189Zt+7OcOPfN90YJLxCF
H4yKuQO1r87e1JgOW9WfOaz9IktaQ00wWWmtUHLcwV5PEdhmEaLEX1h0NbcjXkhW4qfiLG5zDZOE
lJ/hZjUcL1WBhuZg4WhRUqgOdOScR/BSGxSNcK/8fSFmctPYcwrCiFI/2Ic7P6Syn1nxJXcyhDa4
qCJOyJgCeqwrd7ek6S2Wi6mpuesl0CAY/KP9Dw/hBzLpEzLP7t0+fktnlETH6stzTOirRQcir2tM
hvQsJz/TiOIRyG4F0yu98I4ackdHyo6CGDaT+QlHpMFWGT+eW/Jt0EaYdMAbDEGNZPGZ+dLCd+iJ
68zydL9R0UpaIGTFiL9+gObLLpXND8w9NGZpfTqB5eUBNbO/iR7SW3m07oZlJtADl9q0YEWrugId
Fu8e/o1k0YtNfq+fFMsSS5SeJ5HCxJFOsjFJ3rXB0Nmo0FMvO+nkrp/f2p966ZSx2SR3nOqLO3Q8
p7wHszJf9gmnAu4N94nZQByHk4AEquuJ5szcQGwEsc7SoDlGNn3FEauIr6BPyFRea+JfGdSKKDbx
TVsBhrM9p++h+iTcR9XrIixThITgd6iyDC97OK/SSPzcvyLISlK7m/0+T8pk22eGhGK1Uu//o+75
k82jYpbypHZUGmvFPS7GzQF38eaqo05BnR+6X2t3gLraJcxSX9Z6ZTqEG3fcBWi72jHhwcyqY4ss
O7AaPXF3mJftfLPqtJynjNml22b3E5fSnVM/43eAC+pFKAkmm6Qo4oiqHdf5pTf0SFLFdoIa7yg/
DlaUVgzeyF0wGOzRYbWaW/bosK9qCfPc8F2blEiOwI3YlwGICX+2kq2TSWm/vi/FV3nHoQqxunco
8SIphL45zj6KRW64ZwSYqRIl2diroAKsFjPWh400P/HwOJkrgQ3JS13U2VHes/2jT3Hkv9thcyAM
44g11cUeUKDmRz4/HWD1GoQytDYhn/XReUxrWNcRin0RpaG7B4UO147So2n6e7EsEEfx5Cyyfnpe
E/i/B/zHfX6+fxtPf+rmghnrP5fMu0gOZ4+iNuD+1VHzLMDcY4QG4FCUUEQVU1Ws0Jk9gURVCpf0
hXCEvzrPLmCGf56AIE6IMtxN+Ln3zRUjks2KKTBuIX0/wo74evHDNEh1CQp8jZlHkBn3RHCKvCRH
HvsIWkiskEHkd+lUUOHHkQuek9RtDukWNEVWYkSsDliUISxRUkXseX+1eQFUWdoSyrGhio+ZdrXT
9DEazjMB/wiAdCDxhhVVzUdO0l37EXqGGjVEGMbJf6FbFVVmJADR3YReo3O5XEIS+AAbwoyFRjpd
xD95S6VjA8LHnSMewhHRXmGXj3E3l5MfnX0G7elLy+78E+jWDMLP9FUITQv4V3gLxGDUMosJYrmX
cuouPg+RYzPANcaYgIbF6FwDHUg+/wH2qU5n5waF4I+w/SIYtojQGpsFbGtA+f+0i2Fz7xomC4r8
cWB7z9ZPzbDQmwBQ4KfCvy902oAuDR4zMAhUqblHeyshlDoRU/k6NE6m1kcVFMB72c6XFLqeCJ8e
g6maCEiQXik7orHvGE9dL0p7jtqNCcnW0qQeTR2Yjx6lr8b50vQlMaVIHNiLCgqGt2+plTGrA+CW
5+4/KoAj7aQvMTaFeqNfgKrXxFJx/M3/vRzC5GJDSya0Jw00slHCi2KJUWZAdwuV3hggAYIH8Min
g5fjZg6cyyybjWwDCZ9532QgCzwf2ezUvvrKw5zys+rK2AUiEq4DAP+Wf/A+8C4cvJwwFalROGlO
P3XJ19ubrXinNpju4w5u01nxv0d+E4kLTpelhuBdQCWp+OL6pw6a8qNuxkXok+RSTcT7fgpcVgra
k6aa63qU9zenG17ctWHub2+DwzGsjSsbLS6/sqnWYK8n90/hh+cQxPZYDxkOE8r3I6CTg/bT+6st
xtPifBjhAT2Pb4expM5PGWn5KWt4HMCSNJaKNgnnaAldypGKqUUpbpPfD8PVRtlrtcok/vcbxLki
MArBwBEFBwCf+sDHu82vReRIRVMVmNcvQLib2hgzPjSyWK/OxVTVFM53U6On1QFxHLZFIZUYmonM
nW0t6N1LNq8vrdPTohT/ev7REg6c8LV84IZVc81TBQ8nLl/VMkXBsqj42PYn6pL/H9PfvKKBSEPs
RNiscicYcaNylfld9g04lz/MItFsn9581SKpuT8dH5bS3FLCxvrWpRDTOILSCBeF8q8assu2JIRJ
vUnhmru5ZkVQcEAa1+QvanevU97jIzDJRwmPA44eFyQboZ5T6I8hOgP9UE0qUTYwJDpajgyEKVt2
4T2XRqHYofTRbbsQt4Xn4ZNAWOa3lSaXtgDPCkZMq1F6fIyUhDP3+eyfg0aNi4llNfGp5co+6twa
Qhd2nOm+3QmYt90V6iCJ4C6VOZrMY83iKrYASLo9qSUScYkHHrAo1Z+TNgGlwGr//8Luffgj+64L
yXCkWXUyUAUX8+3lYRE2wzosVAsKsvM1BF1UOGQgGm4PSqrS6UZ5OMyMSeQdn0nQcX8F9W7tPmkB
hZd8sqpV/REYRQCTqRANr7ZgPY51cIroiKbgj+e4PInU1ylIS95lIlD0BTwI3xT81VQxYsuNMqmp
TOs9SEA57FkSOshEUniHimxeBKvtTn1PcD1G2pU6UuIhVSPqlAfwAcxdW7i9riARmIap4e+XhB83
Kke3dq0w+jpEmPgS+Pym8FHT1mmOn87s/VSfsbKSz1lypF3bU0kAKOfepuRGOk6TYSRqkkZnUBLr
Nn6DTDnwdbolKK5WamqQbKswCXfLqDi2x3ynTH818KfDDywrmJ4Hf7ctxW/xv1pMZpCBE2+zOSdY
7F8wJexPyA3K6WejcYUT9DA1NQnkrJWz2eKP5xHlV3EEk3ULs7+sI/Ro8FjNiudJh6q1dGBPfndO
UFIf61vA4aHOwxULNJtVLdyxmxD76hun0FffU9zZOe5/y5jW7yw1ROr/0YsVoBNFGIyc165cTIaj
ODVedyXtcBBnwoohI4SWvzbnk8bTVHn/AKVjHroky64Kfi2NHXoptF52Q9Lp0LcUa8KahUNcDtj9
Q83cRw8g7QjxSrhTSYbtZNuIwgYhOd6cFGEnsP5YCEW0CTyLj16vDB13Z2SrTdgnYwZ5N1QDaZ/E
53C9aPRHQDAbEi8C0G5sVFtemS8Am8uMThAs1zJX3ZJNNnMCwC1bewLa9AoFe2FHOgerfEBkxJJf
mefufru31Ffuhx8a0m6TZqUvyDiRpvp5U1CWSUkU1uQu5ujDIDV+hB7s23mYbi52RbAPi7iuo8oi
7PmdVhNuT1Itoa5ipFRB8JAgiqppzOo2H33L3BZ4VtzNXXBcc2/DsOWjmDiiU1QcvIP5/TYaUh3z
Wi9y9yzcSsU50lFOk+arcgbsZc3fQjvZjwTlCtSDKdKaB1CK0j1YUE4ohcTi52VmVrpgl1TzfcZb
j1mOTs39ss5KiGQfE3ib7Wc2fKzXsVTRGHpx3ysZXhh0pcesKOWKgCAp9K3mUeppwHz74FgM95K3
vHw73Va0+vTsRzvPYElbwr/P+ayKEkuMt2SMxcf5ymUoCoKFXJC8IRYegWkpspgNs/MqMwEBJXP1
qu27aDuEWHYnfabuNbuLE6kgPYwOuV5Wr3eMU33K8UwW1oIoHhBB55FogNbdmYuJcEeFiMtdgTJI
buPH2K5jxvAuohh3B2giC1uodlBD59oryS6kmbhWRBVORLnAMpU4Fik5jGV/QPnujHk8C6CSSh0T
uPseroVR+G3rtVUyp5N0yNG5rj7p8RH36yHZZgCzZzaLHsZhehzOYKvwfauJGRKb239Ky4RZe6Hs
WUN78PB+ldGjimvlEESuUvsxpDwsY3azAZM6ou+mlQfWyVYmd4Wqt2Lp+tYXZX5LtboYUPWShLT3
MOzZQi8PtrqYwA87uHHFnyfzFgOROfPP9XgMrx7jjsx8VJU+NcyWHdfvR2Dmrcj7+X1g8mauw2z3
utKoTd3utbt0koJjExz0EyOYA1+Qs1z9TNSqem5MUnyT7IqJSz7BG2Q779ouP+EYhZBOCnkYu4Nx
9kBOcMQ0wuZ0WW66o+Gkf9M501A2qHZWLWVoIoWlPT0vBL/skKvqAMgZVZOYarlsd6UtxmMJ9OIg
DV9ND2o7qyH5Nbu3QYV6GTCBrHkGXwcFMfYA+Ru7TJQaMnm/1H+oHKj1/hg0pN4e6j/LfYE9w00n
C7eLFi/wjMIcq7xJXc2ie5MI+7lxxbdNxPG9mffsZJSjAt7IekfGqhs+r4ofBCbQndO6KJtVvYpr
VNxYXK+gX3MIcnBvVe1Hq4EW1ojbkPN9sJ4sBS5Neg23KEYbLVeZJci3FLe1+YAE42R2NNcLx/Vx
cs7spt3Qh+fcXuG31Hb9SDmPGpN4SUr+ylQVXqQCj9HCwy64LbX/Xb1OSF+lKXmTF2PB2dtrQ3ha
DzF8PMO+hWEjIP9fGWhjqXimADtUWGMMVE/1yFgwiWxAgZ2f981k6lFHvgQyyxQyj+I35e8XdOm3
mpRgobnNWNLQs4duSuvVFuMRivdXcAFN9WLk7RvvAmXgDdvm/z+GR35PP5CnSzIWEd6wCfi4plGZ
FJJnTrWDLCKHFCrV/pA3mKxVBmesqE3H/0U/H8ozMgQbXvEBP7U7x7BN6f+IDZWrq0OYTWUKCoBU
c+lHKnU/WZwqr30rXtoWfADfKZG3m0PJ57nShxnWaH1D3Va5OkykPyDkukta4Rs/atk2G1vKP/wG
GHLBpSWxYM0X4tAq2O1Y2x3J8L7dnEok9GZ77e51oPwFlbLMYk1Mr0xCN5LLCRCh2xIVJDv9mDyz
ZADSpRnBNJEYxbX+iO++bnwd172Z6ou1yv5/EsNT6YHXyIs1z134Xia3scEwXrGLlS8TFMeescMW
pKCU1u7DIuuIYRRC0pR2FEotke9Bq2s7tj1SoCyU3Srf5pF4r81HZwNl3EbkrSVDfN/RmA1mv2Y3
+0H2Ac7+sJA21Gx51S9dsJrrnK2Qi1ilLwcY/54mFihM/cV0UwtOsnwHKsne4aUQ1D92MEkfzGTb
JuNr0ZrOFaRmZdyacLgMBwZdATaJtFoPrTXi93woFedjSTFs1hZofRmr1B2gX9L6HkMfyNycJWs1
wk3DyKE+GoFKNVfFGnRGDIqgdsBF0eW62XldXL5DbcnsAncayNf52wTUxpTOCAunU+Wtqa5u6ODL
LB3XLrGnnQwtvJuWJt4+UIXXl1J1FTV25FOjG9YDB/iO8i60xE68JA9hX+3ETrtBmIZ2jqh61YJt
YDaBrqCefGkJ9a+NgJQxFIQMGES5CtdL2vWwWjNTB7fvHQYNelx0pQ8nebfwACS6QCNikQveYa94
OwnOqgfLDcRn0o1T60dQsDOTJnpZe/M8ThVjhixU6dHeMu1IDRYpMJW3f/4jRP//7JF3O7wHicYy
ia5ghv2hxEONOxmgfdtEVZe1ONiTesYPFmWwz6fcP/As/CIbg3HWHRYQrFkRCgGh5MklfIJCs+iS
uDlNyOtgd/tSzlwdkKrGTc6WYXVkhjg44bQ1rKSCOTYIzp3z83lCARkicCSWBUzN7zYLuTiwGZkd
03L42NFG07M0vEoUntTUZeRQBwN8CaVMnqwnbmZKzdOlo0hIlPDCTE6+UQnoSVfsIn0CJpBzUEH3
2qg/qsQAC40w+grahXv4hBtjeTiJ6ZOK7gl5UgtteBS0Z03Y8U/JrnYnf75PA7Rp8RwyLEdYu9Vy
ciE0wQAYaoih+9hVpPftrPZVvZP0GxAF7yxCTd+C8J4t8QRlwQRM895mz7kXS4YTYJjeu1v6G3Uz
NxA2KNfsi0BGkpKdvjPMK843eBmMDkY82Z2yZj9/RhF/K0Aa44liTADgAeeKIAROefz5yCV/bEoX
9KdGxCnsNeLDimP0an6uY6RJnlLBo4F1CqqR2VXg8RP2GcAKRvlfq/XqgVgurNGbbXbDK6lTxH7e
ougo7BiVQCuVmcMC8k8J+PKHR+oDHdKXfC4etlSN3BQDLRsHXOjhHIcsAmwlYlN0u/mhotpMtk5u
t+R3yJ7MOXQsQmci/fYP015M/IxIdavffkmfIb7pHtmiwEYo9QYfqxVj3Hd8OBT4RIW2vvOfcOCy
9TvCJu9rbOCz8fmb9n8TkAVp3fUjTuRASCj3aHrFYbLM+FL5VGonxT8Ol9za17EumjVmmMF+GKzh
LDMpZPNXHMpV9v7KXjRlgxdRRk0UPzIvteJ7j5qwM3Hv5DKqPtfYunzKFXHXrqNt6iZl5rZvzJe9
2Absah6h1zryyKFe46EjSAWFblONKnl3WcWlqDEm0LU+mP/yxizNWn4Z8zXRWK+etYc0T1NZ+tms
yn6NUARn19dGnC54UpSgeU931UlVuREUkohzwCoWLHiwSbsGXkkqgdPllsurWVa358aRyfv5pSkB
MAdN8kt9civz+TV4s7+ZqhObZGA0fe4ZmCDY7qNnXdmIIfKhLiaAsZztwnd/4aHD3ru7rzdLiE5l
rGydcQErBH/CxT4yeeNYWeuV9XBOPPPgUoIyd4ilV5fntdUJ/ejGNcn/B2ZMxpAA/jjMO+1r2UT/
LcK7grMbIQB3zritMSwhtbcJ4TAge9jt3awAT95xG95KVG0mrQjvgff2ac3+HCmAYiILXXnXVrXO
9r7oWmknD8D6ukwQ27k552hMwvKu8LJlcRgRC0xaYn3yqYRkh8ZS8oKr7N4bR8RbrpivaR9wRRbw
QrJcB6si6we/VC2ly5F3srEk1FSEWx2nTxo148TUliCNIL30u8n+hOQGgv59vvuatA/q4L33Shbw
3fps997VMnA9Lj/3qaOmx1W3scKHfhlDxaFTjwW+ULi2ZPDzc3Kqh5F19JKQFnGRfdyWn8TTUvVd
jKh1U+v8YWumoyy9MzGWgDlamPOLzqPnSTFQ+70p0r5cWIqgPcQ/u1YtTbNbHdnT/43gLi9vVkhr
7AWN58rJcKxi8w0rpeYyxbbccLnfNwRNhhp2+Ma5VgdDWpLpkag81x9AIIUB4E2r4djgHSokIID2
RxbCwKRa+jqGzI0tKDKE2Q/Vg32SSZbNeMDCva0JIumgqsxbbq406zfNjmZ1jmfDqKi9NGR4R0P9
ICFrLLsfEfTIDmpfNxuYS4pB5aBKI4TCinEbfg4SaT/FDEzfdoSUQ8olVfF+XodL7DTf1IOr0GgC
9Q4Lb2aMY1mvC3+uuVBqTE9BJGVTLYINsiJbwhp1cliP5pNlVcYIayh/+ZcyjQkucu+Jyvwqwh56
5Bbh7vbuGAcjW0bNIoy2ylqmm7+ejkp4WKaJZ7Q0FnCBzf3SdzSP5n4C4YR3OPbYvaDieR/g0YnL
dKIvzhRQ99eU1mDOVl2klX/diZnu/KxwVlwPONW6IEVyDeQZYaFJI5DYkjQCVsQfKZN7WFb7Rl5x
W5SrNGnGtAV9Nc2oOPyK6E+jlN9vDejnC1F1TbL9qcV5PhGOVmLf+ihcg0N3Rm7Y40GusmvyMwR9
UW9sdiK+ENcXL5UA80lJnOylim8pagR1waPKYex3myrO0K2G6l+9OMw8Ik4H3w8xlmXU3hSnGlio
IQQE7w4izv5ITZ8ix1EApptNskM+DQYjP2QDxqWo+6B96qxehShdFxvAZcZlHGPBcvVodNiYKcgj
y+wEFHJg/92OpOBqa7CwJtxVRcIym8ogOhGxw2IXnGu1aLgMs24Q24aPoReBrk9ns34YQ9Vha+eC
2knZSKxhse1tH/jyD1qM+O25feTRzvxC/BTjveRWecaogEUjteI/HD415hSmXVOSvs5j89pNF+sC
C39yhz49p0WFbHoMMPggLwR/Ix8YFhd8rvATlqQ8PApnqfWRsixX2/9Y/EczacekweNGsPdqNVz6
Xb0myLVOLoyuDS4dCLsOORgHGa4fR9UjYGtoeldNeMMT4DyC0+LlfsBibC804hL+R34A1Piw9Cnf
E4U04SX4+sC2VwAY1bFXdHLWIzMNHmqTvFNDHaulzRz6uzR7G7g7nlGeaQ9ZvoCZNrkIAe24osrv
vQ73ff1BEgPgbF5IPtO8PQRhvjEXUN/S8QOvtGKubEWBNQW/Vq1BNa0vJsoo64KWzu7cJSEyTV8+
bLwA7/AcQtsBHLbcVePe0ofGdIiGh0zOdaE26hnf9SJ60UC0nSuAtrT4l2no8gY+HyKL1ZWhvW/b
H819MV1IBAGi1cdNDxlcQQJU1AEB+0juGtp35c7PCeJ3lmYgdefsw5uHLmL68z46sTfXnoP2xoR/
1ggn/iUCWa1tpEzpNuAnhGnvfIivgmqJKb+r3AyqYteD+KtCBeTVUh4VJu3MJO6EYMOmO5pcrrLU
MiTudFUO8r/1KVj+uq7MXhMOVY/pYp+h/4g+3cIni6EZfeaMttp2Vncy1q4dB6s0UjNq9gz6TdfW
mj281pUEuHdFzq8pd4631L9R2doG8VHIuVBuiUI5vTDRxT0W9iazbRm96V9ZuehAdjP2MKzdggTr
y5icCfarS+1IotDjTO0bMa3bZYap/GoqEX1cDB0PuBnkr80P4GxH+Gfj5pYlYkW8wA5ptJrqBJZy
JKO3RJNbb4dt6LwLr0tmGFYkyP61sIZXd8/x7qdqSTDofJ/zsy+bURhqUK7ZMkxkN8Jk7UtBr44X
5Aob/GkohzT6isnTUjD8AMkE68duEHlsZIBnNWxgFbTO2Uvqc17uZ3Z/vsoig8isk0C7jJvz6JNz
pg5H6VBgo9SRqNvKYghOHoEpUz1NfEs3wdXdQWDLKx2yDv6PdQkxsprKS5YQGP5sImCYu3Y4VO3f
5B5kAse5TxhSaX54LNXTrhdL6D+fnqoZ6JvbCR9HQpEMP0FVUJy91ud4lAHuEgZwqvvqc1gF0r7u
c9HKgvlzMB7IC8PmO4z333tcIXKCGuRqnZsR5AyvW1qnpCmj+7tzp89/hniWSUfTyDiIKqnTCk92
cAwHCtgieDJ7HqgDA8nvMN2AGcZDpA8Ybv3vVMMSuyavGNfnpprNAfT6D8iFpPFQuOYqyBoCjUM+
mFhofJnKiQvsy57JHr42LZ759d6SHdzEGnYtB1CoId8b8gNiSRz4Qct5K6grYnfwpZf8PFsVlQVh
IUgPD+2pmdgvlfU87d31iLBw9LtxhQ4SROx9cqcInHf4Gq/fsJuOvrmv1OLiCyh50nDhECkFXDVH
sso1lGrWESKLnvWr5ITzYEUsK4IKdPB31+Qvzhp3WvIFxqmGVRT2pdrcdTi9Lm26D7aGGp3LK59P
LsN07xlAdD46JFEp/FJO5FtFHVNj2nrjndxOVLmve0WHX3kr77BSrvEpSXtv+0R5OaseZoyaI5o+
12Tof2OTjY9mnqN8QGMqHKuTDTIaPODQCLkquRCTV4D+QfZmmCKXmWszAGl52mPaC8ewlHIf0H1o
kfS/L2HZNXA34P24Q4dkxJQ6WG+esMQQJCs60muc7PAZnav90Cuw+xtoY7epqTcSqY5yIJNWw79M
uqD2gRAIFzwGM7/uOM1Esz7PpqyHD2KiJ9l4bNJmH91vm7PNPH8SPMsiC5dZTZJiPE3I0o0Y5mEc
diMSLR+G9sAhDOjarfyAi5DLg0k+p97hBchQgOKrdQ050WzrGYmbSeQ2zHbrPqmg/C8M6+r80Fx8
epzfzQyYarlPXgqXK2PAhP0EaJ6Dak/q1SBwwgDhdXS085wacxCdmbLk7Ht0G/O0zOsj20fLXslq
vUD2DPMiDksvTpRma9qLNuLkCLj0LePKjeO2/av6PNIfpOsz6pQvOkXDYH4q7u9+yF3Yo8l7utbB
zrCOpM1azDTwgDuzOlfPR3tqGTz3kQVohqLPoyPn+GbONnYO1DYNYwPGBHmsiDCKiAXoR6i7QZJW
fH/rL59ihvUPsg7sykNnu0RdKm3cq4UgvUse3QdbOfAYGoO6IeZfTj7F46+jiq4qYKsLKIdbItUB
nGoHZOjPjpV450Y6ol48rv8PSY+oxl7ZCfJSgifAPiZBccB+yKq0QQWllTOG9dowFTxwu2OXnabt
lSjm7omoiX9PoapA/h/+g30uPeHGF+tZy9Ns6HKDsFRuU2s2p7QvQJinGuU2eoWw4I4IY0o8jw7B
hbD8smu1LRZY+sU92CasllgPTWeFqV1XK6APYp3v1rcfSCMqZTUDsQfNGC5WX3VAB/ETVygZlJXf
Q3xVHKthbD+56WO6ACTSr6inmnNPA8W9ziPib8y8i8AcsLb3EhvUl7yUtJ4FZs+DVQiRMWArIduo
jLsP+is7qKlEilhTLtGH8vXcFM8iT2E1bGySzT4r26WatC0c9JDSyceVWDaT21x/vxzWHITSH2i+
gxZZvm+z16zrPtQgmaSEBCGhgwyh5KzJmbFUcY6MxH70AZlojuDnciHVOv9ZFTMzCLGHj5qb8utd
dz+21fBkfPaceVJLjwohlqbpCXAnfMHHWap07VIHGgrFxdtxn8owF8D/nyv+OBkFsN41OF/BCvwt
J3iJy/znozSQH+LaDZxKmyVqUavdWUeqb9MhI8snYRl39Rz5ARvoybMQwSknau9CtLXWUx/If5HI
0o6isZLM1fSF1/4qp8yiuE/MSFYbPJucKg3FoUj2ey8HhN555rWfS4eBUzpnnX9BkfZfCnNWFe/a
NLvpv0/7oBxGT1kvnX5opjCn/efJjQzpEWxypK3SnsopcEFP5oqb/ld/WMdPG9SQO4oXYEOnsU/F
67hFxtc0HykLNlhm851HIEiBOPrMSPZMLOp7o0VL2FU1FFtau3opbKZloKoe00bM4WAp9LjcwzOj
NsUHrYRoFQAzIL1TWXjCZWC0a5WK92VFaB2Z1s5Lao5zIckdckp5jUhjuYK7Jd6cZBEhU0lFOKlC
kQDhSXRZ2uyDhRHugJBSUSOxHqXC2H2TJ4R8yZ1SFwh1HBJoL2SVmuFPkMgQVYWfs9TbJ8abIHiJ
JqGw/7uwP1+i39e0IF1y0ZyD6JjdHLLIwXFYfRdTtz2qVNcAKph0Ix1f+Wy39d7eSB0ROZHe2wWD
GB7VUca62iKOs7YRrWF8qn+TyvLl0RZ6vJm2ybgbjUDnB3heEpeTHrHdm2unA4CBphFqN8HVSBcK
vEfzlxHoxJMheLi5RZgBE3MyvdUASaTc50TeFk2q6j0nAEZaAqlZjb5MFUSLr2IWRaKW5rknl6HX
SujmFj9OBW5pB07u8PEIQYT93nswqLEHHpzBCfBcnRno28tAxpmRq6YkIECBgnoUF3QJH1agAgUx
EDjucg40XyIF5dSzqOJPs6rANWn3sqmlxdS0OlXOBCMQM3nNYmXeljmhcC1o+hrKRIAI3KKexq3g
0pvAQLqOgWUeZWYDApQ4BKK83LUhJBevQ3Ukc0XKaa8vQDiJPIsPjV/ngA3cVvc2ihYcgcw2J4KH
n3swVsTeZ46690shSDqXMyc5Tu35lnMWFSa5xFl8sEpIxVZ719ddl45lCZmHIrqD5r9DQb5avvXt
1n2F/soMNzEp9NfCORm5wnhMOVVrr8YxwHkWQeExBfkgFuxi4FbRL3gEMDheq5cBFsTjzB2lh6S2
xUXpHlY8xX/3hQ7nYzH23pS3qfBc0fwaR7hIzzb3P6knOPNKQRg7JVgs4EckR6nsmNt4j/Vko0G1
5OA8WZLB7FWGYnPrrJJCxaVXI26aFlpIh7pv2rBPKkFmVXaoEmLHPyICwkZcJYiveLOlDWTI8O+0
hlc3goFvOd6r47LAC4exZ29tLIWf4RYjhMe0oCL9+aJ/2vUrhkSCB05p+yJQlAGVn8hIDomj12MZ
VUJmzzPCntV62BqFYO6lDRn6F4Sf/FAhGYG43ahIrXxKuldAac0PGtYm+eodsQervfVp9U4ECD+4
0IjuBIycXUhHXjK7SCMNUE8gmS1O2ihDV5v+RJtmYSm1nK8U8XqmVYe8eoOSrjph5YZPp9q+4sSl
Y1uBtksym8SgNW4kYmhM2irdVAQqqRCvE7CglEVzoZcv+/ewcZX51Am2PFFxbzeEXDuWtmVHKxTt
o5jFYdhwfB9LMDEC+g3JRzJA/aUQ76RcRVvDYdNcMopHYDIhTyPMkHxrD7Y4q0cPK7GP7gDSebWp
qD92KoIPcw9VsO42otJkUsg7qBTKcmYVm82/ePTMaYkhN6gCKUXbcfEVBkw5AoPiVpoQ4Cg5HD1a
XIncJQOUpFZ3mbC5Zk3TBuGAWdh+enNJv9pR0k9JOop4/oOdTVUe8af7zDSzGRDm33PiQqP7RoJK
79svCHlysbdl6ohBPTcnodstrdsxvLN6jY4AWYPt4RK16IJUZkbf33QmJdVMQIR7muDFGTwWR3qw
oqcjSFTnIIXS744S6p8ZxxDdNxLa5zsza/VkppQAXUScxFjU0rVodbOfMsCexkPpv8wiIO1T5Uyn
VzHm9t6K+tNcpZVoYitGRSe8+IBAAly/M8zd6H0qJHGh5ZI6/70y2+oE/tRdneTBKcaKB5rH4KwV
cCKyOOYwxbYJOw4sG4NkvkcWu2pqO6q8GZTORjYquF4qB3Tuly4W/3nl8jHt+cVkU2bHdm6MYBC7
VGBjwMqyMAh7I260fGCDkszinlmm+Co7Fua0lbJRPRxha0oUwrBG5FaUIRsN5kqC5QYQhfSonr7n
1r8ggk/TdAOONUdARNRT5+5r9PD/NXwG3G+fuQ08jS9whJRa+0HRetUzWdd+dn71P5/Ixxw6bgDD
pG/AsD+KgdUXCFNkKH8k6U2dL7pDLbbZLqUpJHKU8PpX0rIvJ9qiGfprDGHiEIRUbtdck/R3jbbG
Ec2urc/C7HioewI/azthUqe15M96xLftnbpqSODR3pkdnHVeag0hzHTYjHgn+zxCNt3NkAd3sF+K
eLDpxaKr1Mvd4Th8wbdFmBwNalHKa5RgpmS+n6CQGNi9QSCh0fyTl0VCU6mo2gNbfIv1Ulr/b8uS
0qzIzWFFbMulzENwZIRlt22I2Bw4gAA8C2nV9UdvCAPv4nInif02vYsY2f6gjo2XLft9Yvf6Qz5m
kAtjOmJBhkvF4lD/umHz46XcvYpN86YFXVC6a5iZKiSE+/Adj8nHDZLB4D7nDnKCXC7m2iq9KZKl
fLEMpEDz7EslRFhrmG9COJvncKRVbBa99UmDca0LE4ihi7QtRjwdgZwzOAc780Q8Yksmj+Iwt4zF
awtTUHPul3bM+zewlaV6ZFTmgXRlCSc6z3z2ll3Pr62Awc0hgM8OFQNNOH2ZEmHzuU9ntJaPvhnP
FqmDme9NKQVmcRB3JEwSw1pU12mmPq0KzzZC0pC0MeyZZHE92aiL8JsBeF4fMRuG/PeFVxxA3BLM
tpDNUMG+ciKLgC69A/g0KgA2YyFiPH3JGTMJP31wYAtyRuV5cXZ3PuNfJ3ZzSPq+6vphPA4Lcuit
EtZfKLFSKzRDydZAidkrad+DO7O7znpC0HaBuQE3hm3Ko1+nTkwrIXQ7blsQko6P4EX6YQiliyiy
I53ZsLLFA13163fXEXfB6ePBOgK5LQHAMgzX7xHSA6QMTRt2e49ZlaEh++yqvr3Gk9yqOTsTlgTb
NKAOq6G2S90J3JMnYCF+07zdOZUeQjj6ggMUa7rpEGDngeRlDCEGyBvZuX0OpE8+QdduRBKE++G5
iPUunXH32d6zBRgm6I5upbHAFsEl/48kdk+oyFNWp2jLueJH2bJT4U2KscO3IBO0J5bGZXE8nw/I
5MUNySrLKLuf1W+F/sTB8G2zvVhgiV+hXsPC71grzCL9GaIFyAJy+3xDWdlrPlJOblgGaeYN8a+w
l58nogjSRyPlIov5H1boHjPC8/Xf4O4fglxQ8OrNH9YqC7TT26geu8p2bGeEro4owXg1518z9ysb
SBZR1jno9i2NLTLtfS/mXXnmTWTWsRghIW2u/obOqPskvx36r4fJo40rm1/yCNqB9/u3xiDnToL/
/uIyyHF3CZYxXmy8nWBrqJFxls0mKgNWk/FeNC2KGOl26O38de0qhu9R8TS9ST3dIfaDUG7dV0t9
cqZicbuvfFbWEYkM1fKmiZoKRzJYH1YqpZ59946ylvnKY1if71CahbEflY8OC6TyW8tAXbV+6Tzy
OUu9enuHK94CCSuxoZvFScKQrpCYA4DculN/xAYpHosjRZFWOOGLbwXQ1YwxqYNOnW/u6S6wU0du
CXhG4GmTaE9HJ8TbNqXG8EgspzsksU81U5N/IyqDW2LTkhI60Bf07k0vaWakSvSYu300JIbcgl7R
hpAXlxHLMcleP1JiL47uYx8HEtTtAd7wa7uE/2hb/WebajGcWRgnIDqYoVsFVb2whkjorS6ZXEWT
zA0lOKjEjPHSWg/OIG2DId4cn90ROZP0dHwdkZq+RbvZwuMpxcHq7UKfXsu6MNPyG71KomqjwYs4
YTzzw/c2HClGu1plKBecvGkGOGKcPQWLxL4L90lJoBu2tJ/iZPhC0to/T+//aWujNFK8pbiOHZCW
bwG3Pq4zLqRb8wIJ42kAj3prg9yoatiZZuSOv/aC+V+136gAnQbsOo7+oJ/IGpIxM1EMPPDgHEwO
n0RRlYFx25xW3OCca5ndrDeq3N7opF/MZXY3I7qqmb6HkszgpDO0lpSh3dfgH+ZFAdVm6ARWwTrR
vRE9pgRyIoGAttWXZrw1udlmpmFe7aXo3OpX89VW98YKWCogteAGctYifAuzMpyCZBknMRG3Imlm
Vv1IQlaOTGfSX+r82Ur7IimL7rGY2QXhiRlBG7yRuT5LA0W48MeshDse2XKDvGViNgdLYB698xy2
FMb+enLCH8D/h2bO9CstvNHY5pON+JwzOinVBHowvN1f78ZhcXpITCCKn8rIwOdaqHIiBWMNj0Yf
GEr/bsjTzBz7qIhetf9/58n+OWrejPNqpVvtAFr5gNnlGdibMVhkACMK2eLRgYmdJyMzwi7Rc+pN
XxVjIeJh4Wq7GPLix/IbGG0kgcR5ULLqhuouuUGDKIxCcwpTNT2nLfNG7K3MNF4CCBVkww97NaJw
0Tx7o0UVFktgIk24iUtsH6w4nlme+2ig3yIExDyW2zREr5gLQbO7bDMIA+U7IThcAPKlfr9ut3LS
TWKGDN8gzn4lsyITQmWptYXKEBEoY/hcSL4cHMUmT00mnEY32yfEezGznPxng/kKHrfVHCWzjL40
jOySm2ZZ2F6Rmwaa4OtT+HIjeDOosbxegHwnWiSxpJ9yCeklG7isuYslyIx38faRntDqGWPuAWkH
k2az7DDJTh+p9gjjNe5ejnrxuHw9jgxTlNDXFnpFx7WSRVk9PbhPF+C8ZMlJ3qybpY9gmhq08/P+
KpPHCZj1VnoPUYsdYd8HkZ+9qIYQLliIscc6x/AjnuN2X+f6EZ6Qur9p8NhTDvLuj88rYLM4ZBjo
cf+VQcgoJvsicCtv1dhRU/aNsyeRrep9+0miUy/CGwQ71WEHLSKZNWuREHIgRU9bkxAGkwFk2MKK
ZC/QvCeoNezUze08EIvPGH/OMGV1MC6a7SsHsmkNF6bmD4yjapvFfcAKt0qMDx3ZEDKM72TOOToy
h9SARVlvbK3Gw13ofEUrm3zkfwiLMpU5hRDQQV6B/vF+5NM90rb9Y4R4N0yC1oSJp+3b2ubcxLzm
LIpj+EMhfwJmZXc/JKUHC8q6eeaNjIFOh39A787gjsXeZ99KMDIS7T3NSe0NrxPm3AGBo6bG1v69
Tx5kU1XJVwZrd8X6KeqF8dzcc3PkKCGtgHl5VtuB9PpAufM5gd+lzPfYZ5GPximIZSsVu5tIQBoT
7NTik2rZ2DkwNlzH6VqN8Ju6vqQrLGMVOk2SeqElXzUrTMljMgWubwMfvsfFLr8Ktl5n9uZSLuFd
+6gk4meNfOFpg3J3lIAG9GCgggf2L+9B8aXNoc6/Z88IPLiLDsPOVleidhGKevOW8qffS3TJ8NiP
mg6H3eHGYAVZ2fx0azkQltIOPJq6+4SqteSj54kwch9qCVJ1I9GkIcKeByvFtI1Mxksdcw32Kp2T
mcLQo0MSus1xnuJNqdIny3rAmkQ/2E5LfYFFlnLr1zElRuC22WffhKa0mPNUPqMG8auvwyJ2XyX/
vmwzqoie9jZ+7WFFQIOiq0QZUk/A/+vC8QH63yO2qg7STeDklmIX4QmqHHcW4kWV4+WC2KiSohGR
ATuO7BGDnetv4WWKluEVAhF7D1AX9ysIu43LznrqtoxKth8OAFpVcm0/tzHZ2CLSDA9/POZ5TWHh
Z0ICVgj/fxjJifcTI2EkTwPoDybj4jXpbZ0ag1lFAQyCNA8BvBv0ukETsb8mKp+DPkUSLDbBum6B
YGBOiKzhIX1Q4sfZruTe2kMoOEc+OmqSB5lEN6P4begIrAk+2H2Hp7YbRkFmuk5/ZAylNGpu5uwy
KMBSXQHYjyCvwzHrbTsuwKMSP9GFV0N6G1ed/v/zeRQv8v+rIl/haucbn7bOjOyfr0og7NXltmtj
xSHFAMKm8Y3g8bLYpVMv67YUGQo7TjqhbyGe1Jhbf1icfDXE9I2G9sGxE73x4kHe2AI93GQjVnzU
ecwRdEkVlbsFlrr3vMPRLFE0Kr8MiyBOIBs92o9seS+VQdFG2M0zCu8OpKcdYnHWsb3R8RRkz5Wa
A5gBpGiy1kkgukUm5bwsE5n5UtCbm08oZ3gG/CPfE9NZpXmziixVPn3qgozQqgZF4Us8O209nOGH
/TpOhnaS25k3szyoxEDQHv18C4RL3jYXtLj3ewvhF+IUwKdfem8Oyfj187EPkY/eUxGclMdRnrm8
OWpWjSOJWisx5C9w92+jf6kthRHxrfMVzTUK17CMdEX39OU1gwgODRCL98AReA2VQCfvTkCGvWyG
Nb+n8f9Ek/oFX1rNKc18jrcQwtZLmyjj5DHj+DMpE6qNWtawovx2qDHAlxm/Qmo0rYKyW2NGv2ep
NZjYI/MsMFa0TOWcNSVe6wRnEOb8d39BQ+yuTTgJZiFchoSqvOgqNG7ovBrLUgLOotz6k5tpVjCe
W4Hk5rsXw7f/730GOxClZFnhVMADj9efHCY5JLXVpajjfm709Hb+96qXMBigao63ImAOSBFJZny6
K03Qf+TL0iZ+0WrSQ32eDZUH0TPejAEPlvBrmZR7F7mB31KEAyP/OKUIaHTpk5YN//ZsPn7O9FBE
Vw7td9wlqpGxGyDv8PJ86vXcV+0D88XACyfynVU77i5/SNkSfR0FEhXg8oL7Bdz7kQp/0I+EaOzw
ZUt5AB2iOWZskrz4VBuASobuWmzscJtn50GLG9lxllJ0LmT9Yt3XZqKJZWB+y800ZqKcmU5Ce7M9
dq8/MXxH1yRpt8jCmQRLxmHo5vfW7GusSYEFHAV9MkJEyW0xUqVl5mEUp5BPyfd5YO2yLh3aStQ5
/nV45nHG9yJrqc2rsyCSBExRDm3cRUkXG/UvoMQ1aTHTbVTMiUcDhmL7LWnCiMIrFzzyO6wQZBfd
CMiIroiNs7gfYxq2NixiD5eucVvUdfase2dXBjC1FGGsirfcAaWFMMcygOTkESQicBBLbEEQm7+r
zSYKtoMbzKqw9LaZtnTpcUSuiDvGO9A/4ioTXWs0W6yUUcVA8EYuyCfjon+XANFMfLpGhfKmWLSs
y87oTJlKKrMmnUHzFIAuNYp2YKfYKfmq8drukdl9HbwdOQ0YfShhtTy7292rfIyzsXfhCT+TYjdc
F/WE7/VPEph8Pcgh7MpLja6CWl03Sca64Iu/NmueiGI+X7PHhfXb4U+GxpDcyk1ZTtJKjYlF3rG3
NpOeUCAyGMXQNnTT0zkcqxIo+XRcmW7STnRawojWayVB9F9i4PQVmdg1lX7/xI978MiDfFCW8nWa
jNuEvB//XLunjekE1G1nDLjPoj219phnwbGhDATXRRoZ+pyn+Bb7Ty7oBXq1513RebdjXPCcEjgu
v3jogRhbJozrTA1nsCQHr1pLMXvuIId7NDeg28GCfXw9B/EwUdIdOszHCWADuLpMWSV2RRdVFFiF
bLUwwSWHaDOqJZ/2DJ1XT0UO92za/eoL8QzKzGapx+i+WLndO6hAAEiA7PK8VIDojtZprgggB9g6
OJdzsox6B6n8+nlSCVD9rYTRyy81HJ0G5X8yzLPL4ppJFSIx6swu8OP1dcDIkKbc6qIA9vRtNiEH
qhLY6DpY0WAKclaNcFwkEKWuZ4dzINUNCLsrY+ILlSm3VlrYRg9pFpVIl7MkptKprH/08I8wULWa
jbJeGNXVVQ+/OU0qjz+tsXWJlqAqQg98aleiQzr9YoO7hAjieibFSUdbi+WD1Ybekf7MZ1nDmuq8
8u5Mc+Mu2NrSjmA2hl83ifOORMzvoSOntlpEKaYXOc44Zy7u6SLkS931NyIUjbtL54vlNODh9oHl
bb9j5zpEeF1xOSPbIrG6SsDxi3AEobvKKmRHwYnoeChmgdw1TXxxkZPVvpf49/KJo7STgUmqLVdK
j9P5wciuPulhcvuJ6Spil1fvhko9AXrNQ5wg821zbEMENhzgBjP2dxAW3MCL4epSqxfDDmoBhVyg
APbvtn8xCIreY+R+EmFpBtWl1vRLlNbJ+OamIgzmhEqrDN7iuRT/U+GtySeR/VMu59REBQUxIeBv
3bmQbuefWg1vQsmwlSqzSHKorVbQYj8lKfR5DS1hsJOfMSDLNHPyv2SXK7ufLs3hpTBifoCiDYtE
8gDNvEBhwW3Ly9YqtB2FRU3O/gORg99aYO8Lv/Ybi1lklLoibtlilzx7oWUwda7oqPE0RcqGU4pw
MpZQP8Q5pBfjLWWyWre0LvljTNVAPeFqUPAkZhoxDv/WF+y5XOzbKdHyZWaCGfKCaz6lBALKVs2B
AHRGr4EprImXMyINlpkjyhRBrW8ZB2Lj0b36QHvM99YvfD15DoadYQ7jsqluqvXQ7PWeLpRv+ath
Y57daVZ+HkWSsUv8UQOI/NNy+gCUteZuhFRZoH4xj3aDqptHbnns8ReA9NtKaGppqUh2Gi0AFIwn
L9U2UpGZR2Etlh0Seo6JohSRVfLNTTV+yWzWbXat5UJ7cKpxMByJ7zkYdo80E4u0FKYtCnudWL07
LWMQS6IdlMBsH6lNxc8ssecV9EhQxMIaFYaHpECDplNCrxZ3UzoB1KyxtyhA3Ns4jbcozq9QR8SN
gCww87BAfZKzxpjPbMLoeRZmlzVR0sLUYYO6z1rmt2MQBTxR8m48RS8xCC/B0gUlRDq5+R5eqNAx
kOlqP89VtBeo8mOKlm+vf3EosCLJUnRhOmPmk/dhP1fFNzrE2+qTz0ZG+YFqe6WlwLDu8n+Uf+hL
x7bqVbxm+xFGBYwNKjDAAJKIU6v259V9K37HKzYWUUv+zpoz0AlUBcegwcvfi3Pd6Q8h1hs99y3T
XhhB7H5qzN8Jn4ecqssdqf0oDSyy3VDM24eBtoPvAAVQqi8lzpjDsLUBg3PP7V6XK51OpVI/uf+P
o8P75/7CIWJFzA9Q2HdHmfwoVFdQge5eE6QiNPZWKiOLyb9l8iY+gCWBpskJYvYIVMdFT6moE9CK
AefSsBc61AhaYOTAr3AqsYq0QRPKxOvnpT2npfeHgKuJCXhyHSOiS15R1PpekU9B3fEEFIK/B33p
TiOuYAfdHckX+fGt/c5wImRL3YodFsgX4cr4vCvDmbZM0d7HLAgcf0t0oUu21kgM23xgS3c5Qbyp
BvcS0aELfGIMHAu7v+h/qYmciN3LuMZ3wRP4j3ZJMXsbsozNPBC+0Tgq/JPzUgspmKu0SkGND5lz
SVCu7cvz79VDkuj989JRFo5ZwecaOskHqcF6dzJwJjUB72QaezaD5h7aSdkSYKDtmotb+8KSaVuw
2GP00MWkFVtokmjSaATzYpQmYmcHH6cJuRBoVXEK65T9f7OEqjcD/tVHeTLb4Rc4pdU+mLMjMlQI
Bx4chovCBWyufl65xW9jRAg8DntYzA0YIuc7MrEkmQCsYDMBtLhp8KcXqDeQRsYPyTuJQ2HkhSR+
rmo6k6vjk7llK5xMGjJb9uou6x+7J/0HWmLwN3C9lUc+ONunyte+wZlsynFy3HpDJfl7ot2XK80t
52VP0OMqcGH8+z779MVT9p/zMINJFnU3/qFr1QATjyAY6OUiutN+CtKFGucCKXgcWJ5+VNceC3aO
3OdBHsKh3m0VXhAF740XN9e9hplx5uvUXKPmVfvuRwN8E8pJ8SS7IhLgz7KbCDhE2mLIn2aPFVa4
BvJA26xLgN1H8DCkcjj+VkdKTsaMkgrtvuQY/0iQSjEwJLVKqkdBQQcretaRXD7aRfBZu5X0MUxS
xofn1MlTuXqTXmkYSVxsPr385NZM26fA7pgatWoxdhRaQLYZxwAYAoxxm2//7ebhRPnAmwrzS1Mn
xJattaSJgimEFN3s85jtiZJgY7R1IyWicNB13I95dYH3lBSd39cmwId9Isww8p6aV76pKW/Z1ymB
2qpeOD93Av8wmB0EPO/kq8rA7/neLYgeh6DB3sZO9veQY2kwxa/sC7qWu7sh1g0U84dSQuv0a+vs
VT9OVUYMmj4gx+7CCyWnoDo+MU8wfGazh9aBaWR5uhKgdNGbvOcmloab47F7awfhEFp/GCosz6ht
2TyjI5UOkqiSlh+lX8eaTFOHkh1ml0UsLkBWwXMzlCcX2qeGAZzq2LLX6fhA9irKRtGmb1jZ46AX
YpqvXEat5WWzATo0fs7s58xHy3gkyqm3lA9V8vcqR5L1IJOiQUUmMUj0n6MdiCfhV+GRdtB8t9SX
jFEWlQcig9oAKEQpYRH/tHWfIcZOEkbIFOBbaVS/pg59l6YXcuimOXI4eUCT59O3vZU/i985Yk/M
n5ohr828EOpVhwVkt2lyEvXdLNDsGrH7rkMqdf7gCcCmCKpoBRtTQxy/0xg7Mnv6IqvPSisCJGm7
OhQkiM1ZoNWb0Th534zpa6l1pjkDKrldtXTqiO6So5Eme7c8QEi73QvnJ8QxfI27thQywFkdiPMX
Lq64MUMJ95DGxjC6Kb8OgFqNUJnyhcpIvrrKJ6p9qaxsXfSoP+pGDmwwcO7M8blwq1fIbWtsJb6L
2pRyaeMY06w/Uxhr8jpxqToUKwPWcRU9i6RUHHDXqVK6FFk1DOKnzp21Ju8MeCpd7NYNLmse+MAL
zxLNkEsOV5WV/8fUCMpiziwT59OvVEc4L1kwBY/if1NKVd2zRltwlrpS0WRb67hULVkZQ4IB7RoE
2DEan4Wu+fmf0OZ+x3+azv8mxUn264MBMAE27Q2dmd5z9ktAwilepn+SwiMsmuUMaJgBmeAwIu4u
mGdHhnmiiI4urBcOM9Ig32v6yE6lzVi6i+pirLdRXrDeJxIyQgYHc1mt+uN1iM95QNX4mJc7wKdj
AboyGLVsYjprW5/Vex4ZJEri22qmstQJ9x2hDKWCE9ZzWpGipQfBIiOdOM9wPQ9AVAC0vLzFUAgn
eLtG4xWbZTF75g4h3FDgXYr9fSo1b6ugh++oMDYek374dUblcryMkVTc1x+Br4jY04lY7rx3Qra1
IexkhjiWlzFBaxqCpH12mFSgYqicf5h88nHja4+djzCcmkaepGQ/nmwmTUeNY6grSBmatwldhXZG
LnJWGDk6jsy6aEqu0z6rUsKoLEa4N2Yaa3PCmWvmunGFZwLBuLFQj9iGyifBlhu+C+CcCXr92dGC
P7o48PTLUiqy8Gtyh4c53BEix9UQxfGm27qlH90XUhqV0mpkorrg4pFJRdFjbBRlWk8uuwqtmlwm
pkODQpVJjRKu+m6VpTLj8ouJzRVSYBxXVRnTImESYJKPgNMlJeIrX4KirhBCv2AB6KJ7I46WrIGD
Cj2xVqcCTRGvJAOIzvJkpCOSFczhXcuOa4GHzu8CqhKi5foiF259v1pKPHbyCHesm3slkNQQ4tTL
OMLVbc54wc2pzN9e+2uVnmkMIdK5eQHAa65puYkqU7AKxkZzcUOp92DBj7+1pvaHnJEf7ilfrkRy
Xq/62A045cKzDgrR8NsLmAuY68756O3ft8EDXsj0d04oYBjgkrhF5GmXo0pa00kBCvoQhGgyn9Wc
Uz7R1ht3Q+OCmE02+ZgwpyIybxd9L4X1f+8bIes4IvKXCRjYIZQUc2PkitVhd1yvVrgU1xnVEUez
d/4rzWmx6x+XwNjHcsxBovN/bVFvF3tOqGQgNxmH3fjJsvr09WlphGVe8lNFtj3sUu9ztFtKlDLl
yc+sHbtr0g+KEqFmvffgrAR8s1jOyiqAdecHWHcOEW6Wt/9uO1FpfOJpzw31xZevaRq6n6Tg8WJA
kr+JYCJ8APHcdjd7nvPmUh0VzMW4aTIicq2ufPKCe7IrHr2jhspw+H6RwHWIONebwxEvROdST859
zKRtV+xGKywhzsDtujRoSw7iAoVKDRyzksJalIrphvRzagPG5vl1+LCuFXdZGDG1dEQf671dfo5k
F7VdRRXUPc7lDKaWyxW4KJ0WabjjVTbnNpV78/3AHhrv1QbNoSxvFVq5dnx5d83YF2058bIkom4d
a9EpPsub4ADSES9Rfaff/0UEIPdhCLYMHZ0So0Y3sM+JvtTINiIXjoCP/cS9aKtyKv7k5R65NKV0
9mLsqwsJ1gjg92e65iGOYQAhVxq5xnv6DK/ZcaubLALd4/lLTMpXVY9q7xdw0QrsCqT1qy7FIAj/
AYqfpiKwYnengT2O+/FsARJxXdowP6rjTLS9kRmWGDAPSVky/uHQTR7H2RNJ+ihtM9sA08obYcTg
FNZrJZ+wbFCwmvXuYgFiyhvcQIanyGcHSDhTxFrEi4j69ZlqxGbBKDYqIOwrU/eKwDxk3icCoVN8
qbFD6aOYygK/LJtnZeZCKMyVop9FG+eHc1YCs+GpQKRbw/kyiA3yRYhISXRei90obJhdT6cWY2hs
nvCiR76RDZZTjr8t/Md2/aNM5xWrbTee/9ceiL6Tro0KAJx28IulsWWp1g1by6DPF/4umtLK9JSX
n8g9vPnZrcxFbaDbQCAch/31EgzFahbMSK14JfTZmn59YcaTa3vp0dqBCot53VFzXs48djyHYJsG
+0Zg5WXtV3hHSZTIInKIJW0IIddK+clWhbQs7ZEXb/xCqcvBg+Rf4oS+ccLMCajR8LtM5d7QHE20
gp7/MKrtZsOK9B9ZyYwS5QCqDxzMmC+yGu2brDxOZFq+bjFzC5jwQ8mFtdi2otV0Su1YFBz5PWli
a7e1L6+hzpAgfiGTAjS9kT36p2pKVuM4MHyT2HSRDIXcddzd0q8PNeZKGNYEe41nldNEgJIkMYwN
pRRw+r7c1L/yTXwv+izkyLWgqAx5DsQd/AgjZy7MLrLjerjSPxwJud6z9+J0lLIyhpcSkd5XW/MI
Y3bwKzKvT6ujPZq/zbLeYjIBwJrD9I8E30iNs5SsWL9/dDFu1zLKc+SG3Y9/KbbQ9Kdpj2CZ4doY
SijX87Yz8InEMnIFAYdFe7XdD+Uh8XUKojdBcCErtsOYD+tINhCmpVyP/s1zRufxsvN0fSP1mehl
c7F1YL8sotYoDL3iZHTth3ddcuRSPGWXvCWgshPG7sWRuRI4OHusT1PdO1XygYjI+TD4NWkpus1x
xdJg5q8aTrJ7WQkQ5/1UKh6e6TIZX5zW7s/3yPyMej9hIuXqPAiv+CSbRSgVoQmiOO9cGN9/5CIN
tI+Ar6qhSXFG1mbId+F0sxbX08R/jPx/GKfP3Fu6LfKlJz+nb0f9Fr/eN9X1N++rZBwo430zhWP5
jxDtsMPM6UcmLGt4GCBSy3a+q1NS/UC0h4xmm6yh8aeU02NXQ8e6Fym4gN/vMUoWMj4+hgPEKHFo
D2PmyzaNtK5VAkj0BbGxtaiSf3ib8HjnFnmfGsh/3L/S9z5ew64gor3PKJWc7+43+GMvcScyCOHW
udWoyw+nPtzq8pm8LMTKPmGlZWWS7Szu6tXqvay2IBFHdi4JQCK1i1/1U7CXADUBCS6APkwKh4jK
h8PONjED/bal5t0Q6XSuotLYCIeQ9rDekEOfCbQGbU59K8Ua56xQiAE/0cj4EUDJBhb72m3aW5Ax
9hao162QJsYjmkyZf6aXdsKyVJD/EvpmiDTg3oQgGCA9dSCazvhOiRL5bZSzajqUMYoIf5CNUtZN
Kkq+hAKuDMraBeY37sDBSBA2P5doo8R1i8tVpqDoVIqgjfy2TI+IMo4vBnn7s86bfoBF4cXb4PGd
Gmz6e7qTqyBjANj5Wds6LF/ic3kJufrjfH92kjHuJD/FbgbnhYvs38AwUN+8fOhw0MVi0c9hKQKc
2M2Mf/hyqBwCulvbdNu7WQDCkDgCNV+1ndEpjGYsiBNFKzzMKLmOiWsYP9lJI4UDyghSaipzG7W7
qDsBpE53yrPvJHIC/x9UynIrqFDjvSBqIGodDYAdOyuhhRFTk4Ngvgo/A37Vo45HYbz+4YOK8C1u
L51PrVh2z7M1wrkxPtzuAtjrxM4S1fN4OiZQY1lngUCXstivCw0qK+Ch586UqFa0pA8Ixhf+CFCo
LrHNjQffTsaHxcPEVZVdQZkaH4IJHO5bpsWeNbK4UYvqgEWeLTqPywHsixH67J2o02TLmIWUFjiv
y0RvkAZP5ghjXPOD3+bYOIPSYCevh2M3c8sml53dg2SGFhHX1VK2E+6mkFnFh+BUg2cg0Xi14MrC
RkWtbixFoN5SHOqYYqaBwtIo6WeO8TICOpTlMcGYWFE/PIe4F4+3zchfg/mQShPj0aHLlxyFEwjT
hTw8z053QNEVQ4/OoKHFQpaPmEBfEHqBZqZnUL7V155n5iRG87psiSQzavDLUXLzYFWiaCzb1pry
evbkvLT2m2O7YIZDiyYvL16Pn2HUPizEFaRu9wZPMecPkmGu3nCEcLWru49kqyVLL3c8opOnsfH4
DBQKMZc4IBr7Dq5PFr7M+Kw94KsJVKTVHXE+QP6ipqr9cmZ1Xomb8eAH/1uHjVASkCaL2jICabmU
/t7ubdzgUPdNg8YF72VUv6wkFLkIp5CgILiRXZf717nNZ31ZVfNeUrU41bSLMsrcV58/wzQc/IOC
bt5lwuLa43C/sFYaaliQmvQgO8mWXKGPS/SH4p329bq/oauyRfUjOee26Vh32rrl9keqqMNwCcST
mu1BCOEoRRJdZYZpHEi/qV3Y9TNAvYWRy8oBQfmm37xQwoeZdBfnzp7AMRLUN7GJiiIaYv1Z70b+
7WeNDbTUSSlSagXWsW2Se6ulCHmEoKWhCFPlFm6gZ+SIRU3xrUkOxcQrGOF52vU5DbjdzDKTW47x
6JOT5Q8Jdzv1Iv7jL0S+YHxLY8VdnARhuMMfl3HzxZwMeh9m87NPV6387TukyDd67icvLRplwmYl
xs2AV/GiiNPL+XNiSTLJ+/009iW4TD21ZgsQeejLMqbb/hq4GEYaI00wT7oTiMLVNjA+ONsJ4aO9
G16oh/n7U0LUTeSWrEpcw+qPwH1VfNC1rCDBS46KchIJTstKMMDq1QKGyAFuC9jzQWGtYAm/Zoip
S292VZ2udHnub6BQXZkN4QzE2g6C4KB8xJlmc1bsvS11DBvY+uPTpjA10fi+wc1clGB5m0RBjvu8
fVrE+Pczy4CXiZ+cX1IB25dTGXHjE2kWZV4Gs7ZsN5VepFn79MH1KsonQrzQ847ap0CA9oJ3XViA
IJRx0dyuipowY4uXUMx4MfjKNmMeSvV/pzqxBc9a63a72nP2IEzRTuE5kv1fdCR2Mrq+y4R0Rk1H
tX0sqkAo6YCvzYPhgRQpVGUVW7U4uOGmYw7u/fPZtuBiplUTVR7AdPGcrDbqoUD+Rb5tmvTFykMS
1u5gTkigvA6UWmFt00qaqEVpzq/AWIadiRtxJU1ia0guuTtergu50RVREQxPiCIb/84JBcL5hwih
AkzGvM1aaCTjoyAcIi6FeSQi3bXeYr6S+d1HK1FLpM7DOBenNDAEVP1ipGUEBKnplq0mArJnK5Ia
8bcFFRmXzccCE1qWfG+0mEml7D22pLT5VEAinGv8XUANxuTyClyzucJ4o4fxsFLPYK43a6XCRZP/
jmOpMqursNORnsDhBHtMnBWB50fBEoM0sZ8bbAV6/uj1/W7U0xBkj4A3XEI0W90je8TGTyf4G3Wm
hnGUBDXAd/+FHzEZA8nPCGTdGj8Acvh20zFCNOGkx9XLjc/6rDK6fKvKcosxrta0Yob1qQeDzDFy
PcnxuYYP2c/ej4+YL99dxHS/vRwtGn9t2ra4eygTy9kwReWxKvHNdzHyFU4o6oYzfB8lYqEg5ufO
jbRe0dWb+e4Pohrg6Jw7J4B7c86CdbYBLtoj3fuakvsvEZ78dE6orFFuJmi/Xelm77xTvLoztBGA
lBXP2R0UJraB0NrKH+waa1wdf2ZPE9og88z4J8JL6p7bwzLlxXaokIvqIWDKc6MyZ7WhoGY6Q7a7
sNMoOvoYGSo/ZPKXzYQjdnBqrO9YvJDKiSHZyzyxMI2heX53REaEO/gQrZFNahZbZpeYP0R1L4Sm
Akjt/yrX25a3v1xRV2Y4jcYb//VCJFiIq+MYNMTW2qRlY9LvlkjHIrJgRxEKyvntYekxpEDfy0vV
EmxWVq6CJRiVte3nobPxep3Mg7LuVhM2IYHU9GNRjVyKgrlABHNByCRZElfZbHTUFMNXq0+4F5qH
KtgrhiDdyqVYuUEXB85aSGqz9fjtJp0jF+th5YrHTMvMgtIUPiaVe0WCDzgCyX9VGIJKsaGjhaQ6
HMGDx4DXisHJGWLWl1Qdy7/cNH2tpkapo9eCoAEoBR+VWaTInO6ggP7GefYHVNZGELkMbTIlXg4p
zQ6bpbIFx3wVfsGFeueCqmR6TBqxs8JpLEqrAmDbfK7Te/oV2TA/ZWozh1zx/durpOEbVzhIAwCq
Kos4SZ8CNpJC6T9Zwfr5h5EQo0pN1BwJy2HymWzcnuH9NpeoLm8ElT8M/EB7fBhWt+tHGyUOK30F
MedFKFGmQsNWbWqFZB9exeSvnxojyGXT+S53Jeer0S6g8QSkTfO4kPunXI1Ot5d9Oe4dgLAMqy4O
CrQAav0lc+I6G/3rKFMorfvrq+kcLeS4lJH9dfGymARM75XWu3lp7KTyquryRWNLrnmaTJD+vWLF
uj8nyFYs+bnFqQwP1cqypFwgONyGPjVKhVuTdGnuvqOnGRDydgOP25XeaGlIeWAvdf9RLaJ+PQTo
b5tDJGmrjPQokjkK6tZy2WJj7l7sd8dLECpfpp/QZnIPcmSTL6hYDeuDkT94iSQBVwgnVkm9Xsny
1lyB8Oy2ZVqUG7XdO+ZwYk7Pd5JpUP2T1W7dHM1yngcpToiUYdj1+RzRPo626k73nvHphXfRCZDo
9PlwSxusxuTuO4ertW8UPtTvMTUliBkN09y6CXDhqIO2fJo5VR/BroxJdozZ4k5XFdmCyYLoZ6CX
QPWBaUUmEnM46N/2nnneadEnYbf6KQ+fVCUeX5WMk5XucBdfnb/deLMBOMRhnLCegunSSGHQHQd9
IrBXEc2Ll52oB3tmMxd6qAsriheUddB4OfM342Z2CUfZWu3nY2GUvooSYp2BWaEKJr+8LiMD3pgr
F1enxNb8P7b6HBlAjOu2EhN9WIi7448yqZGhytjlH4i5WPfgdVfpr94y1wZZw6kHd7RQzhsgln0x
MXmalSxf0Q+P9uKJEEe4qw5XTTSdd4vLNCs9iy5iefcmKI5Bw12ie16CtEFZtx4aQBg08Xmo6dh/
wyGaaVNyr+jOJ09IqQgpQ+bzjpfV+IRZ+RPn2VdmuuBeaNFwjMuxt9SdN9kehf2IAWE+JU3/awIG
1UrGqgowS0lAg1IsMdZqz/YkDIr5i7PlT8vgke+BDKZxqczr2hVyXUPqvLF/2cqHuWL0j092o+27
78yyTvaaRFIpUpW+z0YSuNarXkiJJUdur9fSqjVZkVrOw33H8pyPJeMLISCbEyvjuX/YAOZNKjiF
RnCBT9vfIAMPP3FXnChCLSxT/CNMEmIL7XDLMpvk3UOITRSc5Ri9e22SHibXaqQ+37pV4A5j4bCM
0TdBdhwpx/vGrPjFuwP1bmLVofclrRlGymXiBqQgvLHwQKll1+aGpMGLZUcpAYD8p3VPkV+6dnAw
clFG9JatHufbiFHQFwPOUNNp1yAP5rwvWmJOcLmhNpg5TMqyqmV6U9W0Vm16Vw2b41zqn3/ySN7f
o9IF/w0pBGjVcGhYt2FNElIemqLU8KYD0ASXPMrcho0P1e/0lYhjamGvvg2EdNHoYRzJXeJTnMqU
/XtObRrz745oTBlijw3Ub1D5U8BhAKLQtrnkWuNZcw6CaL6an/LJbtx9RhpPbTKHDvw+20rbFLTj
X+URRjHC+evgqEP6owEecbqEBEsUNjFxk7cs/kVGlHVJVHeT74yo4eY0gMeHvejGIov9ETWMzFFd
DbkYoFZpK+HlhnX1atNJ0yAhetwb6l/rwP7frek8dev4xGXfIBaCiOz+ISqepd3LfqxXpqrklND6
ta+W9wqGFE6SreHpK6d1QBXdhN/5cGf7Aq6IzO3lFC0Zzn/Q4S3Z+zDF/BfgHeSFDukLitjExMlX
NmYD/1r/95V4GsLxcXIOBkI56YMo85sSZVoPUuk57sRMT60KQOB+WPF/RH7XYg4PNX2iUCGPaO7L
BcHmPWtfBSEN/0PfN8npTtle3bPkWYg7uVRuG7dhkFYiVa+vb1y8Ncskrf50xrjhgQjXaM2KxJxu
m7pxmaSC6/YDVJsgfYv6Fj3whXt4ObXxCn4Uhjiw3CF0tHYGpW+Hqf3hPzUSlHQBXDITveVhK+xn
rG4z8FSlNqwR0LkjmuMdkqB1PXUHCeK5uUhfkZItl+QKtlp3vnXadCEXE5enjf5u3SurYDdoDAiq
/HLtKtaw3xNqC/paZOQ1FraWx2TfFTrzVKCaWZ119vIOfKkEX1VjHaFToy5cAJmiZwe629NqsUiU
/ievLF5xSHBU2JK92LUG8JlzI94EU3f7iaPCyhWF/2A8si+TT7snYczccdQyCad/7NJL5Wrrq1MZ
DJQHgTd/dD5DsZth3inG7ExTLWWso2N0q9HyDPPpATCsietEGAuOTbVo9wfyc2BzJdpGFtM+B4Pc
jdNuf1jjqqg2SZFG77kL2eyT2dBgCq4DDrxRPrJNE1I4FMOb9oQTiNvHTSYFFwpN/rzBwJKbBP1o
2ZiMp81ChwUl8zhbA7rU0hYbI+vXFDNlWGOCkVxe0A==
`protect end_protected

