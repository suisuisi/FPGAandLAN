

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
E7QXSezI1NKn4wecPKH46GEmlb9nzvPiNp7CjsIFK1lm5z3RANjb+gmecESP+TBysVTwNfFAOL/F
GlaoULdnzQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFi6SgH1w8rzW4G0fLyqSZ/w8OjthdyWl2P/Vqe5owouQGMrAQlf0HrqTY+eyO7EEwX9Yn3DDYU7
i4QvZSwPA9LCeonGNR46x5ZKQrjDz0E35ywfbiPVHRcaI37RevHgVkmFtj874p/Z4N7cGE53kNrn
Uq5J89OdwlOS0crhmwc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DElUvLFa3440XL2bUo4X3CxiAO80cMFl9D8VF2yZYdWv3cLqHTJKRxY49qt+puj85kIfJDxdD5ds
8WCXArH5YrLxmzo+h2GnWpE3Ion7tGeTxYtSbCgvEXBNR9pWuJQHezi0HocBG+vaxAxmLT5GGMcu
kEV/Ga+Y/eu2nT55xsZX52GPHKFaJioWh6RR2A9yC+cmFG7+eV/hCIeO3SlIwBN7lPMshiU5W6A9
hIVzXdklOZ3MMBowKWV+LHGytD2N9Cl7MqqLJhK7/d+fv+Py3kXFQ2zvHNlJCQKbOygyK7rkzN3N
dBTOVuG/5cAR4IjhD3Ez1LNajVBqeRb1bCSnJw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PoEHf8jQc3577GH22wzzbN+Xc3+r+Je5kxpzq46YSDf4RwwtJEgu4oig+8mMg8cvS5XmHcDx/ZFc
A0d7/DV6Rsg1ANL0Kc+354PCjmGpxWkLAfH+CL/KcJk/1poL2B9UHd2YUZSwt7xioiNx8mkEuKGa
/EhmwQCzP4RofRSsnS+N3xRV2gDlyk524IQ+QhS6xzZr2+fVEUruERDccjtpWc3727b8JewCFbc+
MmOhYgmllNMRGI4gTFGoekcazBFrCnzkTrfMUsK7JzDe2e8JTwqKSGIb9TdFRCNC4W/lkfYzGg8j
L1EuKWaW5XLg1PLWRKqaDcxOsZ2Sp6BvutX11w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GYzDwwwVcqfFKbqcfTh76yYTpnTlgyHZmMVVbWjdwNl/gdjQJPJ8FtsvWtygRGzbFYNbuA/99502
digUgEPD7rFgn689/c82BnwX5wi5SgoAHzj2jzT0hssD1Un4my7/N+GlbGcqywNZSWKuLhMF1a3h
bzU/CjgyYGo3l1Ki1kprlC5jx8W5BJ60j/uNzuWucV4QrjbQGo8Kr8fhKoXFAHbP26k7trFY2JcA
CwGRxffys/ORgfdBnfr1w732ppnL6Yu6Pe7Knzh3zjPD2ix7cCl+FCxoRx+r0KOCZqjA/UTlKWfY
yY3BcNP3hDgRf5582rhEYC6XWhLhsrRBSqpOdg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fEWbX7aE3ItbJhwVvBUCIwm9nwx6jL3zmqRq+s8oLCrNCK2LKFN5dbE1J6JKmSOVD++dlIuQAJV8
H9x+gnCuNUvzQlcf5gajwIOp33o408+11FeqlxyruPc5K7miSNeV032ZbrBFFI0nGztx7zq/ZRzC
+Tq08f5/EDY0w3yZfD0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ikx71sNg+C6Ox74De6LKxBeQ30HMlyfx3FZKWD0wAe40ISpT7JYa49Iq9hzmDNiFBRKXmSj2gIB2
qFWVDUvIfXDhaJj74D632hkE9W+/ZisjbVnF1EOoj6CglQ80VdSZ2M8Q7exM6+w1nsgrPvPs6Bk3
+vZlNoA3WRvNYBFfLeTyWWYRAN4yYUz2qDmbo2axCgXVKw2M6xfn6e6ZtYEDNL7sz6Fa1Kq0gm6/
d6tFg5cf+uEQmdOh80vV+JEncLUqh3LPiVM0GmegJbdXhocMkmdba5Kw3KAiHkv8ZK7Co/O5/oSR
m8I3YdO+yaDQAVEJxBDc+WxzNcJru14pkZo66A==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KjiRPZxY7uDBtsGJw0BgB/wMRzca+O1rKZb7HDvQVX63615VrREbZVFjO7wXnHf6xOiids+u4//V
IcO/1vmqVqSCUQCQGHrfhGTS3sVVOVoFEZ92Y7aaGyXKdF/YkjossPTj+stpEqyLvk4+FbtKsaEm
EKXMQWryhdvz9a9Gto1k76ov0teHt7YrGmepjNLcWQREPx8hli3B7BleiN4baXIM8HneQu0tdBBg
cST3XvGNsCjRQ8Miz1iCv/wMO7PJ3dQvf3bL4d+hrz6s5mKXZoO4pSUyN0ws9dgzQvxWWkhkQdro
9VIzJy19U/YUEaDfRZoh3YFgy0K5tMtAUAOPtQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
jxcE2/MjmjxLrNiuaTPmjpDITg2c6qtJO0UQX+eIMZcuX5+uElisr/qcsOtJ1Xd46lwA4zt8AMxp
mEck1vvNyc2GAMzCl0cqIgF+AD2/FBU4mi7gTpSoSQTH1WJQt5HC0YI2aybSl5auVu+H4Qvutihf
aqqKVb3e69BfjnYj1pudGX12Si7IxpQgRCHfVZfLo9AbUb3STGrYTkVAjeNO3pYqas/dmEJkRrY5
wsRqyU+hv3n2i51CYaDtzjFsI/A2gprhamFd4fSotHLwBXyBhNKKg2Rw1jPO9HGX43sh4CZX/5vN
NgF62BcFudzgHg9RQ15KJnV5NgTyst66YkbiKNUu2e/QECX+JfcwITJkyZEJoxhbteySZ5ZtlDnz
K/uSnxkfk99uwT4a+iajKkYmcJuKPRWOYuda/tq9DejvApbgqXz9DpnFalloAX5zqlN7pM/ggQa0
d4o38FFt7fvVl9bLBMBx8M/dG6tdAgSAw8L0mE0pEuzXhpESSJCsij+7cLe77f04pJASEBYQ66vn
C6FlXyyDteFwjZ2+XkcI6hZEkziisqF6RimxVn8LUkTSWOB8AU/4jWsLyActeCxEJit0+WxZIHVr
XHNpHZyO6vsf44bE99fPrC/4aoD33QpbVeknO+OvwbTe+ySlskWk1EWo0cFfcQsYSVWwybqiOjzd
5cZ+CSGN6ZywgTZ6XO0sE8mR5Sp2yEbLTFAYUpeieIlCoSykmsNrIqfeN8O8Ws5561brMOmL8E/6
KEQRP875PnmE6oKg0bkinU9iYZb57b7DIYJWVXZNoq0QkEJHcpw5v2eYEFMAN8JbCl/iVmMdBEKY
PtP5kYa4a1DyN4EWf4tOOxOZGsB96+X1hZ/duPY0FGf2ZZ/+teGAEoK4bFRdeDyD2Ykreo98i9Ix
2a77Iiyj25xz6lhVbQ6yqGgIwWLJ1a2vHKtIHY2VswJC35BpgA0834XPVdDkDJNHt6zm7w36IhVQ
/j4IgeWXk+Kq5wiiyjRZUzJzRfJZ41K/SFdxEAlgeiUyWeOK1NJ+vP0XmUqylByyUGDGXRHSYWm5
jPib3Y2YJ981fqEAi21NYcOLFVorJBWxb9gmiB3gQeIUGgGyMWAT9DpoMQ1c3ZekTDHsHoYfvkHF
j33BLpQHgd+uqT91h7wFNAZmQT88qAW9LnheI+eHi9PCu8tYEkvDFd05jbCqfhURVDOxC0bSiL78
XJdCUeAHoHH9htReTliGiXtl3GCnipptakZYf3wcKFsGVYPpQKOoDAXnvSCj6NNjxaJE5WMazYnD
OkkB9/WOrKwnFuu/F6TXRzmB7jWQJaq6lY+G3Frfb9CB9uLVJZQTg+XbL90wfB7KYJzj/HD5cj3U
0R+dasoPN7Oy3W11e0zANPRHmp00KR9SbAC874HPeHedRjDLiUpD2uGBiywVwpoISgnLqiMA8Rte
LgZ47hywsOorZmPMI1OX/LF5WCaD/o1GNoENBMZm+aW/+FJ+Bn+iIr8eWHH/9US4MzzK/29C+vMI
D+rt9ZechYHI5LP9y+IO5ivq7JmbIBaqPvRglPa3ouZ7rBIpIBbDu0rIv/bbixwoHCYWbJ/mBJAn
RgJvENlWPQI+snzj2AlRTMUn3malX1IUo1RkRhuqkiM22MtWCKIwO57ZBr85TJAqB70TrSxmXjkm
zsQ4EmyFitJrdoIKFYfnDrQjXRPFDJjoCA1XIkGq8QsFqBR9Letjicz/iYzB4GyVUNjjDUyg7ufn
GruJAGstWykP884aWS/emvLVWYmwSnCkHLWDQ+xTBFxplPH/2IVPMss0CMl45IBWWgtNZ6VBuccO
I+dIkMuHtkmiU91OdH5Ymz0s1AqYBD5QJQMsyDbRsezrek2xdIT+SCq2jinGwtKqY7Qo8hg9z5jN
J2Ysoy+LAoGjCpkB9Rg7mqlEh44TlkVW6OrsnDpcwOt1JORmEtYZCjAnPr/hewkdLVCavoKYtYbD
2Zdhy99CBtjva4j8lcSDA5YlkgnrF4VRjaidNV+0wSB/pm9tFH0dP8TZYoXLK3ueTZI1VQCL7gk0
RI1kWFsnXnSwFsvVdZ3Y1YfJ619WMeFm8CM7QA0rartw5fUuDPtQ7XXVTVZXvtV9fEiR4i/D3YvH
FZv39AGslIs9gTR8mqMDBg0H/3sbLCBXQEkZ+JV8A/n9ZvrmOE58YW5qkQxgCt24ArdmXZVAMge0
XnaA/sNVYJlA7EDNkgPBLo91pr3xxpCOVC3+GjJFmbSJEgGS6RGADR4Q67jxFH7S1OCGxfcyAx6s
W1h7IttxidYhjMfSkWLxKQjTDD+8W1KsPOsgQA8aMorWyYK98AVaB2Nly5nzKRPr+ofnuvFq9/0L
xP/GrDzD1CaIIV4qgvfySCcpRp38xQkI1WqvYAplaE2aopEvmlzhDvCuShW1GY5itSiTSMwmGiM/
84okf5AkepBslMPTy0vPH56r62YtsYLXGRXIi3ggMXK3rYfhY5y6WEFplAckJFrTrT2BZsoyMos1
YrSRkiFe31b/RONCQVwDe6A+tbnIlxCfRhBbNwULsVChAtNgqZ05HKiN9/LzvL9uspAhRmltAN44
M8CPBnLdk/YqWnMmTHN6iLK2FZD8KBh5pbSrWhU9ECpY7ii+mmtzVkUVcY6Vx8t2PfAWJirtxt0W
24t8Gv8IJvDurNW/hIDt9dM/IcYh1Ledh8P7xfmDPCGEm+PN9T8JhvgAAmb6w494yk3nbjxCLiSK
67Nw2Rwat05aZV4dQivecKdV1lo2p9N3wazwkcFSG/bheGxVSJLVmtr9QlLPmkUU4dbwcdNwm3Zz
MCobBiJE6udKD607mztHI1rNnXJRlnh5Hty4mXvU2Um3kZ9EUNtcEm5kSMe0kncwezdJdgDdrMkD
955LqGGt6uIPQUgR/Nu5/Rxc94CRhlENzomGRAnMrvqrK0DCvsxo07qJViCmLk54xDFTen0q+c1T
mGMDDBGVqztYw95SfHRw8y0QUqhQP3ogWL0Hy7GjWtbtBpRdn29GQDdQmVEC8Jy244IMnAbGsw1+
j+3mvpOKWgc7zmaIV+pHA0gTnji3fZwO1PCQp7ndgJ98Mjv06Wnw5Uirb4dOl3I8DrIgFufIM9Cy
LSpQAyx2wgv7aEKUT/GClsZC1PpqdJlRqF/s4Tkz8iI3ZLhaqQ4UpTFIu8drdWiyr/NFT2RGW35e
R3HLbk8NNuarxZXgQEqXKFFDrFPTggmMx+WxCaOfaBLSDPpSoL24/E+SshFqcPxtuTubUU8XYXR8
8R3cP24yxTh16Boyr1PQAd6M3Bh1xcFyFgTYZ7CXkTU8GKs4rw12qdWMFlPoogDvrzbsd6R5k5Ib
fO8eljjloUBPa2T1OLFZ4fbWb1bVlQsET9Gx9lGTWcOiXEjVdksGnJHuRw5dbRAydYtFJIAYmq0G
m6r6zjhUXV0O1/HPfNvjvVO2c3nYyB5t5p693vC/uJjcoZUHiT3jVyALD6RRLgWZGy2rAAE+/lJ5
a7wQqQOiswOmduV0QNpThrwQR+e4unZ9ToZpgWJkmeuTHjcT9PXfK0c9sKCCPqATJ/LuejI3Nd7o
FhTCCZkcjfd4HR+SOtSzCbEZ002tH71TasgwvYdE86X3IwR1qm44pRZBLRW+8crjHmQ4sUm0QDyh
5sdV5z4yoyhI2bmniq2TfkKzQo56GdMdQEDuLmGHqiRli07beunIt2rI45LIzryDg/14MSamHZKi
dx5UzwHVaXjfSmMUWUnROHwJU8/pXxsoZN2BKDtE/1JlvQyrFSUSnFrZmDYFXH+Zk210be6SZ1+7
2eQZR43z5Jdc0qbBfXTsFWGAvrBeCqc2R/7RqoxyvJhPMbILJA+vkzuGNqWPcQhwvIDXH1NVvB8S
M1/1A7yQLRIfD5rvacfCeewP1afoaqrQNJ+uSeqQS1u97BagKv5nqFKl+yWQ6F1Sp/JPzg4EDYRd
M/dP2UClrmE+Jdjyw5NNg08dd/G4QbKH7vuCA4Sh8qOnkXIbLTQH41ROtUBUr+oNDa2qnLZ/jBVA
kiLv7pj9myLOjuNPDes9TTrxdhZJtLSaSGB9R7FdoZgXAZ8/uXpzb7II1MQfWCw9RFBaVJ17z3hc
vea7HIaya6CZaTOKc6vK2PFtQAPjF/SEYaQSxcHNVY3nTmyfSd3m6WM3iEDIiC6cVMyeW2lTjmdE
u+p5O4BZcYbNHu7N2UD6Yc5RNHEb6lT5Oc428GDCCdkAz0uOFlY3ldXiVJBUDeDYVaWbeHQXmAOZ
vcIhEUvMGmsSGhxOa+HYTD9e90A4LFjiswC/beI9EEPQx4xmDYyqzsffRSR835Dbu6HFSh/vGtVA
+CwcNRiC1ZhRZGI8NybM93Dwrhq9YosaHqn4KtvWUWJpEJvE5JKFgczqhKGczGi1PoZMGd9KgtxN
dxR9d6S2VCltcKg9o1cPD2f05ry5LSZz0kPEZ2mQU2TynYX+bW7WcI1a0Lxgyfi30uByRqUY6aJS
xAurJ8kjbelFVEKGwUBFhA7BqMjGwoHz6UPKS2jPhXhxerDfbqryqK70vWei9vLwzegtJlZqRAzW
A91hhHGswjyIeaLR4lHbnq9ExJUUSk4n9/l3AuSUmTXJrmitLc2NoEY9pAretyxjkkLvqe/6r7xc
z89Fm2iNUQGnqaZ7ItdlUumbwV0zlesFxXpaWlVZbl9v+xq6p+pM27J1ZbpfSux3DHcAaYy+LeKE
IbgtQIYLSOCMjplgUYLoVUWGhSgEoVBeCGB4y+4bpjhOB5Kx4Fqw12WBPHCyKj4NI5sxLZjyU4La
tEglzkmehi/GbOlZrFNNw3CxTyhQSFBQZOPChLdQB/Vi7LdXhK4sg0/wCkYHQwqkJ038JlkWDcCy
qWMTg2l+n/4yWuc6JUOkNVzypoHMh/VfjEyN5+b8LMCkz0PFd/XGJvqgmto9Ha2SJBq4/sSUXt5r
inzLNMCznLWkT40oGztwcfM4rt0l+aIo5GMHW5gdqjd5A8I3Rhny68vbc0yWYxKlGd/jUo4nlAI/
QOR2f8AK2fuFYtiKxtvP+EIFDyyRjVSLG8FY3LxGvx/PgGKqUgiVd18QFQzF5m56Z4Gkz/TYCzax
mGSfVc03qArzPI6CPweupomb2rlHD88dLoRuVIfFk4Z+evZq2RtQvGH6YIdVQbULEDnokMdxkEai
lyGuoYM2biYj+un0se2OuhewX0q53/DXejCHEgZYdQ7fUc7hfzL7l1ZJdnaPEALiQnZgqDu3P4cF
UgjF6LTepDPt0uUAzAm77mTUBpUkLUbfe6TXSRgExPsoX/D33CwSo70q5M7R0RDSxeJiTbnwuBZb
i57W4R0/bAG4yDhYP7uxnRBV9ZW6tMnwmP38hrKqQSQyfGWHrc7WlRkVJvx+SXoGG0uqCR0ZcCDq
DD1EHIHh3hycq0K1rFwebh9KVeivNP0jj0y1AYBhCsQQCl8yHntzlhn6/a+5OpaeIWaxz1rJJyck
Aq3OGZotx6Jth0u7IwM9woaZV8AZ4Yi5a6kRVgBimthnXhNjjRPG0mieEyHgmNUp6TVLOA8ftRXH
6tNONe1zxTLvEzz8DevURyKaXRcXZiqspdQDBXaSoQb6QWJxAF3tOs+HgoZComNjbYjsA+A/fnQP
Qpm2RqhRj5g3rywnYIxtpFSJYJDg9IAP7gXjHxabU0EknUKn7KAlZuREp8yTSWlUJR7+22ATKcz9
sm0V8fjWXk1WLpEryqDuFv/2E18pbwi1WR7TajsMJMwhJQ4FkkSl9JWB9zL2Zvf9yM1LKBghVulD
wIXJDNN96Gm0RHQMfixW+CZ8jn4p/a39z8A8ITE9oHSXA+1Fcq/99zqZbfVTj7RLZzlroxVIhtDN
VQimrvKMYR67CS+vFazS1FZH/ywgjBxcQYeNPIqjCI7SnIrhzLFWGXgyWIX5upNwB1AFDcSnJaFh
zojJIzUb3SQ9mzeM57aaJ9HZdN6r2bLpm7Fm/0EHD5fG93ET+4mZOwCnNN4aU92GipVmO3QNh4UQ
4PzdSJwDL1RlD3XDk+MkGEW8rU3XFN1XcTZfU70iytBXGSs6s11h8xqyZPyJGeK2gLctQqlHVTA7
npz+HB8Imgqq7ObMwrYFyDx+8aYUrhBuEcBh4vsYhPg2nkGYWbCcFN6dDKoOZb2iVPCfmuF4AhH0
+2tCIgBGrGriUV4emY1yaVngklBBlb1a9IHAYiNTTIIxbWFUZ9NzK/D2UlQwpZmr9RFVS4z1aGdI
uXxdiNfPPZLBsYqQpB3kvr1J+sbQl45gzQ9bl5Bxd6Qzh/6FtLh0Hqhc1V+VjYdAHsjNB6D3Ct+N
PHyIFqT3xAc6dfHtyn/KrnW5aJVBsbpNjZJV+hp4g4gkSJIiL/4M660PlfjUsquVPjHCkOpaX92c
nR+BGqepqHq1hPMkOC7vI+MQxvT41WmZFsSc3yf/k4Gx0nT9aLFtkc5L9Cbvfy780jPfBKGSYTSU
mP2258FkS2JRm98nU7ydvnYd9PRWiwYNJVsez6u9Q8bFc9I0pCbSECLen8PMoaF2vV81u7L4ejkG
zq7NFWUf/uNCKyuiHZ0ekmBzwiJ6NajQ0ALdxNHZ5s6JU5Gj0yS+Eb3qLPxmINEMA5+AyIMwJGe0
Uf1GcaobmBGLNbD7l5ds5rSS8P3xa8Po4yv3RZ3JZCtQB+lFTpcXVcz91hs3JAJsvyLV4l8y6z9q
dxvRWXrcbEKYTdWoZh1iafeJfx/1+c4Sjds/7c8SUVwHUmBoBFz+UGfevxL2w8GdYOIECOnZ4NQk
nc/+tcqIQXuXBvTNkoIk3WMTZCcxqib8mq5omfeTkdY/3gglzyNqwtR5hJRjGAQv5nD2tHUsNqH5
wehCU0Ck6bWaXhDgW3VImqkHHycTc90Jx55+sweb3LbkCC0dldbXxD0oxaFfnO9hd6NlAEZJi4x4
dYGwhpgC06B8fbvZdJ/Or9ARuQ+Ao7McPjiG2RefY2Wt6QTldbOC65Wcm0XSnYRysDYbzisn8fNO
itDuDY7yQrx7yyxe/NFhEbFQQ4XoVuOZefpX0OeOo0imJ4tnGrsbXJOHpDxSfXNE0yGALVk/94RQ
4U6TYi7Gt8nKXtFWQiL9Aensywb6o39ylH/OPCkfwWc9zTIhNsjsKZVbVyE6Wo9wg1p/3xcbtOno
G2d+RZWFhmQB58qlKPbm4+yXshk9MpITVUkljS/kRQfSqmOWAMtint1BG2oaHpO6DY5Ii1AVs3y4
RiE6hlmupeOJSzbR5Y+VFwlThJbFIBzGz7tFslLqlJtkl/c2Ns1NdW144DtqQb4682tdafjeIN/F
T319kSGtLaXFF+CpC6d7AryvxwTtXdnPHsKjV0eJOjSiwSwYZ2W7tbEfcPYuuHNrjALWZJhGjmUz
emfjuHzRFAakCQ8snp0t+OtsYCmDIcyzE8K2arRG1uf3s3mEVM9YtutfvZc32v+g2T8Yo5qMoKyC
FMHEbZ/INGrzrxeZG+ai0aGhlGBXlRLRezpk9lqarw3S8dzMkoKN/bh4EAXbDskBABpf2e/zGLDq
DiALWufT/1xWXn9B4PphAe2bbxjsRHbspNgZ5k8ycNzhIm8JyhtseU66r9ve+4tJpKACyqcmc2s7
9HOUZx48IRtfiZ2g9RQriSHzNzTKI8BvmUIV7A0V9TRFqHKTnud5hXbalog8rugzb6Ss4tlK2oeg
ZZkDaRb1UAZuf7EEsx3aiHOJ3caBplewpUe+/n3PhZN2lb/QEc2dTaUtw97E1AIBrZwnHbawTyGP
0kMWmA28hvNW0J0D6c6z1Z6ZymvhkToaHtwr8O9DBsZTNgQlGkx1ddZoENycobztacF23MM9LY5a
i+5oC8wZtD/ZlCrR0Ee+b7e8xVRJ4O0rY80WsueiDaFxAp600Axi+Wz+6N2isxLMrQ6TT1waHRqx
suoiwZX7TIc1il4ewk3pXlNyYqsZ9dxLqQc7dc7lOpvWlIA382d26O9WYWczVmVq/fzl6lG42+7p
NZPyWnu0WovLt4fDfguT10Mk2vtrfreuxNPeSr5huuAXpPThMeuFT6FVjGmcvQ6hGf3xhXdqCsFl
SZw8KQAej5sDboATSM81cy0UY21J9B4q25OK276tcAVvYnzm13rnWV1+8XCY1DdnusyJ5gUNdNaE
FMqJjRyktCIIVImGQJ9cdaGB9N9cEUqVPVoMVYWS9rPr2aQTjNUxG3kClJBGPl5T5ZZS1LqLGm1g
+49fVZDdy1HcTZ8AF0j2Up7HkniiEDIxbVvbnSN13wih2QOtI3Wf0Ty39Zy02V5GJYqNf0OHujjX
2aIZUr3VYm4a5kbSUHecj7pCC9010QJGptCsDWiBgoKe5EzwEOY2iS+4W6KvcJip5ySNsBGj+KFM
1Q973NPo5/GsVXElmE5eD62z897T7Szsr2acD3iaDxnR0DuTFEx8iW7O4nu8704QYBnqALNaSxsL
W6YuE3Ha+KNgSSgUSSNO4ypGG7w/OjmfYJ/SRlR7JEZzA45hP4U9pbKLrdc56W5vpQrpRQ9HMwVx
FGxSLiWUI6MHAADaqd6g+VT6wKBlcwQYc3qYx/Ob12PIpj/6m43kQ8+FYcFQyHGc8fQzJH0Myp9b
tcMVOcmD6bRcIqlHgIJg2VW6ZKsVcVAdbatw34LiDCYhaWjNBYR5W7ia2E2mGlw5wQVkw+7l0EXz
UxzKc4Rmu/GNXxjoEIULF/Yjo2GJzIb45NLC4F5Tusq0dHZ8pVgVR3LXdMdVsReU2KUWzrlkxpzm
jfyAEvet1yAkL+ZPs3/hEH5PFuQWvGMWTpBlz4RIJU/rD+eigZRjctN73z3+xJ54rt9x75nf4ewj
NmWiClI1ToPcpX4p88yrk21pIzmUfRaEVeuAOAW+U6rSSCWXUTq86HgwY4+WQB0Innw9I3LtZTgc
i8f9936xFLyc6Fek7O17icJ5skrcYWmoosLHsc49ABKN1FAp4SJNQGYxFgpPY1eZIHvmUdlLWR+A
HcJ09KigjNfmJGrDZ6oyFE9jx0QycbqedntSTtcK8V+QktvBVcRwP/qTP8NcshyQnA9h2q4LiZcH
RLx3XDrDKP3NyJy31ClB9fgcDpaUYPTrsfw1hTAOOb8rpy2y6pGCrsEAFF9MAcEiCZs9xHxiWn3l
7SA2EdCngjLaJREewQOjNffhrUy1GK4N/q9fkI0tlHD3PuYLtsbuxWcauXOX1BEDweOup9xwBfQ4
vbl2AtZwe3lT2PEO0W9b+fP+aR1vO234atSdp3s8QYhjeC6+z6jif7pWP8t3w0bhftYQLcXmmsyp
UNhnw/lqTlvXo/7UfCdrsm7VFkf6ZXN23WeL3xdAStoXDUVcyRgSKGYlV+jrowy7sFv/vaajxS/7
WJAfQjn7xPpL0Qi1JwvDhLdoORU0QjHjBRWyVRgpEofy9apBQR0lFav9gnb0G9jW5W4spOMNKpio
DFkpLlfO6ncNM3sDTAOQ67eXyzPD6lfMw3F4ZwJVXYjVzuDMwwGpQWsQixmnw1oebjnApa6IXfa+
W8R8qlBRsMLYp6LzSOWeAYllpeRR1nZOdmW87svy9EryivoF5+5WOm66AJQJOLy6b1/nHjF0z181
H5Cbl50WXoXLaIlFoZ8Gr0BPcclNb8rWKMti5QL8hVkbWUP7qukwEnXo2ZsSfbK5urnGYoNlwSjJ
6mnvJipDwKqy65rIcw6zjnZL7okt6S2UELdPsTj1eldkUcyKvTZ2y9R4foq6kSFBTApwiuI3PCho
TCgJ84AV6P+tEHvtJt/a6Cclh+jzopWyl0NwDVSCxO2PmgezF9madrjXbCoC2n9nL5YM8s50rbJU
NKXaD4V1m+8lr3UbhtKovhzJCtv5v0y+9R2pQcuQzbrJ/Wwuofu0XmTAVj+qGQMznjS9qZ5yK7Ih
ug3uKU+j+Wm4hzO6QRESvstR5Gztfp/sBD1/6HxEypgiB3D6Wx9Gxn2dJRJ7J2hnsuM5oJ4m//Ml
zJIX9fr7L1RJULxNi5lj4qTR3I2Z8xN380Lcst164HwU2EL9Rq2VE5Wq/4OF8aX7cjmhjmNGjxLG
vQo4vVeeoenZHNqW2a32N0cadWqzz/YaU8dy26xEfYMwksroYHKgSogTn1k1aPSw/5zGp18Wvy+a
/ZxGA0QMi0LS/QpsbNKc7bzLdlDA7i8KO+ye0xeVQlpBRk5Teoj4dGr32UUiWULHkTQVPk30imaP
pN3IE6Unmk+V8ty2UVT5SZs2iK8mDgg84pQcFIIyll16kTNuHoi2RMsHEDwBl5fY0STXm9cX8eBZ
/JTnhP//VR9FEhXYeqF0wg9b3sStJ2PaNmvSoZWPN8WVJm3dzD4tDC8FEmiGchj+3417T7ysmX4Z
BeQ2+iaDWkQvtH33jiQdIGtOj76zguq46zIuXJjd9286OQdAowyTew3wCskTG7TyDH1YJIWhbfQ/
XxTORf2CdH0GuImzQRODj619hKNz/TcSza669XG7zAdcil0WcSsmnzKfHYWWksatfWE6W+Dg3i1H
siVZvOg00GMeoIe4FYiviW6PxnXjpicT3Q3IkA/ouNENQz/cJPmaNX3kasz+aXHLJhwbjYijnY6B
mixNjdJT4Ee0KFkF49oC69crNj7zENPw4E/cJ/hP2Zj7rTwWpYRwg2xfbRFazeAy6G5keQTJvhOX
JMW+GUuV6aznvr6wrthmRKNWMkMZEhkSbDehR9+Luj/NqPLsMUyoI09P/tA2xXndPOn89oPESEbD
312wtEFL0QXl3q1vvSHIHxUdZi2VWokjp/8I/1Kh3XBbc4TR93xg1OW76F+zfnc8++Ot+uHNi18S
oD8c4v4hlK4JtIUZUidpPHmkn4MN4+EgFbY4JpIu2eBC4v0Dzy3Xp+LpJ7xjHD8jqoX3FE6VyhcN
uT8VuzSA6kUzy+ElK9CtpdmVaUUElxVU3UnAOcv/n3pdquI8JlpOYpVxCO8K7/yx/9OoRjdG+SvN
3eYxJtzb8+ESWzcJ4GddaGcqbXOzTgHj7JRrBPQvALk1y17ZEF4011rqGmLBGt9x8rQkiSvNUgNj
avEkbhhLDfUQpNLqNyaX4psbaDfux/ccrAZCXNV+S5w5T112JYq7JhQFeJ7WSMOJFUR6zIu3+WPM
bE40lsAbEB1YSPp06x6kqmdQfe5oYrA+KGBhOTtlOSe5SKYjC8I7AYfmyrlmw5vIjiiz8VS5GkfT
8msS3BtLUAAB0/xZLMJrixVQBs/Yyq+XxV24Y81xNgflY8kheHw2cPKgYoPpdojqstqX6hzcowng
2u2VdAIISC4kA6RRJtY5Qr4zMuLR4wHNe3sHUdILu7+QHuXkEUSZThe3px8UnyGzEhfwIRZKHY8y
6L+fdLHqwcNkmJEX6zRa9Kqg8dHxW+zLHiQUb+ZeuTBOtoYMOzoETph+ib/Je4uUEsIB5hsblNkD
94QxOAOst5HlZfkA5ky1R2czeMGwlYLk5OdJUYVRuCO7wSElI5vv1UCJslYhobEl8I504XdTbP1Q
FcqA0qKAEYv+FBkf4bmfv1GQgDBUh6MXODxVn/R4HrtJQBj0scQKLho6ujD6JZ3/l9FeLGapKvHc
0wuh09yhnuLyYSHzE56fjOakuSCR3f8VllAHAuYufGGx6ojVTkrHM4xabR+cIUtBbcyuudPes5c8
s03mpOpHeTk5hvE3xAKOcQCmpYieTRjisuKdrweaUgVZRKMQfvZmX5/iobmRtgxRPKmCWdG2DGb6
T40HOpL+cnzehxvCpvIEOOQd+1LPdIDOHj5Cood23c1Q3/iisurDkRyJsrQva8CGudqegNXnXvgL
xAn8eIZ+1I7b5X5bHAQ2D7BpTmpuuunnFcrFszT5Co141mCEpcWWmVv1rCJQ8T6hQmTXTJLtEqgH
2x60J0KeoKhffsihoyVR4EpgRELAUwAtshBJC2LwE0vJP3bIg+7p4OtmFRQYzmdxIDHJ3QUkGNjD
jxBkc/ji3c7+bb7JBeiRuSvHtTbzGKrVgm6mm4hIu5o3LimR8AhgI2/gy6px2gmcYYOOUzIaO5xv
KoJhLZCtZVoMOTD7Q6EXL9q2nNyM2ktOTIxD1xAYkBiFirXepDhdkXe6rK+JpBVnwDPtJ4qGeEDj
mUsJDH5n1RA8DNO6NawRnJw2FqdVsXqw98zI4bo/XAvB2E8FPv4ckNV18lM2QaPXgC967pw7GvQf
rowgeLwcigq6LXhbtT6Z8nph2B5/+uuPxt+qsLayXy0Dr4nRQe5C8BTbuQymaXGfRhaQTCU/fapr
5jVRlVoFs9f1WNWwF4d/nGlnniWCvq4Zz+Y4v6dvs9amxpuQ+oIarFRS5nWXCQGC+kyi+KKVDihM
EvJTHDVS6RmjRQmS4MRAUVmvt4LKmYda2MOwx+oU6hG4NKCbcpTTiG3Qs58kqk+/r4ys3WZzO0Is
k1WsOjqLdTri5pQxM/kKcoqhoKKHlBdrJdCa63qyVodphDH5IkoDglFskPswNCitqDCSiXt3HQaS
OTlV06Vmj8aBH8eAIWCL5z3lr/o1d9NKG4SlcsWMtG6vb/mqiDG9JIM7AG3xseauMWdACBRQUxS6
tKDwe5ZWINCiQRdUSzoD72Kjb1FigWcN5tICe6yg/uAd02nBsKFWxPMwgSzppla7J3ErYbhHSaUH
K6Lb1PIMwoVF1Y9sHTwM8Vauw6EOWUsHozagfr4M26KZhtT6YHAG8zFCmB+2RjsvbP6mhhbdkK75
3Yau01+ZSA8ONFjE96DJVQZNRSaEb+xxH2pt9euNZcMcrikG8uuR5fXHtybyuMTz4s67kyqYY78C
wdcz86Geb0jsdluBBXgtEl8v5K9K5/uL7Wh5B3wReNc68rriZZCSeKxtKKqVOMeNg/0giVCInDGW
klpfaHvUgDOgOfWAhNWomnLMpvIGPo3AZ/IglLDssqPsd6Hh23XKwDvvp2aMTddzhO7B6FELm2Ho
yGjPiFWJCnwZ5JmDvIhK0O6E7aGYqj3CWCNbIln4GFoPzC6A/sh6KH8sv+2GWznCBGd9r+ifY2dQ
TgmobORnwr1oSpfucaO790RfhJUETJFWkKEt4EeTpUkcRp13k1Fgw9du8yPV1QuWZlkcg1t/4bwL
hsDQ+wLACh0XlEEDt85s8rrcViPK4Hb1yTDZpBsniynI2lr+RlGRD5mNMVey2BOM5YCSGURohNIT
3Brkb60kLHvreYJl7TEHksv7apZpm1bNW58PM3FDl6Ksz7PA560rRovQjLvnI6wMlznKGDkwyRCp
0XAYF4cyh4219bJDYQZET69kf0My4dbGrXHN04nOMBeTG7S1yI24YXfT9TAFYEXd9UIe74o0WFYd
bMtAugwWQUL/M9i4zMbBgJamM5YsF4ZHw6ZoLa4Imf+XHkaKTk9SQvFN9fucC0Y55ybF/M7NQG4Y
ivMjjNnZpcdTyg5rVfHrzl6e62H38rg6XvsEf+VGWSAaJM+gC57xum0MXDIqa/X9CY+wMIJ3ZJ94
dlEGe19rI8Ghyku03odbZLWjRhWHoA+li3xmRx0hJ4c3kw5VILN9INRPTyctKcLeDp0ReKCR+tGl
8dmXjwbTrMSvchJWtLELhTCC5NCP6rYGpzC6LfwLisPkaWD7nr2ZWkB3VocE+Zs2stmJ6ocw/1jF
OyVyrfu4so/WFIV0gO5RoKe1nPHnBoZ+XBVGFE9j/bHU2M83/s2P8pn/ldZWTdGXunLrBxa8wn67
sdmzaWfsiFGTWY+0U2tDHLp1kQHX58IScjL2A8SnefHyLkWX54OESO/jlo/QvPp52g25R/x+GdAe
DNTBQLSShjsh3S+wXqQE8CDpP71YuIiwLTVjFSoEu7Wt+/roUKTo1BbykoKkFcCfu+ok/bbxqZXW
D6XmlowiudcmN8/pQmWLjAYtd0IUH146/K0hRBpMwfkAxMy/NQcpiVIkXDgF5AgHFpEOuy17c2mJ
nruqbp0y0GrmbvN7+ZM9lcS8MoP8jsIzuANNxnQ8XU0mczY07db6ZCcWPxvg9foIhgPCrA2kdEJI
Erw/S1XvQ1JO4UtfqyaBKC55xIU965jiRguIZ1KUksrajhV0eJmL61F06fhYmEbf7fJDRMlnsHjZ
BXLmzOEcK/VhdjXVJsPOMurSdKyO02clV976tJEMWSyb9XiY++z5dlVNPcMOZV1JV710Bna3xqIq
/dF3whxcADpqL0b2NGHB/Cco58UqUUkPmgrBHbirFghNHKjtz3ZmNk6qrjlAmlA3S0EoanwoQnXM
s5++Pa2BQduUQPmgtQlmv514eNEEKj4RdjDC37DbTGHhngG6TpiUILYTe6Dk+ElVdx91QH+8rogx
u+hdHpXzXqhyL/yyordx2S6I7RVNea0WNbE8Za8weGPOGVA0FFNLdSi7ZI4G46dNMLxGjiSZu8VM
E+OLU5fXhotV0oiV+ooXdi+7n34i3qcuidXe55evJBR5Ts6zHcjYHHH5bz74VWD6aRKZ4XZ3Hu0A
n/dUunm5WVyheatnYPBTrikOB/mvWVYcojKQGqvfTtkeDr8MFi2OmTOFQC5SyPihIL7fWqgilqG7
zvM3K1IoW0miK20qF+8Qf7rhyaEv2h8iniww6i4fJp32xEdjoU5BO/3o1rrfrAYUlkPz8BoDGdhI
fC1TMDKVEc1zWT1mon4edFzhtbx5HPW6adRjOGia/LF1B7cG6C+omR20c+DQuAxfcxbVIbdz6nvz
ia0G6EqOS3lBJK44NrYSaPCm/gAZBJ+6yf3H8fzBa0ZBSU0cawxuAnykUvvRgxfJBsmfVvypLXCc
DScAatdDsx1JMSW5eWbOjaXj7ARQyLUdFupLB1EcpVVZeTZulDFq5x3pwlHLz+7ourlalECwZEup
CSzmEcSUQ2ZxqBvU5Py0ZXJ/4bo6uO5wB2Bd5RqT4M6GVBcAWXoY1wxNUK/6C7WCfwgxhKtSGFFg
Dt8hiYYTgpZHISq+HsvlcCXbzM/sVSO820ZXT+dqATqoeapAerGSABOIg4gYA5aUwZtAYVTH/nN+
jAhHCV8r1mtPOFiL62gWvTBmUgfP7leCvYnqpDbwVEx/HQvbN5qW+W7BYsHnaTZpAcLl8TyPvDB1
aJpMv+k/fiUI5+nduPtcIeldx0P2JyjmIvCn6iFqeLyeni93dbqYuCcZYaWxVONu7KaEdhY6D04a
jUeMB5HrqsnMsVqcQhRWjoDMHCJ7RPE7mz9zNIUObPO1VrsVQ7kpvdFkLYBYi6C9t6B8QsAHd2qU
jyzpgB3pkQzhMLmxmlNiqvegeQ2OzLeAYFr/1FFFxUzYR2mOpespLQyG4SqrsFJPuEiwXzQKMcwF
tZMi2XNK4uEn0IwCNHHp6+krv4qfYEBHWCFeZ2gl1gmMUR5jRtzhNziezQcEPMGSVsW9RJZx+yhg
b+OuU/1/GcZijHx4qYSgnyA4Q0deFIcLcYkyt1Nw4G1NXngJL1m7Hy8G3i9r3atJygNubUbKovzT
WBkookw4BN0ptyGYwreT2bceCsTAwUDPfyIrenHZBZYHfAWG0ViOEsvl97SY8EbZPDrMDNES6QfZ
WWoe9fD6V/8OyeTLH6o8SedvbWqumFPonOnSYO/qiPSRpx2Xhks2B8TWSy2yJJHJvO1ZapTKJ5ER
REp0ZxuU3C2s8sOYvVCbqZTz2TpAUQ1LXDIOJtmIamjVAhDLQ4RYMXyZ63iaRN+sDnqcb9Xh/lRs
6h77tAksd2u163nH4r8S/vTWkr+TDJaCz26rr5hdiQbFF4KSCeRzs6zvbhJhTykWpo2y5uIm3Xel
cPA2p/31LBjNd41OaZOgD9BCB6FgvhKPmsNPozrD+1Q3CLw/TfdMrPSwn/z/cL71rbURtoM+0SUL
qt31KMHQj//WziOnJg4DPO/vuk1F3cYLFnG2O6dfaBNQm12UDbg38dzzBgX8KuHP8aeAbM5n+ehy
O9Xj3oOhBhqWjCJIEX+yp6G7/ZCuKPlUzRgtSgFCbqaIrCOPLzpmY4DRhqQreUarSmfph0r+H8AH
PKUd6721yJWFQj6fau4dec4G46ORk3aZ4+MEql0EQTjqtY0F41VxYNuoE9vphwE/a4FOGTkO9w9I
J3RUYCCe4pX7MLLQWEp38qU9FO1o0T0u26fguKYXshUlMWbOJg0TtXHW+eWJ0keEbTgzt+9uBDrc
dOLiQbrxo36wAhbmQkg6hVqVYTStDfZZ7tCeg9BcEPhPH5926kNjQX5Bsetv7MOy9v9/3mWmJVcx
+bSWsK8luWPEhUGyfZnQcYxwdo6Aw4ryKItKu63fpvXFrCWDbev08D8EjDOSvMehJxGBOOtKZnz9
H9W2quwFTmL8ANPhCtF8A6QUWPbMWqllwvxcRfkEbM4ftaRX4FR6uUKiV9Yo+K5bTHca3URE8Uf1
JNpAfnQuLQ1/TIk2lRVQHsT/HYsaFCxIT6xmPpRyco3Hgk9QZylRQizdwxGuOsGDWwFJw/yCEUMv
48EHmvSKpiT3a2MzvGbBaDFzx76LqWBfwF1xDIAO9NiJbsuXBWkcF7iwJuOk1E3iM5lVyxRrYczb
iDWBsVJwT1u4XH6mIy27lolsbH0ZgIyN18DDCze+DwcjmiVQoKiC0RN2f1e9jFiK3CHVQ3o4wYEY
XYsLvosB6hsgXtgx7mP/e1icsedjUBgCz07gI2NdqlQrnVsQLMBtfvSgRGS46a2fkqL1e5jq7hCT
rwcIBkgdYR28tMSaWl+Y1tvBBMHrZNs+Z9JjQSsLSxVGh5asHVf8uE08fIc7FvQ/4pdjPl7HN5DC
M80GdGLBoeSDjChlSNIWGbVdTo/YmmJr/ptQinZvtXJtwdm+hZnh5HldEwOH5H+1AHPZwC8nSRkX
g+Kqu29H/uqn5uDZ6LPluUbEEPhQGMIwC/ODqAihMvKLZZZ4jnnFSVt6C6lYAI5MtNZfU+cn5X79
KQhErd0nUzNVHwysVmQSrgzVO3+dDDkv/rlxIiogDd3uF+Ap14/oIa45SgIYp05FAOAW6GbhOv5T
AqnKdLxS/hwQsrnQjUJHLmuont5L/lYuXaYcfoHI6NaZ6Z2CcI8GDVLO4d9k26NTQJXY/raMYLVl
Bi8UWiRic1LCEwsnBEUEDnsC7EhLQ2Z9NwpO/oZQa5dc0neoNt4rMqi9xUmxfE1LzXU+cQrNvw7U
FjfaROO3924tB/uAfaQNH5VhZqaNgnixbTgrNs6mbeHCjAUA/0C1xlxLrbOQZcy4Od0E4+droem4
7z1KIC6m7NZl2ZdxuSw+AgX3ouFf7pjKM2NOwM3lOEf+dQvBPj72pB7N5hnCdgPo470bM+rli5Ms
m92dUxfoEGLQZOKrdkT85gUdwTEU6gMl8Pl6+QBsBCI/R0Z48IUt8fYgbV37jsL+oWFIYcY+TvYJ
hLnMk7l5e+oZo2iK96eRGITpUu1rUIZBpZFj3XwPWVkR8WArC8gdODSe5z5m8jGU3VtfwqrZwoAR
Gbxa5G+UeWjbLtjiR54FoIis39RRnEFDSOqZFLf7l4tewye8ME7DHZ0LC0VOVaExqjTxE4v1LqFv
gEL2fZ1gHr5OAgVsdv7SJ9kDu/bzqh1Fm4ecpjfcQoh3eePj0UD96AMGAanPZ44gp/NBb037efUj
E7yuyhX9ZuqZubfu+V8NalC/t0dsdRsZhHCRWez9HdJ61xS6LGU266uR9kP5i5N3lEejeUsSVdg/
9d0uNbNyFWqvhAUBJmzQjuBY2F+pEZ0jsvrECli0vSc5HuJeKtOQdw0ec5ueCWg8W38fgjGlpr/9
/wVfzWDXz6qveI7xmb3VpXU5arN2bn6zscLNSwTmHKWhrGcQuFh0s756UyhGOoEEeE9gx0g92vcx
l21RX2al4/QwwqPCKwED3DiCB3vtXz0wm6ZmvFnabkiDSjBfEUBGt+Zq7J59e6Hsbl+L2ksZeLuB
VEUYxuPoFlB0Bo5Cnit44MSyLHCxERvQG+MBdO6wVZU5+VmPURbghWunZpSfl9GFlKCsrxdepTFv
WwG0pW47xYncw/CRofr4ClKhcg3C9W7RgI7OXQfPLuEx95qJpvDS8ivRYWgEslIOCJuDcPbPGves
RSZZYVen7hdLbnvFqkPSsnn7KxcbXRp8S6FmUbzcW+NpeJeqPAbIT1czn5dAUGnpQ4/nqguIWPHj
+MkH+TNTxZ73ARQMhS9QGSeh8u7ZrFWmLo82GCJfWSd7VAbbJQ10hnE5oRRelux9MuMscRNjHuYg
jI2Mng0F1OMjbTXMFNZfj3GyB8zToO5MXYuz4vGwtljZHG3VfHXmSLGUqMeqWrvZEHU3tu9dg0tH
yRFSlVg4DcWzMuIyI5etO/EmFRc6KAdvdVpQ6+Mn2MG79PchIU0LeeYmx5+Or5RjfLKQgx+tR3Lg
W34nzCWh+41eweSx0kzol6VLu3vLsZoaGwiXcHtFWrNwPqtTNG9rxdYwNV9Ai6qMm6StK5FlbxRZ
ezYCPOMigXyKqP/XngkGtUaV8iuOITb0GYzZah/TlkloWQHwp2QpKugJ/ZrB/N7Bb1OG0VcS/sRd
mLhG6wqsAUGvQ400P37a98QefoEUrIbRQZZq+CqmLyE5u5RiNwdc1j3dcPp/7MR/U7eMddNCakR8
pTmf6SLt3YasW/+dBMTvuhwp+9I1sAi4AxLsETKS+y3IER606TIRLmq/dZCdBLMuKpV5EyvBfurA
KLFrjwfOn15ZG0uTq1IAcTUtQGvfICjcmJv/HENiKV5l+SiNhNQrOjA85keU3FNtkP7GFou5IfhH
Na9B47UiOeYKyxveEwkax0y6W36BbS6aoYCTSCQVnS/GutgXdZwpSih3oyyh7SOGJ5v4xBcDjlcK
+h/M+gLbM1OeTiKDpLu9CeqBB/JGju39/FC9AaIs4PuhZyNzuTotNc9hxVZEGd24GKtQsoozmC/r
9dMPVqdV1v/3rGzsDuW9a1KBrc/aQooZNElM97e6i8LMntsRl/RsClyHgSfdBtl8BQUx+4MJh6BU
NGbRjLVXJuKxFZEKZL6+IFRkIpwwPdEtbPDMCGx0kFgdpsxdHG7jBmbynonUnGVdzyfz8OWH/bPi
yVXnHQp7sHOoozI/ZTO9E+WRKhWs5mhM4T3DeV3ItdHJCFD8AcrO6C4HHVeMa1yadScPPGS4KVXN
xFaPQUUnsj/v+wk6zYte/6QR+sNExBRvF/8alZJcWWOpAk6pWe6y9+xkW7W+4lQyJ1U/Mjbfqi5G
h+pKOOZy5/i9FYtaHKVlkedpUJtErRjckXqPXQTygQg3wTUlN6mbvAKb72jCK4r2IZe9VXJ0f/xT
kKh3g1LJRqCenc7dcyq8OfL2mGLKZfLecsfmbqzL+SwPlj3qdPnA1Vhcez6Ws4dyCmOov3w6btL/
QcLlS2J7W2UUq0T6g9xE9ajEtuyfEwShVxaF0zy0/X2JNV8PUqUnDZpv5joHz2PCybFMiLGBh3Be
cvQVSJcblTMFQP+KucQHtAEcs3ajBXOIhO2zGlunNurwKSk0NsL00NpxEOu8t0YdGd+tV++9eJ2+
6wqdPBwQ7eNfAO39b88dBX2vMPMSoUdcb4ztJPz/V86mGKMaQ/j/QIpvLC9HjwyKkZM+irmmhQdV
+UEY3MowpPRfEnyZgYVkNQS6C3p2b55MaecAcnMEkhB1sgRSoybhzzZqnUYb4TzdGLa4e3dBTnKX
pU1ZV67CmAhB6cGF/Fkwb3kp7qTvBxQhavYElxEXnostctZxIKILMm1w9sXlv0IVWmt1hkOo+Y94
CgVfV4cma0AAzmTPiZ2m5hdbzKiPDeKlO//+rdiQp3/UaM7Zm5iI+L2vu48Cf6b3qv6KotRC0Aqj
3QYJTjFcFkv19qvQ1Gn66ViLPuDSCbQ6hxV+fc0nEXjvo9blYXx4ssQtei+5nn9B0irsDJ5ki2AX
AlGwP51q/XmxLkS5AoBsXy5T/RlNykcsxus+6THn/zHZxj2NYrwfL2fEk7LSofDyjaIE5ZL0qr0Y
LUQIHvP5n4r2Mx0XwTGifRAaNt6EshMKPbsaWj1MWoBdxz4eSXBCD4tX0oV53csSO3hQpJDMCUMv
wfwfEfSYJfUslKalrnzrXWKTBQ06ODv4HKf6DfjTEUeRgy4gNt7yWyxVe39wSCdzgZ1UTXNuhztT
U3rskkPtwWO3WyY4daj/nzAk4mdFlZg9URVxVepzveU/eHuVKQaMb43gXtSoTR674gHODdwnFECO
/VW8rayR+ud3OxvIWEok1MaoBM4fkEb0XLBl/jvI9+shb1PTTL+Y41CiDcMTEY+EI3sp2bWL/V/T
MJDkwMg6cGd/hO4PA9wVNpmOu80D5ZZkq47UuB2Z9fMk+WuR+x6CnBvKE8W2EiA/qUYtcb3KZxWR
wBy2/n5MJ7IUefR/RdYHpF55p4ghi3BTyeRs1huy2Tq29xQJc4n1PsYYO+oZTwTI5K15TUJ3d5y7
f3azOh1ZJXs8ZilXdG+8LYSunPz1DoAH/b0zixDtsmZaMKbhDRF7qscEcRo0bNhF+TY8l1o883Ty
bwsxbfKupFLvIJ9vZDorNB+v4MugyQNWh9ANW8w8hmmISIBqQ1+kYAsSJisckShOmfdYS5huEnnG
msbwOMXLsJjWwk6A1VtgPDphwoM0FsAtDFXEmYe2Skq7vHPH1Jp0Kv8w30wMG8J00J603PM3EDJ5
fivJKTAq/L4QxmDPI51TASIqE0RaDeijx5JEbCOxg1QiJs9MjuEv1AihuMUsFnsTcESmdQWLzom9
k/Yd7njsrqW9NvFbU+QFp3BwB5y7LId6DUto/eUrrWhbvQUtZYtsrwx0yta7zDANq2fRXy7cwiwQ
6FEUBVgoP3gNWE7vXKAnQGHxIKmUn//CmuNG6gvHDu0QN6EkeTL+inLCofXtyVGeK6adrqcT/BrX
FR1Z/B6EGCizjt3QOtZec08FZ9eGXWc2yxwRHPT49fvQk/wGz2FuzTNDbahig/YIMDJyBTwelxvS
nwMkkE8kgcVTHL9D3PUmNVqNI80WQkfmIGpR/4dpgrK0A1q0UJX1X/onvG/ytkwyrEHMhRiSUG2D
67kf+FA57JkKmjuusecFb8jFiAMvqQlXw1RyaiT9WdietuGh0Zqo73iI8lAztg2kl2DR5QcHPdsb
WsBs1FdvIb7eipu/G3pxrmHXIPQFdktmpYGB6wW4/cxo2GQf6fZBeDEFRnL4/wFivFyDAA+o7frc
rOS48QrzQoOMrECk/6h4wBQ0Fxmvaa9EXiwaayZBYhyKQ/vjPL3HLuxpN2m+ygTCcjpztvfSpRqY
dCfXA2K1D50xBsaOH+8qu5j0VYf4PK9SFeFJUPVBCjpACPfVeEM3t0ZNwgpSM/orR1aK0cZ9YQvK
FXrId0OgKQCbTov+ORVsok7qGy32oFYVxwafK3AxtlnQnrcJpB8+m7eYaCn9dK/HX4KJSYnzRqxe
hmKc00rk+PlxncjbNpFf3QDOR3gdgrLd29eqbXcpPQUDsDg9b0/kACN7hW6lHgKHZY7G6B50+FmR
Xwr3qwbaa5hE42Pb4syxb6UQcX/IyUcVsU7x72Wzy4Me04ANXyxjKMGvML3Pj9WMTkPzd76jyfXA
jjQ9LKb85SyaECUpQPW5A0P8K0rTQBQQgL1eqmgxmCQNtz+HLAWCmVqK0h3USbbJdpugFUPuptuA
FJeSzV475QrAuE8UmAqQh26I6W10byJxkZRUXIu5joZmPUuJpvpDEQJOLcd1jGk0VNQcYWYnOnM/
tzBX1GNZ8v7CwDnG7E6wx/IWiYNNEdn9AnfWKyA5CsSzQy5HV1dy/thmYVzkG+O+EwbnWBwa4vlr
T9rDpMvR1kQkVNnu1KL+95pvvPiD8uZVxfmHGqoJwOHYzuZvYw5E94NGcQ46n1wCv+1Y/w5X42Uc
gLMui+QumJq6Dx2Ijy+MObKCMoY1EKAa9OXonoKqcCCvxN7X5cVNZeG371TEQqrhiRCr+6CiKWV9
01sgqpMfOkm1ufCS9/lrBxXPNymm+SMc6BJflx4LCi/wFRxetNevQdv469XPFLgWv678C5QCTgV4
UvvG608xe/XU7T45AWFWiK2L2rTH0j8jQAYertR7eg85TSZadeygp1WNGekWFwPEeQmX9Xkc5fAq
VtQHqLjNzQwyDOSmyl2/1YSbP72h+hnT+IGUZbK1A5AeQdsSVYlTbFcKX/z/vXCDbHZj8W1PQXBx
WKR9BZAb8w/p9kNkdgnThLOLMZ2HFruyx3/v2YqqX/959SCUDjlO13JQYdBnRcGtS+JJ15ai/7Bt
9JFb3OOs5WbVKc17VEG8vgqYl4tyaEq3wKI5q1smgOjCp07eoRumnQ+0DxhmMJUIsY1BoV/MkjVe
LsrnX7xipWPaJtkKDkyCRg7GtcWx8nDVA823SrXbmr3T36ojVV8tIfRkktCO/SbZy7e5xN80Ho4i
nr3AcanY3F9ZQJX2d2wkjqLhrpm5xBhsYKsqnSxUoNGYe/j2hURz6CFRmlIx6pygRW/wBAs2u3cZ
2rUvdkmMwga3I7GuEsMF8I1HOZUFD2RE8aSHFBQoQs8ZyFNoSjEkyLfxIv3CYwXFfaHmrzVXRHjY
u3oD2bPWzXgMb+XPRFSdb14MvRqPSKJSeM/H34rvg+OTXtAReWfxXj9AbkTdi2C65tdry88Kfd/K
tF0GTgWqRRDv91WX9JvEY482QlJhD5zgfaFXEhuCmMDf0Mkq0piWWrCau5sIw/hMKMzOwbrvIrHZ
qd8BhvZYPoSXAP8QkY32q1o3/q1ZpmFnnzIyhooM25jZALda1LE+YVntIC1fllppOewEq+/31Kxj
8DfsTlzu7h5mNx2xUrY5dtYpPx21vH5/+QSjc2dcPsB5mqVNc9QONMsTvrxh+Rppegqi5X0VnJ4n
G0qbvm/AM1OYy4CWFaLxni/MApwTKHitKBmQHa+/0McTsrtovvYXxD6VO6oXhKQI7A5b5f9We8CG
M2HeCkIxa/ocveZYIV3tM6bRL7qzLkU2BRJz34vl62u75CmZe2D79u2ew7tlUGcLcEdGBG5h3d4b
bUfh03muCuwxxu3a2G/+lpN/l+3juyPeJaT/ti01ZcE6Ok05448EXFUDRsUsxvx64Aavbdi8FvOT
7QecFui1lLP2BzmhHdxg4AQvKouxQYY0tLCP4+QtH+lX4BDYw7D03ssKzhIohtIAHOtAkuyojndK
Wl+FOtJTqHOj0U2uH0CDB/ahv7c6m00DHro4QBf7mt+540t/IRtSkfJ+yBczIVCu5bXnyBPXBZbz
SgwSFL3SbEJksV9ACd2ZYfc38S4q8UgeStMYz9rFLqm0HdFrFh5Trx6bbrPhP8nsay2KQ4HEwevW
fwZg/giENxm/aHCfhEoOUXss7k2/twJhm0xKme69tXW/aVcCE/Q0T8HqJWeACrld2gyZqx/n+Beu
g5/eoAarOQ/NBwm1y6VLQuqIVmd2quUYjfRmeLruAdmZYWyJ+N5MHx2wr8ZqI2Sl4QcqgoZ04NjG
Xnz81OoRvcONqxybxMhS+Yo5TIE4WwbsXrQg0Q/CmQpXJoc5mEsbFhNOMiBwpGPntMOXytMbZno1
vV46yd0i9Ot+YDIaWK83N00sWD2vEC2u7/hVNj9EBc8vJMs4k9dX53nJDWZSKa402FC3ug5ajXgT
zOz9GMtc8vZH/jrnRYyLYsqN3UC7k1HgUwUS5rmqo3LDSA55smSXUOPbsp6Y3Spw50hYU60rmTyq
aOPswlo7c4g/rNNZsgQhrV2AQ5X2yVkRQB2hctor/+iqiorNNy/S+5xIxFGkbZuoRHkfFgroVUfN
rQurjUMSU0MeqbQlTM91c/lGWhcKJ+eZFwVJsCaH86CZ0EP1iNeNOzUJGPkKMCBxIBkrWHNC/qDf
daazn418UWtQIEkgoeMJbtJmsJTLNl1QZKQrk1YMgrDIOrfPrqg9jgMr5CMfqmexKKTavwVPg0SI
f9YFONyxQDyMxG70oeIjN64Is6j8Awj6PFIlN8MGNIRbAlMHhCjk5OAQb4mMnKNX8qJ81MYmT7qv
VQB16tQhDTH5lUYhi7TWfz9FX56BEM8h5Xiiq2QLVENaWcHGJyXuMnOynx9tQc8HyQG8HY+XDrjh
gNlHXSM1M4lrvN9xCvNKNh2L4IWy4ZvTF5e3lOrINjffyPxts9pQfYv7lmooH0AMB/hIBV5mFgsK
i+qtyUgqma5BqGbP7Hid5aFzBTl0K8PsZ2+g3T3NSeT3cuV5G8kS30IQHmf0UugnIOyOe3QHeT17
B0SWH6L8nneLLVRUfBCnWni3TNr2o9VlHRa18lVaiK+DDJTCax8LPmbbM1jsXRtwyFts7qC+ddVC
Qf091BkpzYcvj9hMWkIb4Bc48NR5r7iaTp+z/Q4eAl8Qfadp+wC0fLskUI8e8Z6HO8Hvq3NJHHB0
A7j972LY6fa2RKxR120EjIHf3l2BAtekSsfSxGhCdyVGm2Mk8EdnYUu+LH8hnGyHFInidKPqkt4X
DFqmsq+6m81rDejYTV60iILWr7iOeSF9IQnZtEUklI+FB77McciLc3f6qAacFw3UHFAvrtk//9GK
kDVcHhPn55LQ4U/E9zFPmm74AP/ckBGd5x83DsGWIC7LidW/yhehz8Wi5Qgkk7hLP3m/ibTCK79h
ejXYcZAGTbFaWfeugVrR3SDD/9d2vYK+nvulvjz+tdwMGBCjXWIvbFT6mFO5KmWq74Uy8WXKw2D7
iE0FSRa+QWzBqFEoMxnv0qOv1Qcma4TrBJnDN4iDGvZ4gcjBHwzcw0hZJagrkYVfO5gmfKK1Dtx8
afI1VDp5OSDf/+B0WZfPv9++6luJZQUcM3d25j/FhpYCXO/E/yAOjStxk0SBdBm+P4LhKRZxffxw
RaeoAzoJTvusV/7QFyYvk54gyNJqz9ZhKYHNGOn1+QQoLpEER3TsjfzNAwnKwt2Ty8Xl5Kz8Baww
sG9l3uYm+00pUOEQpZbp/jOFd3Ri5J7BQYepm/T1Q9vfTfaFrLAuXwPn1k3KQUWUOgevPZG2jYsD
FmGBfO8JR64e8kKrC/Uk7rA8Uv4xy6N2JRsGBYvcUO5Oed4XIUbRFRV3mW14TAIkIg5r87DvGazo
McKb/Vag6nysZLucmjPBP3t1Vlh1aLqkYEdlm0K6/y7/duHYkzi92CfdjO5riq8u+dfh3+baL2LI
ZWajVZ/79u1WkVaYPueos3iAVds31NGH2C5IzmaZkL8Rg0Zv45Xlzkzto7KsidLIKhaOceG5RD3Y
nnQgj8y3hA5g3AsBVjw+bg6M8cIPv/eDgl0p95IBf2DSASWTLJTz8gZdwsRelhqJC6IfUU50dcTq
bWhpLzc05x4qBYUb0+/GH6dr7ZP+TCoPl32whqR8Q2mlpLo7SkMBjzJfJYApRjy70Bfjj5Ax/WbY
G6qPshu/uNJkQaImsCeTZKW30rPYHCQaoy9bcWZPBj8+96HIyFbSbWvsHRqaQohSM3fxcstSIS4k
vRmNtIgnonPD57QPDFIPHsWdia6gjcMDgnyCF0hqv8Sjliy30/CNcNYbF6nzfSjSVwMAlSZRXs0G
Bu8Okp/K0XCgEWBdyKpMjbifhnRqqmn50b4Mc7UAwTXdFNiwJCoOOudIr93L3UO+kHAkTI2TLV+U
FylkHVR1Xttcu9H/HedFAXcxM8YV+5PvZ7T96dOcY/SjB8MRETk+mBmMUKisPKjej0D9ChEyuDmw
GSi5GhXcE32wsM00Dyi1az+2P66Vwfi4Kcs4Tjp76Qkc/Slsc0WSb1q9N1ixr3uBy5rj73gdKLyF
cVk6Ijd2y9ixGFqdhDgtDc4q1sQsVBkKNEidd8masXD7Fih8dQvKaxK4QTqvDo9JYBvF52u6f/8l
OZMzRvidxjvmm0qqudBnOFXBhoxTtEAi840APahsXXnADjynHLDFhc0gAsv05Iwt0YnA+0HYG8VQ
s78Y9SjbtsnFo125KDygCb16F4Ig5nDk84Wp6SkW3QMP8F3Ml+b5v9EBz9nDRLnezZ03NJyh/CGa
+Lt1D+2Vhuz4a7kGQjYfTOIQ0KMKzFMddytU5722FZC4tmNu7sTji6sgFE1gFjDDnukws+vJ9sX0
+WlJOvvYZMlzBO0G4+tAqcMcBRLEidc0gSe+ioEKtuhv97XWgSpEtKN4lOl5BAgJe5JgkSE9z3fs
nSqngfREsuSWHqdSTfBJ529NggjL2/zjrpcZBNbFNrvZH8MBhWm6kZLi77ah5NrM9DHlcZfis7lv
jLC89UZFSqNFVwGroAv5W5FDwv+AHl8m1+RAcXAB38+G1Ntg2kJCai9y0ALpWH5jVOH1sefh7X+q
W9VlpmmkgQmb3cGpFmKsKKihQM521iayQm62dsRrl9b3LihoT6nWk1LlO463b/grUdSvjObtNjhb
rdmdvDMkRVsNb7CLKvHXebi+Ats3Ewd1b/KjEbRy7HpQIGJkkV5FxGnfd/D6/qjnM1OE7ILtXfvH
+wYL0wsUqdSCucDDHrQKZfJl2zFdfDZ329kOljuwMvg8d8C8/uj9+nZRtZdrtLxgCM+72scAl+/f
25kvHofsYP4IfTKTyDLA+KB4Xgdffi3QsDmtzgc0SgZhv9qAS8/9qJ9iLISgRCHVhpWtwl/fDxLI
wIfM0oZ2di9UoMojc0q1ZosfMMNmQYMZn/bGjaXr+gjsJvRCpDIHwH+43HKaQg7l1ICF9yqj65mJ
i/UxHRBIlVdZmpCHk+OML9Pjk7jK1CXNJx72ogXw9g/K2prC4gtpvTp3Zs3rwn7Xouim7ypHNMTe
bwqJ23taqZ/eMwQQ2I+MYclpiEtUTXdXSzIseWCIJ5oIDCgu/QYf2CoHHVli3XczlfcSbtv/k9Sa
C7AF4HYGVk7XoDy1uY6HMW4Phbtm2wJcjYxjPcZdDmh8IXeqKpbXSpJNUtQXWDwUjdQ3cE7Cm/0R
EJnv3mGd2IvlhLaWQv1FRNqBv6r5uVIKFrfmHJfVRKgBfRwSXR3lyNLuAzsyIQuTabHmZ7lAwTtE
FAe6UxiL/53/8gdn9sLQT4alX+wzEf0IZpsFgFwVzz1oxFcm8W+kvj0LCTXAY4qcCbkep6CnUyS1
fOgCQ6pFaEL2+pVrXlzQtJ1y0n0wFtfBZqm4cwHDOM7jg7gKb1BDCBD8S/D0AmGwUPxpKcV5Ss3B
QGj1oJQk2VdmEE9oM6nvyTAyWX3gWtFFSJkuDL0aiV0kkameSmAuEX0SdfoEdBIHLz/R1E/wPCKI
JjlwaljPKS4zCuwvldpTZKY93YTrKxbRNcWmWdwbpJ3jddW4VfGAvhg+kXXGWVYf33wNypJB48tS
4zVA+M270Jkp64Y4ccQEA8zwCEm2BlG0Ls72wlxTyhRwAlzNdKT9Stis/pwfQ8/ZJ/WP2klT47op
CBqH416042dnPgHCluNZBBMlBiga905Su2m+4zW8d9lg5fauTIuvK7jSQx84B8kgA1HQT8ZE/9if
T/88SfEBZOurtStxVrxIg8gqQgZJleNVEJH+6NnB9B+K3VK577KIY5aHLDjO+5w9xyxW6UHp9GzW
VS28m4YpdtAqsywk1p/tNS8OUYeWeu6O5Oi9Z8CBqROlNgGg88Miye4P9y6SS0WnJu7rGvDwvRrj
45qHBCLAaO7h9REUrnkpo+M71lgr95pJn7Bh9RV1hFzbNL7Y1VtL/RwLhM//5OmctpAmHwiXp1Lz
MkGMvK1x4Sz4NUIcUDb+YH0uHMwWsMX6BjTdHT3ziRhrzzaJv3JX4DDL9W4Kx3GzyMpXNZnNSdgj
F71YTOPWryTVgfl81sXRVeG+2heDxRMYooAsjqx3jJabI2rhZLQTL1+694etPsb+sFv93MMWzLbD
tz1TTyCABdhR5Qv0SdxHx3F+bPFjqYS1DbXVdkBj3/myZt+4SLP3AjtHcjQfvqynWKy7/v7kV/OP
ItJoSCKY7ZZ3gzXyIhMNbrQtsk2BkCfwvX6Bn+xguqqvMgFIb0bPp21bcAAikQVl5OkxG7ABi51f
OC1ijrZpxcFE/QvnwkOsyHLAAOLc59ikqz2iFz7KoZ6FzZZTGUfYaXKcxe1vzLq8W3PQZ/q72yIn
5iWJ2r2qtH+0PEZly5VouNQOvoDzazkDdsqcI+O4yW78Op0JgX6+EI6KQHhZ9zUtASD3vPRUkHGU
yr9AIBy/63SrMeF/lRo7BVO1SfF4/5Lfsfwwvx6HCBH+79jgoI430LWBd8nroln7mOG+C7hnFW1x
braSNpu6ck8ZLPKmpjtkcUv199mthqMyLFiENydbuWDZiM3IJMBNuwsh3GLloe16iyIy9msf2wGJ
DkNA02eQRIRWzfKtshM2ji/nUfgKmCueYx9iOueSeba6uREguC54REM79Ouvr3aYgHUW7zUz6qf3
+kyiAuQFyQKF827w0VnMEY7EbC8eLj2kWnG6X+9ZcBGTPD/xcsDh5yujSCXn+do9xYQxyZgMM5mU
6wfVEC8FVNhKir7J4uTfdJ2aIZwjBWuIm/AWbgzuoCC4JDA5IYDDeQEfbzc+/a8j0uIewF3fG2Pl
UoDge1uWcrPQvZphqKNbKSVNFiIUcErvTbtaPgt20Xi4ZbTIWjxRL21DLGh0HLfeTVNdLSyCBLOF
rxfwjZce0Ozk0tT8+O2qOYJc4EQ4/tFbiONQ78QB2KqjqnTrRnpDtojSTm+/Dg+iflZf//ZVMuTF
ddgBvUFP8FzMydCnCE2D2FG/PgtztZY4wV6Ouc3lqVdPmO0kGlbBfCOe7KqXmJ1AN7XkjqJmb7iX
8bt0NsY2+i1B/LedwNa7xZkBmihOA7BNalZwIxPiEz11KXI5u2k+aiBIJE5GjVQa6+CRb7qxyXtY
qpKc9gWs/aAF1MqFDES0ARLtN8RHWZX4JP1Ya9wuJfKyeel7lr5FqykfvMNm/BsIGKa8IyWU0m8q
xFfdVlyej5sM5DNnR1IQwvm2kg18Vov5CV1drpL8PYvlwXBhdDBWaWRAhqSIVPNJ+evDX6Uwv13w
ARBYfPyfkuBuQyGz+N3eyinHgI9PXX6YFbhJai4Nh3U+pHQjJkS+l3nvtILVswbldD9eyG0LL/hc
e+FvWHo5P98TlYWE5uVyZLlGl0ZNKAn2m+aySPNc/j+GNXdy/Gln2pslBDT3s+5V1/inqM7/YZrC
mA9wGEa412xKPzy0ihp2XTmYbBegbV6Ok5l6ncsXr0Krc/45t6BZ6MkDu67jsib7dij7+K1JmwEk
ZuwUc8mMCUPW0plEUePe8TFWntNhg1GadNl8nm2HeyHesTjt5eDbQ8OhqrVmuRRzJRNpkv344Hup
c+VcDO/nPaiAbPKcwycNL8WaZPCSBLhdHYyqszCXXJktBwV8J3jYlsVdDCK9rOBxoF6it/J64FuH
eqlf70JJ9hjXDSbncLPBggzG93aOWG/+Ox7ldrOJJPYIuJDf/tBKa9++q/PqAvqTNzjIar1jVYmK
RjznCxv/IZb4/nnDHbCk0ZIyTB2SCHJLrQmj9E9LBXL3WvFt/dEin+2N795b41zjvHTf0a9UHipR
Yqk5wUhHmx+OBDRgMjSg2xM1RR771sEQQw+Lr77CqaeOc2MmDOAIQt+YWHZYA7TFM5lRTPpYqDoR
rptsnELglTwrb4q7e1KAUnHFuT+UcMFdwCf8bSZCsrJXtH7F+Aua/wBCFGRAHLw2vG5as15TuQxM
lyxZ/X3xHo2XguqPLiWuFgTJpB2MVR2HIxTQCvGJyC3lU+N4sahYjUNXys5p5p46B0AKAnjPu6VF
3AOIf4O8JlaJusA6D34bededpEQv4NmnoMxIv15Pu6e82FYM2UNzzi0YlX8ex7ZNTrvEneNCZyv1
hHX8scrBOy+HzdrH4bU9+yIRP6j+nuj+/V0YKe7QycvhC7rjsDJqBliXgPJT74bKPdfo8TRJI6VY
zjfjv3FgMuYGtrpbSioSLUTlcCArM+Xh+oHYtbCsaFLuz7CqxvTdG/aORKOD9NHIQf/VSaXP2Cie
0Y+w4I8DVpl2Cf2r79yRks6enf+fYabuwb+SS/4g+XO4HEBltpR84J7Edm/gLmmjePjeZiUM1/M/
usVKf9L0Cpw1Bnj+gzKHXhxh1w5Iliqb/dgtkSlqguNawjASiuGx/G0t3Puspw6UjUSQd8Q5HZoo
WfUkEvK/7KlhVN3L62Bdr5bIgcxnZ8H7otx0hynO4npZaLGwTa5+RC3bVNu3rp5GTLs4BlEWOAqH
JrC0uE95NgARz1fh3RrHSHnTAPHKWDCqQ0Muc3gsWHFwXy4JJqNjm/cNKG1c7G70cFHzQ3+TZw2n
6bpN6rEck33sG5I+GujwFU9kOThRvgK433b4/QYj98Y1LIpH5mWGoKtv/MU75NrSuoZZ9dJNcqlA
9iJQjXari0FeeGHTcZ811WRwmv4LLBPsxwbKIMDjUVVMviT69B/sMRZzk+EjVcmVj/cggwUmDL/s
e/bGU69RLs+48eTKRy5wrHugYqYU6g3AycHP55/94fbn0fIHHMwRe97QHbAZ4HMnyxQ7OxexhCYo
9/W7hnwuyZzIPctCM7cV0xr4JJBbXzO2RN4X447bpvulzGhy4UMoUNn06ZvFDZKVEdduI1CskrVg
0VXEyflLj6zP+x+6M8mLM3cOF/lbbi7H90DE9hlc11sPX2h+09r0Ea4dMw4hPFX2vNJdGHMxRceW
PtlAYfdg7AoBGFlEjLyqsxaplykC1mFudeVRR41Qm6tD8iSXMQGyCxgh6NhR1vkfzSmdDndLIDsY
qZ38jyVgX5AhoReZ5O4diSnTMVilZtCdUQay35vbLb0sbbqDm1+k1ecz4PgC8SI3jlJRqwXHc4p4
HnCZ3u65bJTSLWu2ZhDLYey5rLE+M2I69qShTMEy0LAt8UgBGy4ZUWaeoiuTajiC/DUdviDvLHjQ
y/bBF5AiBUsENkcMaZHjBZ0Z6lxJp07zl3xLzCbTS8jNnyy7+4xCUDIeS6R4RhTk/uqBm04H8m7k
eJmnh6GFjYQbATz7thAUxK7VPiLmS3Q891cjTXcm+x/BKM6+k6RvfENp0M6ZtdqrfBPv4D/fs2UA
4C/vJgfOS4SNBzJwuYfKtG3Cf+EKPTckjOTRXetac6lM2yTHssnTTPiuiFPZrC291DBi7yqhcGTW
Jap9DcXjsWhv6u/mW5UUrbL58Dl2Pdu87ZfLs6p7yCePTVlqq0a99eKeLXmpTlVn+9kIWqMw1uy4
ifnWKOEZ8aXoFpJrPYAzeo6dzskJJR4YFZubdOxj44oUKXS4R0Rj056EypuV3LhciMsHbei2wFz8
ocepyqRBCXYwtPwnVPuu7Vhb7gH4waUaooxPGDnLBqrH5aTL+7sGqF5M8HIQlvEy15ONpqK830Lo
CQ0UwSl+twIt7ovkfP0YCI0/NJHkeUW3bd2o5bJXymwQ59FX0xKxFguTcoZ/FJ6rE7SE+vLlejcE
7Xuq+xlhoOmzNLkLQaM6tz4VN0piFK7c/BQHvekcnQZJc71FL2maBUB/PyWvg5uD0svlfqT+a9/g
IjDj3CIeyvuQGf/1SZz4p9c8SUgsT9b5gsNAsrkk+fz84tqVbxRbmS2WbIk8662A6DWV9OwXmsR2
T6aMABqQ5d0Odldin58LFdYJ6yOcWIfgVcqYIPdgz5AU0XPR7udyMGUd+P8d1JHKYvbo871J9e3Z
KQBRYjA/rwdNzTgqTi/4B5PhH7GiV0XcVEOn9ki4GGQoLLxgdf3/Q1PAf+ghgd7asPo5nBccyBmW
Qb2DWYzXYd15exvh22yuf91QLcKM+HNEWivW9FfnyU6bfEA/0ugKMWRwdJh8y/oZ3um+unw8x8RB
Sj8OwM0vLUmpqhwgFOC8LBhZow+1K85fR98uvcGOMO3qdbIhY2AJggnPE5T37iGcYR5sqe+rVUm1
ItG6+dct708wsjWAvABsvC1wXQG/aN0CW9F85TUozNt07sVTYLEFs8m3iTZbjfvVsPPJ50IS7gDL
efkptFThmT+dbyYLUBRdpknPXDxxyxRRw7YBLNdTXeWiHnJYGP+VOdS7k8dzSMEf+LvygTYRZD+s
konuBkkAf4HUx1ibyy1nmX7LMVeIQ++iX7ztl0px6YAZPJYsng1R+kM5b3to51y0u5k2NlLdKLVV
kwiZC3SFunTiURBDwu8LL2SOO265NXRw/0MqL3D33EI7NSJUCMZ1popurqAALVurN5TeLAziuP9U
bUdZzivmyfYUIeaBg3jtJmvTcTp8mOtMnyS4LeO1xVwp0ywsui4rPkBSMNx8+jzB9Mq4IQGHPakm
wnCadHCBkQm9pSAlbCnQbpLWPjb2neWTWIn+elTl4g40t0Ppym4stBNdOsUDdKZoAaM8vKrGxmdu
bWY5qyXIphZeghQz9k7p9b11mjT9W7suxGep2+dVZBUq3W8Xmrj9e+6HyQP4de9vLoHt2OSc4ZIj
7y5ySb9UbFeahAG8k7pAJxbjjHDbS4Hd+WVCitCy9nlo+5M2/POCmL1oSkdfoK1p2rwn3uZi86Du
zsVb0tAN3IsRhpgJIU8cno6QJNbEHQYgyz4JP8ECPF9rhE93LMERyFpVkcsw2RnGpIMm75goC6Ir
4MJ4grUXYSaBlgG1Ccp9OWVikXIDEVdLPOni7+0PXYMULLv8CUzH/RFpyOO+h5tvz+hRFylJQLUI
mGThjNkwJmQGIXOv03RC1IALpyw12GrplCv1n1qpoakCY+IsGziBOQEdFbPEIHsvljAtj5ap3Rjm
oxCF377HcGAkRRcSosZdso1uZz3vxQ3odtJX44CE3BThp+YIuuYqXi+qKwglSzZkDEVBOpny9BsS
gWazq4j61cyNQ3cQeiW1fA45injzYgtcVFqnue0bF/YkAlcnRGhmh+wKsSaIIChl/ycFWRhi7wWF
A/6onzm+yVoVZTzHQWouZ/a2qgoZ87i9k70KeHlFm96yfUZ77lfIWdhj6cN3/cHPAR1joPeS1Gvg
9e5qy8UDDRjcM1L7g3IvvajkA3OG3mkRTEScmlD5n06JJwGWyLbwEBhak1EmLxT4Hp+nVMlRdjE0
nDrMuFd9KgeWzZ7bY01XMQBiOPNO7UwY+dejYHFbTkDQRM8WZVtbCoAZfUTeGWLg2pfkCezAtrYR
mGmRtJChepqwjYfDNkjNGiCe+nKEYXqS683YtJGYu+mEZQKgITigPTwbNFxcV5i2c8bWApkLj5eP
5UXJb3OWiU+219WYN0puztU8cxP6KIOhZoHMQTJfgViUzcywhltZcJ1mD5w6CknkGg0S8aDDiFWX
lQi3pN6lA+jTBlW5Qwf4ISdd9q4J6qQFIv+Vw3EEE8DPXtXHqE7bUadWtE3WHmGZr9j/Qf9wdKep
fCetZe8ii7QJd3wyQRUOfxRMOws95CzawhDCHKZb02wPUJbJQJroonUbAS7j6kaZeZPvGxBd53/i
XT4obC0KgkCh8jj16leQsHL5AXk2j3+0KPAQUfYBuKf3+wCcTaaJZpNPerIXN3iqe6ukCemlyIHg
5zeb5N6RN/UpdlCU72/dbAFPH9rf5Q6XZpl4Kdtd9sz6K2yRtbcyNfSAh01tGz+6WT5FRd0wU0B6
AueIRDmXFi5fpaTBgT/oBRAZk15kefIcYrgiLm12J+qP26Detv8X+jecSx8YasCgXA9swkcqvzyS
ezY/x7dJTwD662i1YWrjCJSEUQamlJfe9zA4EJGlEtSAVCPlmjY5vmVHdkDnfA+blnpn/2FqpIjW
jsTvsTGhEKu8i7m5mwSgVXCKUYQFUAUNfL73DwIUkkb/k+qeerk0AqCDRmP+PiwtJCg5aHjPOEFt
Di1MOdhYphAHflMn9buPHfreGSo5uwbS44gE/4GUx3tL8XvE9TQinTtsw0uY5E1Z3h7qXp8vVpw3
3X1r+87mSIa6oaZmxLi61JykTN4HhjSQS+3eHKwMGbf4Cr6z/3/mun3tiWYSwSzfN0aP+CheDCqP
dUm0Ia+aEM/lIyPQ726mAmRR+OhEtIGyPWK/hEciG8lK9+qQeRdsWXf2Y8ph3kXGZebMSt1Tpi50
js2F0QM/2n6wQK3VIkTATjLoSuq3tzpcBk5MAUuAA2xqfoew/jnhvTsYHnkP+dKSNoRSaZ3njghT
mZlQTzKO8NbleikN9EiABGpwQPgY4SZijIQ1z6t/35Rbs38AlondXFQ8AP9fy2+pogwXmntDM+px
EDGuPuB6Q7H+9HqJ+/sO3xWbLukscI02s0znfgMaQ8dmMzfV4wklvHDPjFfSr7c3Hv3MJ7B9yC9q
GoSHL45SJZXtjIHtH+310JQ2KvFEPKax/gDRbzeQFfJ+5VgWx3hFzNavYAA/dJwAhyWcL1fzpQdT
yourp1KauVWAM8ej4e88W9/ckuxBvlJvYdFPk4GnV2sIMHCoOG066wt2MXbBHo23RVtg8gQu+75x
kgfzrAZy7juFizbImf1WuLKMUPRE1K0uOrCvCdqPz6nXhih33mxXYnq4oRURgrhvY2yZ5C8OF6Zg
xPWUy4nX0V8qI8sdhzsZjMEzhegQ5dt9BQ1FZgkfg5x2zAnqt3XFcfE7pnYsEiq4cgaGd5Rpogdx
95xmWFxf8vQQL5h2nBjLR0iEl55YF2oIvwwvH2ZQWjmvvFT42s8MuDWVPtXfVOlcjbk0oYSAnnx2
MmUbH92AcGfdr7VTchHZfed/XMFSYJcFUGBA1L5AIHIt0P4vaZzhY2XJHxFiwh5bFdN5FEA6h/Am
0K88RfoXrjWAoN0GxRmdgkgFBgie6e371wGwbpongGPJRy1c2fACMWTpwPTdmydfKuNEBlJRfCuS
rJHpLB/Ibzj0zVUwk+FFbiTt0lw5La+JDIwB10ww3CJXBstnVGpUn6vWc92bC5r644qiqUPfxRp7
oCQiK9VWs1wMUfCjyhb23RkKqr5UYfGL2xCAyEAQT9CM1bVeIKYFR++S7+hwiUtT1MgTE+Wa6sSM
fYQIFwEmYYE526XQRQpPfE3LpjVLM3TylQLnGvb/bTlJ3OMkd/Hy14mvftCFQ2ROlDjeMfIDPpj7
dmEkebH74le57lAFNDHwI4KIPFVswSupiJGKW/4o07qqDK8q3rOy/coSSznwasMtI9m0IKQi5WGu
0bhf7btmnrPF2LkItXnXDPSLICI6dT3Xj0HBW36d04MJ6NFpooN+QcmXWpDGXMiEfntSBTjT8rbx
NST/F4kg/tXVp/Txm70HnX0tBT8YO/bBeH5KI0SYIyOsaq0DQMaBXJuLWAJJfOf6++JJSeDp0Ko0
R07iRtPqvZ/bU2r+HU672ct/UjikdnjaRQFUwiUlkv0BnXmky9q7hvWoSGHQ9p091XBv4EEfNvyz
xBXiaDezi/0sHj7TTHFAoTvjIxj1GYCV3iKF5ysarkc06KBzcIs1XaKKpDlQqHswQu5Hp1mmQzRz
LxeNm3L4ET9et5eYrnUaaGSWziF4aYxsCeksWW5BPawgFwY1+BfMNumIHSNb9wjMXqAPoDfEJ1ts
buxu45TP/Ln7YpX1Fn3ufFpLjr9ErmOd4r9bQTCpM4Csgq7FubT27gQfy6rut7P8wi1E0JLl9/lx
nKo3idv6O7iVj4oyD2ctQs4RGZj0bes7KhQ+LffNVTG6Vgc5P9sq0bAe6O770Gs0iCT8oXldksc2
0F2lR9tDd4Ocy6SsXaOZqDizvy3KkATJLyUElZB5COi6bgTnt2tWkitoazdbmUQhfsL22VLWqMr7
Y51FYO6LYKYhCxyWVOCFqMTpv8wTR115PBH1r3CLs5gAHsSAXWAycD2MI/a2NaFin9XYZRNlD5oe
CQxNJUkRkTExqJ9JWKyBdgemQblV/jyIFx64s9I3NegaD8/iLSoR1aplmEq9OUMR5+66tkuYL6zB
tmEat5BcI0XZuhxeUjT4UQvBGIwtu3wdn6NB+GKtxVX9xKnP9IxjS0at/R3otPUQQ3hyEiizddv/
Hk/4rtnDep+EE348Z8zRUVUWswVj80CWNW9cwWBY+q5/pnnvFf6iePas+HyA3tQD7qDmM/ctBCd7
B6c+Xlk3KyB2vqrp+FNW4g2Ug6ouGRG5lo5trjUTyG3WjqBd9TV5u5m3K7IU03HRAeRtv37/8tto
pzxzbkU1LXh07/p3ub+70AlB+IKrPJaZMJWSa4dADQnWXx9b5rZOZ4c3eheD1m6AoaNZENkiM/Pq
XwJm2HCJwvtN4pSbv4rNV7At8zoEePs3D471mY/fZ0vmyDC8VxxvfPQorr6P1E2JoMaEo7u2nTfg
oqwWrjsz9TOansm/KnPDQcjTCYpKuCW6nGRqO7cHt8afIzE08do69cSUGAGk0fF66g6GManO+PRU
rGc8dFywSJxOE/C0mekKgd6cfcBhrr4ezmMckobqj6+yXntFk465hLxsBRmRo+UXTtrT8txK3Afm
yRq7+QOuMlFD1Ot0O7xf7CTZheLMeQFLt8i31OlYdTfyt3hYMU/c8Zonpi1jtXHxj2x8p0krsC2p
lt+kMiPOdIB0EaAEyU1NszBrpeQYssuMSCWFYH0nRttYGA7lLZQx2kfoQ7tyImIS/5h/WDHfmtn7
qYjjMdo0RJGhGD2ecsjWJSVbu78cqtVrryD13+8EGZmwjkzXo62ai14NzHSkmHiDBqXS0yLdKz0F
D00kIi9i5wZHq0PSEuIgNSeDUuvcNwbhVBimL4U4rJvGyUWZMJsc0eee43b7WVajFZyF4cFhQ1t+
hTl/afuAxgcDo1MmT8j5+HTU843kSz975s+tSpOEnjFu9QGdhkh6jPwIEWPQBuPubR1JBcSGfZ+2
3iS2dK0TDWlGP+dCEfZpji/gETlDdvN1LxHs8sSfBHUChXgmryouMkUFuSuuBa6chZ3XOD7BJ/GO
29hvMrWcVwjEH+nSdkVKHhHUxiPA5OfTHHc1eYsjRV4lGbFnVbmzQzYs2dS2qiapjdPlwk4LA3UY
hVWduCAIVm13qima9kGcnMtVwhx9UwSXCyMVck0EmiYoIdk33Z4qGVoQ2AGAQFhQWZ/nkYaYxmGi
WVX46Ifob6I1mYqGmqmnWocJFW3gz+pVSbXJWPPykvR4rP7ruaoVOufGgXJ3eLESxGxEfnIrKjMW
e1NKbzubV/9ILfSUcvb3pwJwYQzKGOrN2pCUmopvGes93yKAuzdB1VaVBciHmspRNvGisbp2W02T
a3gMbt1dAbfRretnxQai04AjhY7UlO/NMGv4MPdOiJMKv70A45WiEu671uYTQcr/8m7zbAnaFDQK
CsMUpc7lbp6sWv2Z/dcP2izot0xlWtnPRkPFthHFiIaDO4C2MzDCj5mvicb9jUlWNigBV6V7Yvov
/yTHKGmFAsN62xPcJq3GAl1x5UBAe29IVk0h+u2xYaaWvAM658S8oli6Zyb9gAxepBvhQo1IvJUn
cHkicQ9jaecuFUwOHzwiCdzoEL3XVOEbDsf1hsDoCWii6niscQh2/nS0/mjmfZ7T5CunR+O/gnSF
luDhoRZssJWi07/FgJIEZamoxmRDlai7BLFlRm/ediofz4BsSb79GMsqrCuDRkhBsad9/k7Rmzu6
YJitHlQRbx/yy/g5l3uaSDfraZe78Qu7QAwHKFMNxvv5qqLnrgmVhBE1dqF9gmtK0tp6s0KJeKVq
fgn7jDeKwc8hLRVJnrgB469fI68imFrpGcWubv6Us+a3snOATlEeGOyJmtV//YTLNBAP7dgt/Tg9
V25mvbgwQxqMBmSk2/cpbJwywq2+ZXxps99/mzzWEL/7GSHzv70u5n22A5R47255mDyzoRLzLyHL
xb071uvsWbrofqTM1xoAGx1CLbZKKirNWPeMXCbVpyOgOvf+YeMH2ycNrPwF/Z7sV1WdvzkM2tY3
+rHz5YRpu2kxT0Se+/lM/ErmvLLPRnwnTlLqiiSJVn0YGJeRciF1h2fe8Y5vR5nxE0v1cSGBtJza
+4OXzwW3IcCa+HrDTbOUMyeWbFBHiNNOi/k5cIPCS+EJ5+xUX+A+cCwZeRixULORoBib0/Nqrsom
Zltf7lfTyEyP8hFV1PKlsFM1NV8lqDP3TcebW7t6rT7QlL69o+457PA3LEDOz9Q4ieMlPubP1NEF
NdIV2QZDRCzzGZkKHfkSe1AFiWBmTuWJwOc+ynuEAe4r/Q2iHUi7FOFXJJXK/Cklcfw8TMlTtFt+
4HdyBnvJoXaoi/+ZZaT1rafFq2U1tlUmyrMOYLwjSvt+LiEUxDgfskjAOgsd5pRj4Sun/aoy17LL
I1OUfad5bFALlGptJqedTiYJXSDbApqV9gVB42ZXqf+sZt+24UrKpTduiA9cGSpuxFha+aBKmGo3
vWudYmaCg8tqKx6o9Nhyco9XMcAJ3ywPtxPlzOo+O7mks+dhnWGWzuZi6pOYHPD7nsruyUCfoAYY
TMRbGsQ+cU1AfouzTcYnGynArBWbYA7RHqFd9jOjgrzbhIzKZpMpd8DO09qfT7unw1atlx/xNbVL
WLiUn5MB8l7hc9rK80oL9IwiHGk+xBTa/lGXG2HV+XHNpNyKsCulHMcqk2LFUFWuchJhISIH//WS
E/kqF0bX8OdElyh8TG6G71DQDsu3X8z/ACMWd9j9ZhHLc81jkRehKOerHb0b/mcFMha5fwXppN8K
q+8m4b1tVfp9Iw1Zu3uxyQ6vCoYIY3TbXE9xBfdG3ZfmY9fF/NJGFsCjywiZ2t1++QuqQ8J191oa
YRDt1FNphx490njtV/bESLXwAUC6TFbDw+mqbkYGJG9+8I3ei3WXl/VtqI4F2COxZ2Wjud69Mhpn
G3TZ27mykDsH+QWyPf9IFVwchsSkcT2tZUo0Y/LvDX4XZ4lea7I42SqcyzDAnCvT+NEavblJ0L61
ICS6q5M6yLF4YzabbIMmxSf7+6CmdNoAPIXUzJFH1dulPsAmJJa/0tSEZw1ddIBhuL6npzvllzZU
8e04de96ZozKlroNjwMdPMqy6gv30e041CdS+ZEJPfCsJtwjrVviQAX8Q7LgguOlXE0aSxR3hbGT
LRHFGzhgSkEQIsoafJiLQABK9jUGsGh7hfQixIZ8Uhtv2WBMAs76tu62OfhC7LtI6qapJ/9UyNR5
Q0+SkxMw7hHZrZn0XxSH/fCqqfWQi3VY6gF2S0xiSGPA8We1QcYhQcNaUyIImFQufI8Hz47ya1Dn
GJLLfekmJu5EhIuxnRWw0ZvB5fMHG9kCfgvhrBgEDfBWkuFdVwK2CfckYBLjTuO1QYxoG+Nn/Jqu
XTgMXF7PtJ1TNSA0ioASyqCdTP1M/cHisCQW+ZDOXLaVwVuylufwZsmHffov+aPbY4NZubhW1kUI
CzEVrzt+sLpcxDR8BkoClYO5IUmRtcm/6AjkG4RBR3aEKP/Sw238Ff+O8DITsAudnKBA57dD3GHk
0ACCnkH3X+reY6XtzmjLi8F/6ThLtDSVZ6GFFWjtDbqgzfPXixr8MmIiXUxPLMatIeoNKh49Dqpg
EuyT6B8bs8ilBkh2eW/iYnb+jTtCqza574S9xIzDdQkI3U9VDatRRQ/+iJXBinmllggZSNS/TyAB
gs1RUie8icUikEIdFwHuhmGkBCync5R4FJeVe5pgrFV5MjC8uqSsfVwuMBD4DR3HBNCQdxS8cfxG
yQTL4o/g0yN5gFeBUXrzCxidRxus9J0xYMy6aEaNH9ybfNpUu1vd8VcF4wReh6k53ZDb8yOWueD6
XwXgymM/qV49+R7CuFS7dRtfzpsM6i8BHGByZ4FQM5Cm7RwQTso3Lt/Xd6rFwxbUfkDJIHh7wqKY
MzgJ8JZhfun8tHdS2CHWySqh9WoWBd32F4yWQ2Vs/MKj+vjeJN0IAfwChpj/BXkCyJtkL+eEXXUn
9iMbzsdTaqBSMxDab/c4c6e8/1KIK2M68D3woWiGCz8AEnvW5j/Ku6ncTD+XcB3gr6Htl6CQXofH
B2G0bqwRD94RwGqFbPoKq7BEOK/lSl/+CYR646Zcf7X5ReEyg39K5VRKHwWhOGlWFqC/S83ZL2Hs
7dio1KDw9nFyLKoNh+TLpkCHE0r4yQ3//GANjpPwInvTj/26TRku2kNQ2Bfxy8BALQHxz/BVGCMS
uK0h+M+4sTVR1i2QYjtzdyNUjm7KuJx6iEUlPmFLbVJzYZfEHrC2DOPI8/ouJHaMCpBGYU2Fn4/c
xqM5f7/BGxOFDSvQn3MqeKolqWHGed0tLpAq0frHtC5xBN0mfTK/Yg7J5G29pQKuhYdbMbmdRe/Z
HkC7ElEGeKgGjh5mLzmcgMc6D96wyRK1ou0FEo2+f4GFBXRafJpoaK8UcdsvhVA/Zi+r48Q4GfrU
BExWj6yf81VipyC8LKc5RU7/EcVDuw9hv4QYag7noC7JQ7+7vr/s8gU3yKvvfFWi96qX95bYdX3j
m6t0nx4bGmDfEtm6E7lCFegWeac/3xoKtDDnxNVkbuITtQ4PmVjEVh64a3bnDxeuwXj0tHObosKl
992ST/vVCBTl5OI621UJ7+0Eb8FiuJjboPA4GCd1ux/p3Mm9XN83hMRllF15Ldm9YFDzy3QSaynK
4HNpkJzNOaJpMwX/T4W5jRFizLvDYf7PcxbIpd9p+TfdJGXHupxXUx2g557prLLvH0Wxt3uMLiLt
PCAYoFjvjlVJiOALHnV2ApyE8jWE/ePik9+NRSaIYBT7ushsh2qhZdJp8PCygg2QTAUukfCL6n0q
7LJ1xp8POIEPncEgAJktNWDNN6F/GQbGa0mtfWoLtK0VadoRxK7RYUf5XmmKmO4q+jKssP+3Cltt
uahtrl8wgkpp4LkuFil6L5FOa+XVHL4vqaQHWMmubDVonwTRI3x/N2u98GU7PHdLYgA8Ch2rNpTh
pDt7jdQ0wlwV1FLuqhIdAEKH2B2L3umxRyuRj9Ex9+saey7g7PX+Q2iuYE6Y1VMSIJfoE88f0VWl
XXffPR041Dw3ItuwQg+W8ne3wkNnQTiM+ph9YjBg7LPQjPe5AbaSkzF4wC32s6kopP5yYghAA7NK
CuD4RS4lIokCt8xos39eoBUG5dMSsQm8OCrEbQVZdHvOAh5i7mha1UApgux+hyR0PiPImGX/ACtA
+AHhIypPX2iRJxQRPPGUKtXiDVmrMtawkYc7a/twOAPtbnOqGgHdIJH48QmsUkimCHVGXsnAZyJA
U6uKGaLoFiAuXvgt465BpqGJm73DklUGGjgNhz7qRyquyaUusENnc9aFA0PdUJP1mTiFVTcwj+CM
heURhBjGzDCJHFsvYAqqBqHX/wezFjnzaBWUYVcD0o8PTrOUWyfte7j8cLM9Ms6SBI2ToSeru8gX
rweCxneVrKbDAO7uQ59NIDzSzjuxyMsaABKNE9GMdrETyqFv2gQ6/S4uN3+hBp4ZX7suTSUf4wlt
K3r9RS2Ax7IGPjMdzMAy8jgC7i+rzlF5ToYUrAohrZAIBz3nkjmIoB9eB+jhxEDpHrz5L1iVsOLX
EqiyArmLZEjBHVu1MdmDnxb2BCZty1CLHVMbSRQahG+33mFTVG6HvtT28IeZZ3RtJ+tSkonn/lpT
OysNZYUzIpjaT2AVK5jLyMOl15dAxtLh6fuCyiYiVrE+1aSwWqvqgwL0D1BYsMdL1KvaifCVcjgx
Sa8LOr27W5s4Qm+3jZzcPZijHhWxKW4XXTr0nqA53O/9W5MoIjjFZXEIEPVxkOM7c3a6I1qu3ng4
7Y68s/JqOkG11sFdsDQmIkASBD7L+fEXR+G92gTTXQ6PKygiu361aF6Fj67w5jtDxnybtM1VGmUN
zIISOwFs5DLkwgbIQ+xCp1k9A+MVyDBfH8s+IHLI6llS0Oz9mysAUXlQGqWTYBOBPpRk75VJ3Pkm
eZdNEQ9HBtn4DpymRsiMKjgpj4cLSXalDYUVUShhKqwqJpjaGPXfmbXdz+TAAJ6BVsoiMOPyWfZ7
eOdydrZFBbhfgLo/HrYFK2/CX55+RO8/sFdIHn+1go/tdvfSP60bY9P1/R6dfZEAOi6QBsPY90O5
rzCB7j9DuNqjPg7e+ZEDMgSLqnCUsQDgbB6Zri9XC7X5XRj+CaKFdneMj7mMaK5JUH3Tw30Dxg14
1AqX+rrx2SNXD7+Ff7ydw6pRsYh/ItcNP6K6vVZMOqrbB8kJc3vb3EQeasfxb6skLODjL4x+i0bb
H4n5AgYOadWhx1k1gcKyJ+5wCcZlG7SlBdKUBUIrCjNW3YLGPcglQMZMlGNGn4M0wM08vlqjM4+g
dOSyiJdHQiCbzTjknzm91XVVMQZhxpi+36sr2634I6iRhVm/bLs6hGDQ+XwADlClH3AO+5K4BJbW
hI37xpil1v8vHBuLqm+1Sf/DiHGR99/JJJGXtC+EIuPKm+HWETiqQ+k9fptekHt4HOfvS9hUuCQF
CMhOMO2DESaXptlrBX6zunn4L3sEunI0xW1z/W2XIbTW2hBjESu3CP1MkzlK3sP9e0Yb5ThxHxnr
LNcI+6GzzGFSU8kskDMK2DnjepraxsPCWDHDuaBk/cPBjmPZlJPuY9flQJq2eZjUSlWLqYsEnX81
nfBKbjlzHUJm2GcSc4Q7LbWcYPWpWByC7VcNW+DFuX7tI4U6+14eD0mP8CVtlb4x3D+cD0vL4LDa
ydgNUzgdxdsPnqFRHNbHRGlZ0dpIk9G72/+zCT8e8UMZbfrO+MjzUDcDtYhNth/eAnB2tsWH3fe4
7a8iLx6XD3tGfp711Bt6oriDQhDL+1Ij1/hMkiM1Tx86oc+8B72wreRBaHQuyTUeMQTcydI4UUI7
iXSJTidQuNsOcZ/SjEYOPSlH0GAhlpLR1JfvlHa9QUeLv1YGtHpuvHkNZDXLmkRlPYB283RSvMSO
XjHHn/poMdG9nu6mZijupBDvGKpOeybGPWGllMsbHt9Hb/vWT7V3ujQ9mhyV0NsG15bn0NjF6PTH
1pEeItlpyo5L1rIP1WtY3H1IdxtJfWsh5+TizS6vKowROqKhsMDcEXxOzqi63EQUpDO36w9LEYcI
VWwrnoJxozhUq+rRg/WtIMoKHTCEQSMSMR5wbF7Yhy4u8zebrN2Z2Oe34kjpQZcn/0u6NGEaUS1v
mfybc7pBXgrS3vdI8riTSN0Gf/TjtQ7iSZ38lM7g2dQMZwv7nd7hrj4UElU3WH374unVl5ABrCNd
g+G8LwJlNBOtX5otiM92/uMdLIPKGgME/P0Vlsf748AKuGcoemNGVhYZL3qZUlku29zm6RpDVd6P
BXUSof0Z9b0ymclPlBiszMY7pPDHkzEbubhn7Gx6VTuCqH8dyPRhB1dwIYq84fgYHh3KR3OJ6e1/
cXG11HH3Nry+w+Ykdyn2cxcXL/dDfC7AEU63SrjeiHFtSbTXxBnT7zZcPzzXd6JSWbaT6e0IkldZ
ydRa0XxNgY/S4M92B0PkBkW3tYFlZAGziod5S0u1ePnLvCDa8rWoNo52iaRtU8Xj/1mW0b6kXr7Z
yA05XLfChCqAIrRaH71yKmqABUDP7vKtGjTYdNVfVbI9L4H5cvEPYEOd2yXC1wkS8x6c5wg3MZRB
fh3sgSFQCclIRLYdZpRbYLHjVW3S2vjjoEVWXG6m5ZE2Rwr9MV+NqmdbGcFPVldy4mg3+R4Yym4j
JrP4upnJd85+G+B4K+1/AEzPeSezMMYM0EGo7rc0gMY+YoJVXJLxDmjtyFBw+zZaiRgf48KuKcM+
LcvWJnVf3jN/cNVB4v3HR3w5R4RQ5o4OP/vzYy8s8xPWhrEOFkEFNsEuJt5UgOLQcy3L+pbVuM1g
h095vihJbbRKqEnKIpUEhMkRGkXBBM9An0TpYz+GN9GqCAkiRN8NvlSwBD8XmB+WhaEmVXRzFciw
yZ+OacRSONBU4396JZi+e7ch30nysWvNUmNL5sYLkYiXCu7VNSxNFcYutqsRsQZMegQo6Fr28437
iy7jEdHOFvtZPVwMHoVNF9bfp+zeTUpjutABJZJNxT7DK12VCga6B5BoMeqhv2SxWNie7AjMEWLB
0cVMaLbA0q0WhoZ583snKNHR6ldyKYe7CSKrFakVNAqYeEq1fVEMS/gejh2uu8kOBdhob6OzlmD5
s7SvKoEnQvRNZXxtvdBX9k8VqLMfluaD2Ak1T9czdtoDStzKt2o68PxdZJQPU0OcDNDxbvD0Jeth
AzZsTw7wJq8ew7lFc+3k3HCM4VL9rqnu3C90LhrG5sQulQCZF9FPW1XKZcF2uzXYctKYFjvGI2xY
77DbUV0NWkL4N+KPPdA1/Rth1UacFw9CT+Lc4ob36wK2pwcSz4FFOmwShV1TvukJURUucn39ZYDi
B5wTHazfNgfhf/HDKhCzpIUR602kmxs4BOAw/WVS5/Ke6HEa/vc+vSrgUNpkVSz/AM28uZlaoXIv
hu9fzM7cBXXQvmmg2rRNgaVbvP0SvZ9rex0yoaFoqwW136h1A4SkBlGF2AkO+YipNyMTBHvpyy+g
zrvaY7EFBw3N4Juu3HvGp6HQOJTNXN9Mk35ggbv48/nwa4MR+QdSMaI+qsN0kpV+k+wYiXTx3alt
wR1JvdHL/573A+OO1lGgqU+Ko6da65NxatJr4STdqd4BYhF3pb6XPCZXA+wDOzho1qbnw/H94AGp
XoCgCyrZYEel4Mgv2r5Kc9lPB0u8WDi6gbgzkDg8fV9vnC3DpLQbteBDknIbvQqAvvjfuuHs6sCr
Nursu3ETl0hPE4dYjZipYxYrypJ01YZK4H6KltLUo+Uz7X21rBJBHZ8cXJlHj4JZtMfAqDcxSjiM
I9uA3JmFhdww2qw+7i0+Qj/+l6ycxqrHPYzOY1lcoZOMfiIPdScW2ycQ+h6ru+0hmahvtykrUFS2
Zw5HqVmAv1HCx5O5qob4M7Qw3Xb0GsrLM//pjA2JyPEhLTrRhEb8lp8nBbfKvQlnbJEQo1lqudrM
LYEYqPfkaylgNebvxtgCJVcbwp1F0aFHWmBRwlA2ZJHGbfuLpXzFMmO7JHIuQVhDKoqscEKjRDsx
SFERu78xnfKGTjO5/IFFbHWe5qA1IUffcMMBPc1+Iq35gieyuJEeF4f5f3VSncXfi2MoXV9CNA80
ZlLXctHfndL2yBr00Kn9x2+zk/ti6wIASlzGX+mLYt/fMUax6YV6pw6bk5+7Tm/KEGfkY8FXJdbT
a/59fdmyLobQRFnxJkJuK83pmgC2xsFMB7oUdPVgFAXH5cCaLPzo5PhQq0/eRBwxsD+lEqXCYEhG
80tOBO0zUiVAB5UARB0iaU7emS9uRwTLb+j5oFYW7JXEnkwzUWf6Zjbvta/fQMck8CqYaJ4a3xAm
frHvtS1gjcYLwfFgqz/e4JnX4H1hyZ/kIXFCP1HK7v+bS9Ei77kzs99TXU9b7W0b8s4SCqXxRl7Q
+o9AkBHEivcKR7DvJ0Q4ma631GYtMzkEfiMGJZlxxdrM4iiVlGdSQTHMDNMpiLskqpm/G5D3RUL9
FK2Mtuvd9bzXOnTMRwIYrTrNNXPn6RlAcXStL4rKB2r9K0S3jLZcpCjxowyGOfpywqjhLSURUlCT
j9zw0I5H4emtatxQ++O7Bn19WNvNJa79/hZF6ndywb61k8AmZ8ek7xALPMnxxBo418mtbvWdIcIN
6pJwU76W19F9uD1Q2j/R3b3ahJEIs0YguAkBnqwBi5ebQ6tULX8mQZ9uuXTPcaoaEM36JWA5h0Yn
72QKlVAOhxXYxmkl9EkYH+pj5gHipbf5TaQniKMQzMz12r9PU5ebTZRiddV0qLOwrLv4BkN/RET1
LBTcFdFieaBegG7VsqkG0PNfgaA+bT5MZllzN1P+QdkuTsE+3fm7WWvqlasSOhwr42Y1yEjtUthj
lTZrv4QrQUu5UvmCt2hEZtrSN4KQm0ydXK03TOjO3Avs4ou9IP9UWDr2xirepPNyLKDhXqB6ZtnG
WfjOYF8oIXTmpDdzcrf6E3tLxcvls+zSqcH20qTNHpQS97lIhaO2gDfYoZUxbu/VEMO/u0PqFoxC
2zi8xFT1Vt7VzEdKre26mn1FoUo/mk6k5PVVogG0gurs7LlqorRNkmUqrbcYyDV+UT2rc5KO8OJj
SsBn/DMtCMakzS29M0pvbaRka3QcoMZh72jlScc0BSvQ4lvIdJKKZpD8gtE6QhJGqH79hI2ZbtnK
lMULdRs5F4VbFDdIgH8WtScQwEvQQaJK9xZfO557keYRvXoizyvuR1MycyrrFCDZBpG2t4W4Jygb
BrDVLLNhS0uXgYdiS/ztfo3B5N85MfuGeVC0cfb0I4+qsi7U33p3j1hWjUrlf77Oi+bN0msfTxgb
YLTlNJC6L2r2qLSV9sHfmonRbko1sQbViIKdSfmrlXFc3UN9OKQA5oaVsaBFFw8DzkHNH5iQ4Oil
tx2jQo53hqipTsp8dMCrAQ/HuJYCYrBl7gowZQkFyxtkTLZy+TGfoJoex9GWEKia1kaxQ+0IVJC4
6keVTOk4QR/hDGGG2t0lsJnezlEtAQD+K8M5vYFVs6dyl4PUHpJm4SDK2bJdL/0+We92GRHhliqr
i4TPsS+kVIZD+Bs5RJxFiGwodfrUi8YlKfllRI9KBqydIbiZ/mCrRIJ/b6uTiCxdAi1kKUV0d76U
BEuuOeehuNHE9MwD9JB82QaAt3WbDkadT9jODgGSf6KWzNuwQDd/TCmbdl3s9hMWjVxQuTjUQLxx
0XJBCA9jSSekmYJaT7lRogmUU5Hv2jS733Ocdy9VkoNQSxgndxoGR40Z0tuqTho3oZ6z7/boGL8C
zoVmT4PRiTYUJyWJEsyAprxTtmda5jhAEnQYbzw1UqKwnmP824lGa+EL0mgShRM8IaIgwyay3LQ2
kPkXkM2Pli4jJWXjWu8b9MJATfk3znps//CudjFJtU5zxVCmXdmSuA4gPkLZHH0Zi2uDt+VkV/wK
QGJ7UPrWoz0zu5g7gNRaRC59xKct8hlF8/7KYJRGAI5U1b3bsh2mHHl67kJAHgJclsui92R2GPIa
ALWBm9msDjfHA1FOHdcP8081cyzkTXQ0dCWLcSZhhfqx8fasCLS++4qIz1L4dkCAoqqqQgFFX5Lx
onkLX4cq+qJJwDg13AEIbMuQc0V8VfqNlkOZFtANUrfre1t20oqYT+8F2pwli6OHyQudvCXIFAsw
ysR8ypeAUblTJAEBWSA0c7L9pXl9IeA1lQLB/9o8YvPbTEvm21+u8Y9KAEkOnk19XSE2n1/Ft/Qq
WngkglMHcu67qijs9reK8P8B55J7scSxSSplCM34KoylxI3PbyM2jPsZNeJmYkGq6XR5jJgtB5wt
wH+8wOVVD0ZR2Vtl7vfdO437yup/v0eTJfyFdM14hPK33qwLQ8EiZWazIcuQCGMYHpYCaey8WBGe
vJEGXjY1yXso9j7OldUqpggDV8mHiPzMyDU5k5LSqX6E/AxwVz2kGC0DC6ar6z7Mn2/yfu3/ACTS
iFCTZR6dgyYEWV8Ty+JlpMTqpVAAfuiYuv2rRiAWWhuYUuhJucSA+8PD2Svhbs/xlCYbfQ8yIuwe
R34neFSv+YJRrmsdkbZc77I19m80WUprBIGHpcWNde1WJz0M45AjAHEeYjiqeZcuMmR2ebJRO5IQ
uj+RE3EcPz83hWeHvlsDGADHfQAMaZgN60Vmdrwf+ApYLm4p4hkSBYBXerDItkUx1OgNh3ULJFe6
Z9MA4VDK3+FcQ3xeFZEbgrbXX47QHRqWRffHHVvGtlMKCsDq6qPl09astPPZOjOeo4Z6kR4o53WL
iBQAYAvazpQEc4h65IupdIrB8pZH484biQh4zbZGnQeK6MjU6CCrYMweL55DTLeGkJNna/UC4a5v
00K//hFLaByUZVulnnEJe9zEYx7IYStyQbrSgfisqRBg/tj4nd+GVYbzNSALwpOwKCV+eKD3xdTw
bJ2kug207ambhxA1P25jODzz7PxA0TxedIohmRokMUm/JUdvqTXL1ViEADN1vhhJo12sgetEtBzA
OCFDz3zvRPS8RtGdDGe9cOv9s75aaPkVgztmEwBSxmQSCnU3tuw1u4Zg89wlycJRhhx1pb/gaJ7X
Ty0rzrrGez9xxt9RXID3b/LpXo933ragrE4KlEcfu0NZo+1ChGdPzbLb9zGMABwTSwFhUP0/03Dt
UeqTyReKnarKl8G4tWMqMC5G9ciIVW2/GSQ+Qz5HA6hdJayXniGxiG4d7bBxSuYJ4BsfyqSeV2FQ
xFdSSeJZbfxnhzp3qvuCOUYOt4vl9FZhmYAoOT0y0PaabL1UGHGE3gpUmeCQgmwc8S9yiVcQKF/I
kllFc4Rqr2i11t0Ep43PXCTavNOp36zhvxDdpY5aOnGezqLkXGlM9cDyPyeScG+3p9swiieONhFf
4q6kUc62+KafB1siXXHvQpU4T8VnjSkFNqpCJdoayEeo1p2NNOH9SMd3uxZ9i/rS3hh6T2ZeymeT
jPYzhgMaciNFpc8yRNy3Faov2QF60Evrdoytyl+uaTTjpmbICfP914JTEcGyjxgVxy1RVskvYTtC
ktEQOGi2t6I+Y5cqa9IgusLOAKdfkDTW2tYWaWlPiOtDU+HF379CLYp5NSM4/h1zV+UysvHJtI7o
tK5kSU1CECuXh7GerFeYbaIzw/Hlixr4b+xr2QslfOJgcjruOYX929fFj80eF0S8jJqZ/2gWnUZl
t7vzHRzLSU4gy/KylRu6jZeWJOolMIAPwtX5BnceIA6Zc/Yu0bOj4Wk/65OWVxBoners2FjBWHQA
FAgAz5b5flUGeIJpNK9YfWtXg8/lyY/pINXpHABgTVFvoTkIJ7jmjxp7pItQk3+G6C43MzXeeek0
RQPhPYfNug0J3N0bOTgJeXdUuGV4gdwASPHCCxFHdNoUSR6q9Rd1Kn8IHkheLAS6jXQyORbr6CNx
dW7/Z1XXiMLgh6nJTKd8YEku0I2PXv63HQEynqhHnJsXc9k1abr7398at7LtuB5ggz3ssE/b+bWh
CEMadOr1qaBeEwmHd1rNXZEt+v+O/BWx2Ekt+Npqh/A+M6O2/O2MYdBI6RSCniXyDv8WuYc5Gnt2
wnFPqZVuf2Fd+hnF9Mb7T6eJZvRu1/cqhnFAZ6KyHGD40C3rjRySNxsGd8TwmYHBmiF/62/x5qny
xoTeIUR6zJ4v9A5WQ9aH6Rh7E0jMxRrwwRAHoBkqIbg5d9ZEmhqBB4BddVtv9XJcDS3sfJgstICb
LQeqQg9xc7s4NVSoaUGxHvXUQZ+pRQlosDCh44SxrF3kfQJQRcuNWjtEzavCvYtdTXYBO9cLdnge
fbOZv+xb4QYJa9usmMGzhiAvSx/dKiXraKv/IQxbExxxKG7EfrIsZrUGQlyRcwFy84PPxoIPkesB
TWhClKIT1zCQ0n0qrY1L7KaytwMJZ7UH3Mn7YeGNIYC4Q90b/Js2QkQCP26mrS6rJ4eEcXl8IS2J
FKxeRq8d9skqboe6m9ZAmLqkNwElFGGZ0VjFrxe0Wx9MCG5l5K9dymIwnvvupGOv8SnMUvexFo7k
pFbfQ1wpeLtPCeuG//Bz6TXSNHxVTsygT7Cay3Tsc3CaD511+aMPli3RR4RhZeJ70d7peZf0EUP8
UO3epqBr5xUW0ghbwJfs8CUKr3fQnmEJeDFs8s6/g09PzQFA0mtysXbomsm+FzlrQE53BwOpzvlY
oJS/IpcgTTwO8+XQFvcsKxObE+4Bq5cAGd/krsGpo7isuqUUo/vHM6VYZz/SLrnX1H7+BigtNKAf
WSR5jXuaccb3zZpL8friIoVU/NhOhienMLmeDmquJ9WsHKw+cj++PNUctrbN7hEfIyFd8ZXPezso
6+mJ778nZk0wWi7zxK3g1QryU1O6szCq642s+tZFiTqN6tLXuUOMvz3rJTXjXkvPihpgO5iui0X1
SXdVXgX6uZQV7IyFbvk815UtbXWsTFPMlK5JCyRPTLBSxa7Nh2a0xrCMXXMrpMBFCnb8rQ3874Cg
LknEYRq6WSm65RyfrdBL5+WUnXtnPi8Hyut/v3gR7p0Av/8Rp5lo+YDMw70mgpB+oyeWb9OVnMhp
bEOlGpWBVqxCKgBPzOZHNofHhksz5XKt4G5WWAxDf6X8aVQ1YE/b2tAp2atwgO5HRPO7UsX00i+2
ITeNG1bZDMSOg+FdebNfmIotpvmp14rtJkvvTlNeSJsJcdQEjovuDBWUhSxE6bV7tPAXGqcOwWKr
uXJWCS7ps1rA6bOTA70bX+5hLoYmPbN3qTdQLoKDOgYxg8jHcUh0pTgh7XYAOXoZjFdvG/oGOEeS
7jfnwNK9doYE1JIvs7lCIAsOfiqlCho2w+g0hedRUNcm2TIgL/Ki9QONeUYn/IRTPUPJYZEmqTbM
rm4y41AIKqBw2p6b3FVHs+1nVNoVukcIsonkJP2R1wjD1V3MViht0fqd+3Tyhu80TvWBOXGqHTIl
LvZXfvSp5n7c+850v17vSYtlJep46gPYnNmf47clEZrfNspjaT6A6EbxDrX3/v8Iia1C/xyzEH0Y
Q1BJUd44jhNkd5lQihhTjPcGbuGVRf2PTi7UuF8aGNe/1jUtrgtUqsQ58KhedXeuM5qbo49nE/cC
zuvYZV14oNPL+w6Rcr7L5EHRYXtCqKex8fwWJOmy+X/aDr9Y1YDcz/dBx66gg7MNekTbV8jxC4Ts
d33VmPnxxxm0oI9xBCXF9GoedTcF2qQaz6BxRSXXWZwaP/huTLDuk46WHEiSyameTfLcUU8pIqXW
iHuls924V6tx5VzGL8AMhcKsD2gVaUKK8jVUqdOZlGoglWqwDEh6uIyx+4wVaRjVnxP3cvPH20wk
+hHAMN7LZdnWusQfnSQgBeJ1y4pftYvIsMV2N1DumUzX/lmlSpnSFs5iq0iFcMq6Il/WK6dHOg0w
8qGrFgqhe5topToTsnFyREU531b9rQTldnc9c776NxJKuWLU0L30l4DUDGdiax9J+c6csRzTL0nD
ox2hBtDQ23QL7tATFumeeepEgYEmsXzNc1gBVC/ie+vZyzNcsC6mG27dj6ncylsjaAo8AzdW3gcb
Uhb7og+FsEed1J40thMAKlHWfY7mvpTQJJ8cEXUf5J7Uubt7Pg0U3sgEctWPsvU5K1Qyq86G+w3U
mRN1h9x3P0cvl46dxhgEmnYBJWXrkgMzMOLj2FjK3BV/XWqQ+EFQ05qjWNfEcgwz0wrrcuMrWGNM
bHHRWXkXHkn2I9SF7tYSTmBEEIiBWslQdH9miuTvz68e/RMABlYCoRfPA+/nOgMLlwTXI1ko/f93
UYb3eE2ZJ+SVCLltYqTVgLQCrU4P1gLzvQED8C+EMaz7FGUyQAn5awOhGlBU//Uvcq7XrUAjq8PI
St2knevoh7pJqgk+FVVPdfnNehVY8DxZdQVm48+vsv6eN0slUX8tQ0KEYBxXlz4n6dWT+O2rRQ7I
6kzPSDoxLyA+I3jNoVr/2F33WKVvfNp4emaG82mmz8yLQLjQng6gLm0/hMyqm5e1Z2R91rX6FCLM
A/lG+rOY8giKUURlzM0crXdWIZxE9A94P9WKf4zkikQ8ETujeRt+3mBjv5twGUWWuz+tUz1VVQWm
X42M28A3Hve1lB/3hkKnCqvh7XvGPSdWbeLxV8NpMwCHLzKCPiCpFr+Xs8s0m5wuwjxjJlx3022n
ibcS3noiz5+a9V29AYhEkRhX8UJPbmCy63n979eZg1DhtbqUmkGEOfzJZ3WgXJ70VrG3evrC/Axe
L/QZN3F44mDeUE3fcTLfegQkypfDhGxVPjyFAt6F7FkRx3t/E5uJE0NO9QQowXX3XvW0jy3DLV/Y
xUTizE62Fa/dKRHL9+xk+sROdmZ6v0qpQJ2VRZ/qY0gCzYCBgCmAD0u8iPyNZb2uochxIVfjkpIw
CvtEuvuPGUxccgaAmj7kj50fZQvG58z4F14kfJRGrx5uglS0Xc1isGvL7I/3YnCOWDymCLmj5gV7
T7cKdwdldg9LzzcnHWDUdUxrb+UabzXZB9GbqsrJtQ12klRmUWB0ImMAzJZXTl3pKlZK8OJYe505
l58G5t907u6s7Drxf82jTsZf42NnoA1EDh07APQZytHMUmcYEyAJpxyFnUu3DhA82SbHzQcKb/Ga
5kq2/h1nN4Tp8j23mXxIFNrX8MldPNUobkyeaC6jWcp66oFZn832RFQ17DwgwXaOLU2lq8dU5g1K
jzcaEI/KxlexrSv3VQZRX4lWRGM/jxMtibvCqC0secq8yWzURJb0YKzGckFOLtyyOfwR4NQibrOY
ohtB7Io6AfpMg5Yvxz/oaBmG9HeQIiClqZWd53teTP/nYt7wZ5Hr0BQEq8JZ/9+69R3hO++EAsn2
1c+KK2DFu+RYG45VSMmJVBsCaiIH/rpDXWRO2v3FVsP7P9Fkp8vi7YfKdczqs1RgO7PgVbFLkLwv
OHl++PlQbDJ+4srS2tcISqTmWNjz1+HxbU3wAOP58haeLWtheuKG27psuiBiRypKNEg7QzAG2pLX
lNyr5m8TjnvmwiUrBv425zW05rH2utIef3OAUYzo+84h+COJR6uKNwzz4zaqIfyHl4aQQiYpZ8Mx
Pvk8oDOf17ngOq78mveoXHBqSo7t30mm75g0evjKwc9E6TXZZaDXdaYAOLruwJTedUO3clswbVMT
wAlhaz+M6Ph7zsSeiuBgLHDnZmScDQ5jZPTB1Imw3+6kWsa55C05yeWUT6a3LEhvZ6qESOxQxvhT
cLZa4t+0NR0GEdb9Sj50fOiC+HNwaBR0AteJIvEgVtYpD9CWa/FOfshqpMrF9g/kVfTQvdZEZH0O
ESmRzutRJpY8UaqNwFfBFKDTbNwtvZilBKXtGxEgTSskMWAKv7iWvxGGhuUrA5fkcOAsrCuoV/1u
P/nmMulnaNP79pE5H7IKWXpOvMR10K6zdQFk6Z9Q1ffOnjXWE6L0zfSI+KR3+yr8leK9HpT3lqH2
pymxUHjtHOsIa/9m9abrpVR9S+jM3QxXnJ6RRF5BXVrJJGLRoj0zlW93y0BXMsJ54qivY5FQtxHx
Mu9jEd+lQUrcLFtHfbYvDv1jLYuXDQL1+HivotnFrCOxybnRf9X/r4ZEjW0XLe43uZfS7ZIB7rG3
jBs591Xz+57fERV3/5+U24bzAJq6GBXIGYwKhISOJujCszC8v06yT0dk0UEvJk5sc5DGt09tZSK5
pJLKbSG7zAD1ziYo1LWc4NBv9y2amaYvjhgHDfVSuN7KdTiMhXHpnLMM3P3+EzQpl0hdzQFEoN2r
QB8+i2l1etMrlm6486bMEV7LTuXq1Uy0LY3AONHSUlEsR++CwLuGuPOdYpZMThfwlq5bp++FWYPu
4qzjCrk8ubbyb8CJaGC6tZBHHijXuUzqiR+Rj3P/+NvJ57MX33d6S4e6icrNnqBpHuS0Hnpol6vD
2WTIlOtYkUeLkdWxD8E4zpBL745e1ZHSKjUnN7iC7oTNEjakONVLW5H3zMsJS0/4Hyl3G9v4wlMj
zVxTpAxe5aEovfPpjVyPzhXPaW+nYSEI1o1RsSfhji2HgKAEtVsJoLAI/mWKVW50fPCzIV09evCy
YgTGMDSCToCgsuHaDpyTzvvO3V+0kYQjncIrkgScgAxLP1D2S2tyNM4bzb641CEyM9xbI6NKLPQ2
VaKmEgjj6OKhRbwCrCtCe+dJsKU+NInLGdad5ZoRmwdui9N3vDFyW7psGs2bdF4CSDSWt2/HByep
eVYyyMwPDTMxd4X87f9VBmvBjM5WxjtA3H7fRE71HyKXLnL40OVVVLVQGIHSkGZEBn7P6pYf11W7
IjzYCJB7tc0+izLlUZVKSIEueSqXynlpEEBkDzmPfWaggh/nPVEhvXxwaL4PvaGAmv9ndX2ij7jL
8ON5QoHNMxczGM5SvJAAyHMk8Jau3txleWNZn19JD5+l4npbcoLbC0egCDoiMOtEBNtRz+Cl7wXS
iE/gcxb8mfFnZnzpdkjCTFoSiWJb39aJ0LvD8cPkGF+Z6i94+KuNc7pTVsnGf6rKGple7PKbVgRQ
3SS6XoKL+P1UMQNdG5JKvOgnS9tGDbYX24jmdsX7aH//UhEt3+98G5bA1QwCHDZ4WWYm98NxDGo9
+yckN+hH4/lTwnpf/U7eOymqzaurd+e069LpXmrleKT2tOeQN4ImeZgJzVbDwKTnc84UtIDZb6rW
+oGyIIB5LnXi9GVcKM0i/hpoxMhj2EQqqUGNkBo0+532oAk0H45rFTqSs1h7XyngvqT6GN4SlqDX
C0STLXcbuOvimorQv3xSTNPeztf6gZ6ovz/x4YWcG4rAYDptHWTD/6J6hss7KrlUWk08E3eW8vZc
irt025j8+ulKr2ItFT0EM4unTMz69icClWlEUWHms/c9sjxF/6CeYO5xqxzs8bmNvzKaGEqinlU3
mnV3krRCGTL/RqysTN4GiLfvV/zn2/6SLjZQKe5aTKvCiy3vrAfWdIS/iB4iRUW3sXyYg7X0yPKE
fdEAOZ6u8OhlxHgMUNCwYORbG56VxilWn/Che6jswwc1VXdVLiahoA2FiDL+7Jbf0kSgcqyMyR1s
EM1Oq2R3tmqSLj5+/SP9yYAf+hRc65hLgAANimui6VOxY8Ubb1+bWUtt8X9cXAZHPd0WFi/CJTVY
LRhsCru8o6QTT9whel+6T++1utmrmdKBa5l1m/IQf3buPmOu8hhYRWjIhEZR/YIid5Cu5tykkuwy
twvZhBjgEFbcoFRVgwcz3REM8FH8yAN5LzfSnwSLzURx+7ClfVD5CuPZ+5drTrpciWDKD38Im41r
pd+mOujERKpEXlfl8CtHZm0FhOHJtCgmMI8cRad2dxaW27iexsykLr+TT6B7w8Gx0bXP8vQ9mYyc
iaMXFIoZ51uHO9nXOGqXXdRCSYJ1lXbgeYpfm4QhEKEma/YO0g3tr2eujN7PEFwtcEUt3+b9qPVC
AQGBuw8pOH4Ask4S+NYLnr4Ha7xURxWg7IH8K8m0dOm6t4zjTpjfiMUzw94mYoVqlEg3zSLhBaMT
+nl2G0hwYDQ2Kmtjor4HwTXe/Qo2ZuCjX1knqtHJjhlZSLqPDLfhJDNEvRf+pygJNpNpagB5dxC3
/xmn7VNwG+wq0lyU7g2bWdgPm9vchnXEuz+EJZ4C+yqJBO+5TF5vputOXtHQ7ZGgwYxlr9tzydm5
noNpjHDjYd/nUV6fdIrwKMp/q3vHR0MqbFCTq0j7uu5uLomlQqDiCZy/EJoH7lJcY+Lg+QTcaUBO
g6z/tzfyJJbY/p7gLVi46/4n4FQRncShJOhJxZsEbT8HUmkdd7/EAXr5X6Gpe+yp2Rq+Fk2wWqH0
DUnpfsCfyHbJglL4l2EESz8c79KR4bxX+Fz2slvflqA8AspBo2VCRpKCYnPbJ1Tjlaf86+ed04UB
VnLjK8PZaOfUurA7LCE9UPtjKds46yHARFi+jUAutMeIX2FIaOqjoYsGEK93YnxAuk57huwlL08p
amyK9r0Grswd6dr47B48jVbScDBz7nAuwSo9i68R45IeB48CdzaOA+ZMITfK8kPHEfIwAu+4oNq1
yO5ECwvO9IfYFytliH7e+6SwRA3sZyg0l3UGlZZ159ae3kFVV2LEQn3Ur3tydoBeXm2SpXhFUA3t
/LbovW5AxsXPtnyeZSi6eeqErhboCYXfw138LKQfA02zae2FMZ6uXa6etyWzXi3rUpnbRVmK9+Yx
68giQL3QArmS5zKqqhOrO3EMZa1vNSzjvC0pCB+wdISiR1uqTQS36y3/9Q9eSqBbTfJZ5fHy8Pg4
LVI36sqdWmC4HSSapDpy8bypaBE5DlvpXwZGenVU/WgQWzbrony4DL5XIgI267LZqXlb+1VzPENn
IPqLqclh/kSmX+EyIcgJdanGY0/dkVhAGeBBc8G/p1k1rYX2GVJi+mEL0DldPsdTiZTDK4yv4wqf
sUFNDztefH38ho7WTk0meyue9a/VvAQ4169S7cKPXX1Tl+OrF/sdwrcRiS1ll3OuUIzmD/LC8y1A
IQXXGi2F1OIUYGRxH0REdFAf6gcYjs09hgiP7D/1u2JJ9EiqAk8DivIkHjI36c7PQwshoguFkb5L
AW9eLLphH8VEVBY157L9O8WOstiBlNTxeXRIadL4T5sdkMN2IcRa9/GsI2sXA8+NwgNJadrXnXQz
pfqfj4k70kb+9MoMMsJZQgLPfrTkY6keX/+lw+dsoveRELyyVN8vjBFNZ7e/dCD9ioHTRfbBMC3X
1xXverxpYAsyXlt9IXwWDf6V3RU7ID5PYf/Qn1ItxixosfNwQlLig/OvFqiv18MwB5jozBQZ97h4
RRMmlCYkn1smOMxm0NT0qSyEsd2+bR6vwTER7jCQ8EjyE0BTXDq+W324kBMNXJCEgSvUtYB8+sE6
BybOgFtxP3Mbk0ZVMB2eNv1HyZuPGnUye1QS6X2Cm5iuD0iMprdS6jiglYi0yhIWHUphRkOqf6LJ
T611zwSyW8ZaHPjmwBway2GFYvcuLmH7uVCaMfsU6+bgPxongT9FYNnYI53dh568e0YAa0tSIKMU
N5g/S280C6o+Wf1e13vb/IYJAjkLe6nsz/l33/XlJTO/h4HNc7rDWZLi+GLQxtlEHrsugn4G5Msp
BvjrPl6pZ4joWL7t6N6kEQAJNRmrzvf/POdfJGP7shoyx8dEjP7nFdZDoZgz5LTPrJU7McD/wnY2
D6Rur1MIgBn84UNYxYt++/lruKGr/wRF2pJxWrnYHQGU0MelkAvx3LqnRpXB7MY3rob9mnNr7n9H
uP/5HMUAUt6fiqxar2jnGqlGatnmP0e6F1A+Z0kkgNxQc5Oe+XZo82XwJ+hHmMdh0OBdVOCBSsXY
KYb7lEkYtTfxhKydFoBqquSBck73ylUhHkLyvGcbkuyyvhCWXovVurf80E30XipAL/rRhtuXIVdE
B83wAuH/rDZRXd6lzaUZPF+7yaNTatQOmLMh93GV6cZ9M895iRh6TSikMLic0tor/ZjHStq09xTx
bNZhjnLDwlbbx8tUiyNreI9odsgaUwgH26YvWmfwgSVaTCatNnWqrbFzddAFhs62B4CFIZCQ71ah
iYn7Y7AeY3KWsemRUY06AXfDLwnxZWNWhE5W4AGP61QsOwTF0/JCBXyHXzBONhHU8YJqx+HYJjop
9pbdGaHdrsAt7M+Q9zQTZuUgzVCepgttg9KxfbWgtcWPRqHo+Bju7O7EiaBIJ6Jc4sftVrN234R5
AXSbhdiqPgHmsznhQKHRHYgGmdmDt1hvZfP4wrYJN6vwZORxmxuf+SFLmX77OXJOcjM3NBd6B02d
K1xByE27DDXpCudjnl4H4j8Dm5ypYQpIuwtOFbDspF3bAoxVKNwLH8w46wAn6N44He1sWny2nT2B
I9xSrNRarK1zqUqxjDrcMdgQTLOMI1AMoFNUcXU/RkWjozfrJQwboNBuWWplwhOt3bTRpemD9GDr
t9NdAUU1GrFtkvH8bbsoAXfmkvTL3dwn5NuJNYoleXQOoiINHQfq3EvVBGzc0Gd3wEr7sROnGzeF
TV6UsgRX3sg2LbLYwhi+A+Vk7nrxqkAoUo5qxI15O0zKWxvKaix9XLtxwDEhbBCU06Y89q+kXgGF
+y5RhtmBMWPa6/zDVi1obHWUerGUrZByc1u/79iuTiJopKsVdSo5+5a+WR5SYF8LjxbJV0njBeci
d5rhLiVB/HW43jO2hYXM+95WjbsFxRHEW0DCvl3Ce5q12AF5TeigUQvIzNJTwJlEZSXsXfAK+CNr
goLiNT5ee9qASbw+dOrY3Udncsi9C1iQW+4A6wnirwaX4I9F574EfRH0aK4J+KI/aI/bJHv523A7
9HPKUe4ImI7NVvMcXoOcIxsaFmc5xIIJJUTvykCfVf4s/irEzpuJKO6oxtock9dG6W/mizqlCcLw
h+gaV2Lih9pzTEV0CRqSPb4h3lwL8Y/JXiselZIUO2zKkmNSx/Ee5sbs+uPT+HtsWGImqieWZH5V
VNqLlvnePS4oQNpq/z/zI9DEQTaYphwAb5aUA0uydK5lyUjIe7yyBunyhYX7FSFXtH2FVrrIcvtq
1ZqZEEETvv9ef9XQgwGOBjgcHEwvPgjs/TMyg4s70LFOBXtXOl+eS4r8IeHeUD3dEW5rPnkR8BMp
4Gl4XqLTbI5SLFm0VjADhZdtwOjZr6G+47ESJgB/25wAtX/q3OXroD320k+8j3iEcPXE/mqG1nWf
SKUKuN/XscENqcGEHWT58waF8z/duZpshAj99UXQWxCwok7AtoZWvq7c3ojeZFl9lsuQz6HmINuY
guBX/+xM23T1o78VJkFXDEjVSZ0U4/Rfv/eTH9lva5pTcrAzzbTJJpnkQ1Vy1mOIO4qFuUEhmZ47
2FxVVdu/jdLb2PugDg3I+SFaUoeVMqqoUrjtJTNuklhtJHIeX6eVN4W5X6sWPSRx52lCNkAJhs7T
Cv0e1Ldj7TQybRBTMO1pNTcMDmlKr7BxFH2TVG7lJ+QNP8ZppXqRnuTV3GqUSfxpeU9uGfIipiiI
36ZjZLy1pKqVE6I7AdMpps5xWZS4ZjIjdpPmCzaTAQxrtvC+fapvQXJT9RZb4DTbvjxiAhdKQaM6
TZnACX1WkKP/xmBMyWBMFNtjENWRKCt1iI+YKgb4Xce+0QY6anvMtv2dlZM8auY2pJWrbrdYL53Z
6etaSFYODtz2zmXBXYNo4e9Rv7SdyhJan3tBLRsPq3hbqAkWeRjA6XtFfRbb7ezEXx7pTDoE1+NN
B0gl+HuQuJoeoSKlax66FJWHKxT0aleDvdqiXyUgbwavHcttdjbS7D61/G1FuAq6AAAWQdyKQfQM
6LzwacAuPDlEL4k94HktK05uLVp4bzUEEqmypog3leHVQtluHVBArdmfm7g/sqWWrQ66dTScNaiZ
l0yuNV6HLUeYmTxvJQR364VH8iiijfMiuvXZz80NmhUffC2kq32nh9mxaEn+UBl/emTJvyZAqy5h
YUPbMMz7ojI8WOpvKyi8O9GjU8E9IOtVcrmykgLY+4DZ4PZrv1ozzbgAyd1zQiIRHKo9ddONj7Kq
I+L11Oe/Nks3dFVX/1Glb+GNFVEmKDDVQgEWF2Zve/DZkrak5XTp7hBwNdDTTpEblinVeiDdR+9V
mqrmgUwktQuhQX+r2dP24AZPfDZnsG4+nx+ScvjgQqn/1ihSOWkeoB1XOppu276gKwcLZjYSqwJa
19j2TtCEK8VdPE4TV/4bJNKUQIP9lAZed3A9sJmZsp983X0H1313ZnpMHOF8ssilnsbe2uLTNd/d
OCpRpV/I0coTORRXk406KDSRHywKOgRNH0s7zzk0B6+TcHfqzM7W7RzLMcsmLeC6T4oVQPnrztiU
JpBmdbppHnEeGP3dYHybblbOeFsm4+0ODjOgp7puzl89WLLlUK5n7Je4h0x04ZDENKrNOHWljjxx
C6hjC7a8AfQ+J1blMIN5Lwe/jpRc9uDKtGKkwPGE235dm11VOAcgWluZtcS+0PMVRy5MvjiFKCRT
8SBJJ6TlgY6021vSq8j60B88FuqPNMFEfOb6BGA2Jt8ivoMUC9D8m06YHQHqwLxAhWgU07wtWKxh
tvBu5YZDQJcGnDZA9itg8yxb5ojQ+D6cIb0LpHZ5a1g7SHjVYv+RVm2t9OBnfm91NCvnjYUjJKC3
LMUvaLJgmbnTy82YP0CeDzk091yHTGBNJzKv+WmbSs4WtWCiY/ORpkeJ66n/QRLyr0IpURgwJ59t
cl5pIaOt/+znm70/zOjKENydvFE9gdx/h5WMRtz7Oc/VSWe93fc4BClXXxq/FX4B/qeZL5vtBX98
fjQKk75/xjTqKW0BNc9iGhVXW2HFJxqOkjop4qs3qq7s/nk4DLso9jd6qed5GcsuIp5ka685abww
2691xNhfva7ePs82/XKLyDpXxktPRvYgs6HvzbDRQjFfVzE/+CMqzLjIu4BdHmsXiqX5rt9esf6h
02yI71KS61uxqR5g3djl+ukP+z9njduYXksNYf9Aypl1IjD2wdgiWGrGISGzMxTdlU8VVPz3I5Vm
aez7n8oqbJFj2pNlM6eQBbWHVoAm+LfJyOWg1tStZWc8P7YpQUt6n8UQ+EWp3EF2SCIFqErzRnVk
ns4nGQFtqKx7WLlyA++OaoQ9Is3Cf7GgDxNu/2AB3KAg1z51Fnk+tnQuCPtBL4nI+0I7eXP/i1c3
J3rsmpXsqLv45560FuAH30KuxoG9l+iO/NpEkJqUxUwll2nbmFn88f7URJ/UHzE1EiJr1eVCqxtN
hmPp7bnwvcyKPR7Arnpu1SizO9RCArYiLy05nyGx4H0EbnQvuSZk6cHn3zhE2NrKjQkhRrbqo61H
XTvvXuAL4ULC9eB68ZfrOgKOXKW2dSWGIv73sok9vTxjnlsm0P2Lhr5bGs5ej2IJQ9DMedg9+Y60
dtEyTc7NJQBAJlQSD7IYA1YNYyWitHy45SOmPbBvJ3BMD9EzNhUMbCmmBsSGGKmvXgVRa+BGhQE9
LHf1XPC4GGt1C8BuztheCXySkclTlfzJ59ENaodc+9WtCTc3pLcpBfb8b18SiqEY3S+BCoONYSsU
vsYTd5jXQNZlC4gxQi/yBh87VQfKsnutlrx4IRZSTxxBelmmiE1czAT6z6w7wf6QYFc63IGF03JB
PUbCg/sWqNWcjeFb9cnLqjfg3FcPF84G95oI5Jlexsscva42Rn/UWP+hwoQG4o7qu/G2H+bPF56V
T9zGV0vin+8CqKjKKONFAQtECD+zBYnYoBROkB3HC+KNd66A4bJw6nzIP5Q+BEEAw0rTpBLNnzKj
KU3ARcMk5eqfW6vGiy9LaN/MCJIVd4xzQrS3bknMEY5xoNH3w+4SSRCP5aKw0zXB0XDaobMjDj5o
DdlxuEYXs1H4y2bWDyLmdnlCUXe9nO45gYgBDMgPOaSH31fLnI1byPrrFy9KJpgOp6kRSExK7gcE
dHgtuHmSeLkzB0U2h6T975pDdhiG53NX5BW/NepIK9J1VFKe4PJK6d9VruPGUZc/53jS2MViWZV/
SvxqkF83MDwU1da8GscKoUNDbWGyH/3hxoB7nah/jiMpjHDWl/rh49XD89El/VQnLQ9p12tL5pyv
2KvKeQLXWX5ydAPOketjd/SZyzmv28caw9pP7AZ/afpCOn7sR2LAQdfu7J9RVxB0Y+L3m7ni3vBS
q1mZhKpyENEkfnJ5+JRjcdrpiJ+KTkM5FyBstmwTpxsjatGH+VaPt0Ma+fIPcHZRSyPo21FIqFq9
1Mq72bBz7gG1boU47ANkjmhE8/U/rpU2Bi3KKYdGeRTDoXJ2Df18V7YMv+ndPlungdUQPM2a8RTy
Hyx9vjdjhpGYonxJg1MiBtQNvgYsrnGhiNopv4jCRrLhtoYts7lkEcZWySqrM78MsGiepe3N5hzY
+FoU706FeXgolL432L4tL02UJ5G5fNAoUIfpQiCxLRH6+HS1t6nbScVHQGUHxu38Xcbegx+NBpzj
xkQe4NDIHx0ZGoOrxbZwX8Cbp0+hZKyhUN5cXhWOP2hEnW6cl67dL7NFt4AFMTRrKtJPtwTaHA6u
CK2+9HJ5qrXR1Y1TF5oygdJQW11yk1iNY+ZLkvGslsRwAx1uhYJcL8c/O/05l4ExYQlKXoZ1nzaC
uOhSG1nD8gV0XqK1Nr2C6p+Mq+LlvK7mBdPYjaUwe8tkJTLwHu12nQT0KCJmH5fYmE2OOc68b0Dp
YgWNOvl7D2+sl/wpRt1hKSasNdpyF78/iCqikPXTuz6wdvdpUPWhKNi+0Qsei9YuYOXy/Ksti29D
oeGRHvKKIcIC6AZXUxJOh/rSArp3ZQvwdsSLyZpoSeeCzO8gLewzXWrNHjuP/Q23BWp5wcCJAwXY
8hAUMWPgMEVLz3qLBzoTil5gYW4oLiTYc9dbaKg+C36EX8lEMlDq6unCpwDBkWHfQWdbnbaRGXZi
yN8YADN6TjBz/+RunIhdrgGBzETi9O6r8jx8ds2tf8kukVnB121ewazBQspqtSjkm+QZS3iXHlJt
xfQWcBo27/tJTQcyI2RL218dETjlaI2pnkkJCl3o7AxsLTwybsR1Ze7EWkbrpoIU0l+u768kfSjl
VR6Ui9lICikmAvGRH3c8IMavkKS8CX+jyr3ssNLf6J925uuca6BqvBh4si54av2Ht/a48phtIxi4
P6Gk/RaNhHLshe2xfDmahisDaM2vCU0pJlv64ggk1JN82WUeM80ki/45DADcm5J/zO3g+v5T2qrG
UOC76616DdZHFY8w1DlFgiCq9q9awtnmxCrn5re6bkrcY0mf/nBsFZtG+ktO/xcAEN463AnlZKf7
ixNC+erWanKbqSdidSzzaKqFSxE3RX8WBkNNjVs4lq18lxefILOsj6K8YWEaZX5dEVK4xoPOh8CX
VZWlLbfyoUtzgzjvTZJ7OUoF/sAnS5JAaz9OL7dJBVnDnDQNiiKPSVlXojStsOnJeph1+dobHsPU
/5eCNXlgBsR03VKx4wqv30GzCycBDDKE6r1upCJLPN5O9qa8U2lmoyCGZh6g59bmhN4BEXaBd+LW
Xuokx2GtGja4W2XWX/dP+wK4F6cklIELs2wLzUY2tYagW/ROpiqehHgZD76ZmPvMO5lJa7pK6i/Y
diTaC4aYIAOFJmFbRcdDE0wmDuyTw2eSdJO0nY3+yIUy+iVLtq9YX9u620DH40ycmT5uJOx2bBxe
rrxMlBbsyjpAj1SzNRLadqkONgk6Mbv8D1BLShk6Y5qfIB07CD4nFu1TZJJl259lhjRuLHYCYUES
4auwGcnSIJCMgYBPODb/nFuhOMc6T5FDp+vFUp/h3XyI+enPvPA8/djgDJxL9+y480QxCPMtyz2i
zLtHAWKQPsGMhr/n0MJGWm3JkRhPLmOzOYcuKfAFKTnlYGuCATweHDcKjGEuwQSTHM8F9fV2dftU
jw3m/YMuC0VzfJXtGAW3Y1lkQ8ZBB1EyCZ3c9aI0ZUSVLAFj8LcnibIMjSHl8tEEbF7lBaAluIYY
5Lnw0WmuH0aqdp0RN+MTmeqElA3au2MJz2JNUTuKkkQ0tymxx0piOMhdfAGDDmxiJKep9f6k86XY
s02XUMRSGlhRb66WKVfLjk98+vkwsKCwVLvHpohWMAc3TA8MwZMXPjfZK37Xo6QeyP7nQ1JvN0AM
tWPoMppNzOykj25koRw4ctNxB3SzoPB0nWt6Ehnb7/trwKQwvJgzOr2cf/rdID17fOKLZQxC6uwy
spbBYS12/wY8j2jMImIDS+Y8AUbUaSr9sbz3fLr9WzqnSFm6PWILtG6aKAxuOiCXviLhR6r6EJ+E
Se57TYU7wScfhWTB91RLGWyfRsvFh9K+t8fBRp6+ZZ1RHubosVsXe+3LGG/YIiXAybiHwB/X3ZOV
RKZLNrelthmMIHbpBHcMLux7Hjjq+Ml6t7Z4dfLmHb6GxaNahks5vpA3oVhKGNgZUpe4rV5ofeCx
HvhsOD54mCxxTI77e25G4bXEY8FY0fxbA+OFHKYKFDNMYI/LayL+78U1AHGTKHeTynoYWSVYENXf
R9mi2CpfwP/rp2jZytNZjEMg0LLTBRTAxz7tFsiKxT3pZXMdtXXMVoacltebqp+mOzUhdkDlq1Sv
Jxj8LiQO7f6YN74bK4hLkRtkOUPk3+MRrQPgyLhOfh7NMCM/0lk0ZB3MwX/sAJBbUyZQJHBpWnkt
ARfofweyql60m+KVeTXE7fM0ChcnWnqqUIxTWvZ0J+57cQ0a2OR83Kw6q+yhxkR3lGMYv9QBD6yT
DLNxc59G+6hqEjGq6QQHQNzjAXSUn/DZ0Y+7sZovltPznQV+jyRs7bXGl3Y7WhCpI26BPcYriWb/
E9JLFtB21dyokXdXFKZC+cDao/TeinGJz5mdMwUMwrePSkhV9qlRUI+jx2keSS/F9h0Y4bma8JiP
20FEg58RMEFkPX+5KTtW8nqCRAeMgEqFTQ+7iVj65r5MzuZU4xIRN1jJfskwiiKDX5vpEfnJGPFt
y/4iGV+rhH0hT1NY/IZqdWmQocroQNdPSaOvR9VcLzewe7sPWpumnq8iiwEtaf5MCGHyE+YGBE08
CNecy+KmSh+6kdXiCUllykVjCXSrJhfxuprMzBaO8g74MpUYRBzHYEPJPaXLxXEbJrhc1R7PK3LK
zWQLpwSJMFHImf6qKon31Vz3sF5vpZ85KRewNNjztTMlyAkO1C7Zu00IOzC/hq9Ok2bRTLI5j9OV
cM7MFMXiauwfid9cszkUOvsQ9IEdourdtNe4BL6D6HgqgT+pukpvE4IGRKzXJRLl7oU5S+5xhFxB
XENcIHyAfxPxSc8dcHobwX9uaIUJBl2GbkZngi3qGPgVWi5jNJZpx41jM54zD3CgW5YdjS8NFqKt
OZbFzu/boPuToZNTb7My9Pmq70dglO4PspQZg8JXIy27LeA61SrCy26iJDjyrmapVfuyJ7oh6LR5
iw40Z3zy2XVLMPCX7x9/vS3dSGGIM2mUrCkIknPdI407cEPmCTk74VbJNgByYTm5eMeSlchhYU62
7RErIaiG5FBUbfN6UR3eoUAwOixXtxfyWtyu0r+ONvpKiH5uKuVeWQvrqUGW1RjXA2yFO2bOl3dp
8TZbK7lDiccNzLE5Ns5xhgZVhsCF8V6U/dKY/pjhdLPkZNdMPPDzzJZpsZDOHCxjYPTpcszwkA2o
71joSpayFoeAM29BWNyWzXFKenOLIs1bEjqf4LDdl52+We+W3DgFXHEGGPY1aFCoaARSJjty6Hpv
ULhR1cSM659eLX9YeSG4ktqadpOOBjV4+5mvOwdL9CGJgvY11FeLcMWB8npIAF4G3nvp10QS4BDS
c1Sji9liii/LRVacKRofwx1EWle2v2BXixAEVqE+mfnBoeyArRKBPpiXg1F6OfaeIq/smz91tTDt
DqfZ2AD7Z0WjIfo68YSrmybv1upCz4XVTzMkKB/dueClA/tdhCy5OsvAua/V7qdg/tVsBkk87IZZ
DaVDZq9J/OzcpS2tE+SFTqPF5+CdYFdAulotIBkmi4cRZ+DjYHIT/z4W5deyaPOBk3w+NjH+WzuF
NOk/7YJTIUoWDvS5FIRdBvFUxMy30nXU7UdAorTCt3WR0F4XFMQv47gBGDytXlwfv9Pee9Q9gWfS
1jUaldMN14xvPdUtGAvgDu7YtWVHz/6hdWaO2c0sQgrxA9K4ry2b1XXEq92VgXvHqbolkLfRNNng
tkpr61+2NSFdAY3Ib/dUTe5kCYjU2yayBuActjK4qWo39LRwN+lbTVlCOz715fDltoGzdSTUoqkE
cIb2DC1NamPUzrNVoOzjwXIbIwW3IF5mjL9gnaDwfufb4goZ1Y3SNN+tavHlHucQOMoq0ZLEbx+y
wUvQIXiqLxGwe6tfgFAq9Kn3gAPtha7/kzBv21iswviXp/+988vSqctnqs3Vfjyo6PmHSKvqw2CJ
YA5yRDXUDtaGeidGDn/mTt/0DRLm5PG0bYEMkGpaWqv78Mwaf2plFBUbQ92obm7MOYa7y1IXCr/H
NIWHmYHAVdBZCpMmuFoNUnmE2wiIbqRB1C8t5J2HD+SUVF68HkDprzV7JnP14irGssp5ZVvZngPs
5dOekK8UF7uLYr41C3kwmllpRMH5cQ4REy42WxPwghZRT1El3xN7IrU+TcMK2iFtOrgPtUkydzJR
mhlNAGVKwkzp6X3JKDxcdG7RL3PN1EWFzK1OydEEUv1eZ6dDCBYFqQxz/pUQD54ssKgxnZEIr32b
xpOBPJ+qW08kWJg1RFQXWn+32wlFjGqvMcjW3bau2alkPOzksiVvib23xTM9jbQ8oQfPtE8FS6NS
U7TOeGq4jkf1v0bT9MolZURnmgfHRmbP3j8GjTCstGdP7L6y7yd+578mD3f9R+4IFK7crOMJw7Os
GJj2jISZxy0+TtsF1lL0qAB1Flku/3t+sN56J10DW+58JQHBHxn1rstZAGSMj/bvNxBgRifz0KLc
p0WaVVgva8tSs0ROdtqo5ozLIwhC7LvQEFK2WG+CZWzX5iI3Chv1QH+IPp+w6y0tJC47NWFh1YTQ
Mtn8UQWsL0qNFtA8WCQZdeDhev1GX9yz5SYw6rPA/ccTVHehe4hDZqjhRKoJFpdNha1bAFadAMBZ
nWZA1gUUCstrE1yE1xIYpV4tjm91W5g0ZSS1r/exGFRnz+mSaUuvKqbat0E9bISDYxP/+5XmiD/2
u+0xOc7cCNAeEBMhaOyYlcm/WpPxrTlXK0k96oKYdjomGUQjNWA0JaEzw14MccRaOwJLDCI1XWsn
JF2hrla/mRIi6EPuPVm1TnSG3RBqmbI6PNAmNCgb1DbNJD4zg80V30ZgoPNPW7z4t1q0h62FkH7W
0LkzKm2Gz5G2VmDm8cI7dIm+IJAEtnG7+Llhio5Y2QbDATH0KBCWjfPnDKeQ9ZlmfC/hYnuOJ99E
ES/suTHyykl+yQt3IsxZO1xzv93ifFbxjEXyKe69JB512YLFWur0JwZ12vGwgEcqV38ARirji+mM
b6bdQdcYkYVTiFOw/I14FRwYrwNLV4Dm3HsMumfUCOzq+R246fXUro8j3U3d+AToDbGe2Fg2OkFZ
IeSGpan5bXNSGb4Nep8PKg2jP8N/lz2e8X/Exo5VN61bKFReQQqsURjPbZAmxXF1U6OwKFc5d9ri
9ouOCdEu40H2Mj01WQxs80tr0fAUIua4ZRmM6/CZfNv7gbJ2FjugaLKtmLBamudRv2rkOeYDxpbT
q1+Fmj7grX18IS8gzGIyxsDLazsgF3uO1siA52geIwvv0aG4iAF7CHPkGonVN3tcnEycQx/hZ1qO
RwH6ZpoTvf2OMmvzSs5g1NJk0xFn54yJpmqQYddfmJY+XwJ+OBk6d9PMOxCG3ZVIKVoUf2FN2hV2
Yc4lWYi3yFV25l/IdvriRRW7jI2QgJEBlCtQPFcLi84e9Qt7oKvcXPaGR0UdF7bUbCJ3ULlnBZjl
76jqJuuHLDaLHqsUek4mHGYWaabVlfvmH9hO1lXPWVka3ZcliVLrtxb/oXV/Cw1lGff8a/fFLBDH
QaKhJx1O0DXxwQLycPaeRZBeY4e4xK+tLjIEvKBx+x1woG9uCq5mALlrGHcTgFXArWxMo+dpjuCM
XdWUjgLqGr2bc+NWSD8wCnDfp2Se6udk2MOsh36xCGdovzbBogpYSJB9aF0DI6Jw0tsJGFN7wDGv
oB0xS8mLPga+hvhj9+aqorBmpjr4AuPH5AytdYSZPnjNq2PW7ebkMudA39FXs24f88y3Su5QOK7m
HMgY/Vg7akriO7v6r+QdASArvsi20R3c76UH6HULaj4odBU/zNFaE45gtrdAvdpqz5qaJ0HQWDWa
41tEG4IUuVlPB7+dlTebd4d/D2NyHEmwIu2by0spsm91YLDbiF5PlfMGcE0Gvv6w6c3vqhOkVsYd
3RVmyqYkyzl4dgZSzcaoqNPn6myuX3sPP0g5YRmcTiRDNkTz2SJkjqC6dUZ70m+x55roru6oMWHd
Aew0g0idsSZBMs/T0s91mu8/r8KgeG8HYeUldbWt6WbVVCToK0VwODHve8flgsePL+2LLdBgmu0U
HYuhHJzHx3YQKgQbGw941RI1asnQLvlDLpGLhbQwZz8rdFd3WBp4QW8JInlGp29MRhCx0kjPlM82
O4ALDHuTFQV80/oleRONJDA6Hw610MohoALJ3QoFUbpPI4eFG5KSv9ncpQGCnpRZZKse+vVlJgEN
ypSqFFlh1GSvzFU+kQ49Tq1cxYk5o5Preu4eb17HzsVTQNUSghpbWOkFxFLSmLM+KFj5P9qKfHRI
0HGI9qqOOFyrWh3417ohgX8VYf7eK7Ps1mA5oM22bzXOh9aW2v63mEhBlrq5BdmAI4bx0xZMSrMG
rYpKP7+ri5dQLraTQheiREZf1KAFnRM6WNS/Dc7N6AX8p7G7Ts/hu8axbPWLO8nxKmYMNJPl142+
cGQNBgDP2BTF6o5sHTR9CdvQiK+KQ42CKN6SiPoZvNrg02e/F7SgM6RxeQMSW1YWVdbeO6+ZPACN
j5Q8yBAWO71i8ChOmQMyJhbz+sePF9vZdwGj02gBGRHnNWxePcE30jB3mLt9WiREIwlcL3+AFObe
SLD9QODdd47nShC5j4BUxSLEVEPnn9RSAp5bTIdnVfJb3XvMPPqa05IvxjwIj2l7etbgc/z5pi9q
bYw24sCVhhfjukHPuI27epWTGd667ULYS0o88zkF/LXNDm3LhoYk1TEyBZk10l2Mgz/8YAp3kP97
nwjN5atI/sohCb31JaUUCOoEuAG+QhaPg2CicgXP25A64n25/H4QrgB7ca/GN54FsNw4cZMPQyBo
RJvc6B34kgMdw6FVH3yTW4pLrRT3E7U3uG9RuMB0xC3v2E04OEwZvFh6DMkZYIbvvws0OhyxCFao
5XWp38lS2kH50d7qbArGXHIvurj1eRTgNk42CTIw3BK2GP2HV//BVFRjpcs+P3Z/xbsgMdhIzec/
R52CaTHObndZ9JH3BoCjv1R1pYhKWEivLhsj+5olmiVHgPb47Yrjrl+wRdb6kdpONmBdRXTEKQoQ
jzpX7E69Gbc0Vs99IX/lNBmggXkcWQrhFCvJM467hsb/u9gahFJnmFSS25GS5JOCBIJniVKTxSYn
aHZXYcsDfmVKS3EPmkXe5MFN6IOOvdT6nYtH0MnBwhL9VrVR4yi3cHRpoAAhM+Iu5NxxZDwQfVJj
nzHGKApWjolbzRRkOYIl+tbaDJWdg4S7PrkoosV1NaE4QwzTELwY6mI3D/RENcqSt1DnJD/xxIni
bh/kZpysQxJ+qxGG9ofJUGiLCjYx1orVB5tYfn4jOvEOER84FmHYBsWEXxb5i37x9oHuDotJeLjd
p2iEfVxs+vBqLWXJ4fvFiCzA2ZvGMD/44GAohy0loodMqLMeNyn+31cBBMC2+43WxAjzg37jtrj7
Ndkoyn0+bQlL/bnggABvJ59CTKBJT+KtygRObpKkXxqiKbsLuks664gpj/X1sqcwdtE2Cj3FtTn1
1URSwoqJgoDQ5UCTfHHBPg5C5GXlZL+KQg6loKl4bMjFbiFpcyFfDdJgefw0/88K+5BaCtqYmABQ
NwqDX+nUwEfCOV+6Mh6/mWrlkne/1xqzx8D6yuqnbcer9F0GR14r+Qvcz8qFPLRGMR/16dcFyahx
hv4Z8yk1SPXKOvTFCIgw/IigObXjplsDBuiTFmbSyz4xRO7Un9/9foHIrbt58r2OMyOWgkCoB3Uz
/PGMl5VnEcCi63ggbCT4MF7YsMYoacSh14hKCAAcceo6yXmBuryYhrFRjEIsKWjDmQkxSkcDz0LA
coPz+v02YMONW2lwHwA1hKxiGn/mBcTr5+1wI3YqCzdCCW0LNCuqKV5LDxtaaLyPY7V5hMStC/yy
HtfuMOSmawkmoObrbgzBq3DVeTcXNziQRfHEshMY+sjKOpWjttsd5XlVrOE/IjY5WgFST+TC2X8G
ZwiPBdZSkBK0tUU/Bo3AJuQcVm2xV02o+uFXRXGcbKGZyL8lDDFA3sDbkKHLHLY/CSi9WJV4G8v2
z0Rh85XK/hr/YjMiVenejZ1bopLN06g5EPA8CB+BUHEEFy/Sw+4yzQOZy2Nhn2mRHeaWeGG/QJ0n
eEsmJzFQl9ebe1idP6sg6rfthsxb6QLE8SaQpbengbCrQqXxxO38F/AikAbe8ordOMkTpJpz4fH7
vG73i1lVuhmoIfFm8TC1dKoONmynucb41A7MCzAan06g8CmVxE0sj1PTfTlKmk1sChpwlba9IHL9
mghVCEVeQxp+pa1PJqdUKWIqfxVWxtcqdsWbO7FWu2jNoIz8koWpEGzpVfcuSUTH01X3Lht0uIQk
OVzO8aBj6+OPG27HVA9ruuYtLHUMqmMAE+wFFY9IbfuqsS9QyUh/GGvuw9leC1oqrx6+wJ5oMx0V
39/fQ/so98id1KKloSip4SCpgLIyKapNPfZVQekGFm3fIbikRRRGJduYAf9UOyRjx7oCg+h/Dosj
6xQZ+0jP2F3s0oObxFtf5TwHw+tSdVBsxTYqyV9CFDwkN6LWOrS7RDROa0Nb1WdOKO0BaYXrAJy6
oyCOtvbvExNW+AVQFSflJZIY02yRbEg7s78XB0nFmZAO6GiX43yaRaAUoDBS+CAzWt8mRerl6Ksn
fAkzEE3TiVqZKzN/stoJF2X2zXrkWa//j83aPgwfEUWvA4IRB7VMiD/A/H30Yrh0lxvgc4IZS6Fk
AeHYYc7manALxgw6WZelPBFko555TgC8Z4JgzccC8RZZrYPjiTfL3mYwNYGUhluV2cs115ENCwd+
y9wrYXtSrsjGS32XjgC0XBzIRG5s0NyjBytO5xTB9qt4uJIOMNq1Xu3Mtg9xLYeFgAIwHs+gpPbH
RLn2SGu5skuqnQNW31L2FYSXNORzNCFryBEu+CWY4ArNO+xU1wK7/LjVWFAhZoOE/ujwgjUNOi7+
e+kxhluHXNrHS2JOaIuk7dKCMrVVIJwdJ2z4Z4owQEt/SOKzi0XyMwypJfTQoTuCAmjMhEEVSB4I
QT2raaCdLVdcuFh20lT9s1NtRVu91JKo1Z67h6ArQ9G0A3uobnD02G9ER9Tcw2azaBqopqOO/82S
4Ltn30H2nugA11RllNtm1WENqvHWoY+TcrYuubTVEL2xq2Nqy14HWrNrh6jY7+CPZDouDr/T25Bg
EyURVqvf/EajXJG5QrJrxlaNvMgFU7T8zO8qlX6F1aIzpcpcM9x5MVxc+OufeLsRAvyQr/Jb+q09
+wyriP7lZScIpWdkOZ/E+Cw3vY/68HbpRW24C99CdBN4lrccGwTM7yW7Zt9B3ozHBYBuP05/ammV
HZh7KR/TJHgt2zeXGuwGmelHbqLn1+GipEyR8Wm3q6CI/MauiVV7yb7u/C8t9O9svccvJrPKvEap
69VGbp9dgV7UDXyKHavvlbfIot6pdhDQV3soSQu2ojcQemN4HXnczoWij5bEcUOyq2dfc90d/Swa
j1r6RstzlruieNZS1ot93FBERvKxDsJvG1SZPIOSNARnTnnAQFKJq/OQpnmWZySZz5Hv3jJINWlT
6QIGrlCfYHV6/z+wa9W0Rqbt72vpnY+MjLnP9jCffVUFCuO4vM5OPhHG4e05QglwD7RLrAu7DasN
Js4adsaHN6NwBAywhlZNKIewknNzh0FEDg6zCAb1hfa9Zo01CBnHjsE2hvadLB7qfxsEvlwylYWv
Wsh5TXJX3kHthCISsB6aJPlek5n0lNRWz7/J7du9FXZ3v5HmLFoil1KmnB2St6a5PDaYV/68kyuR
+pPYW8zKnMa6Yn2ORCSiPgbpKnTwpl4vtrEsrMul57dU4rwVjSPgZ3nzj9qB0wGBfu3gUcDQaFty
EciO5spg8E7EpXD85msL/L365Ag31oXABBueH4MnPCN69N8pmBNao6qBlJQ+sUGUoXq/LFsZXoiv
Ib6v6RHHtwocH8/siIxGNP9KkBR17wWpaXdWKr663h0oGDeBnIjHNPGRcBQlPSCYPjMcoHo0j1cZ
eVkAkBijf7CQ7oah55w3vkixkpwxDzwOWwLBZkO/MOS+V4cAoN6E39ItS0CvHwHVLwReaG9SB5QI
wGtjZ22ryEMUsPG2216aqU6NT5cd/u64SdJOsKo/IHQTBYcPB4L5g6S28vUMP7UjIF6NPHvuVjbC
wJt6ZaCwGpbWeAQ+GS0jLBxjBwRUw0zRMhB/hPEDnGEhpILSX5Fc2eVPE9I9d3zHe/tR4c3TKbU/
DIrgn60q3mrs+Aly4B2ZDQQvpPhBPF0mturfuUWPg+DM2CNdeQemf+hHm0fykeYqTG/DAF5nkP45
ejivSsdO76fyqVWajrGYLxUqx3gakZMziqkcPYjF5qj/lLy04o8MzQdsBcJs9Ijg2LKBA1WwJmV3
NG5Lm7prNQN+PsuKiu5sWPFjiPQWFKyy9B4Zi6yQQLrxYrPucPbIS6ZlB5YdBqPT2bcIpLAPAMec
b0c8w1H3OaZ/cpSKblvqXxFPJPu4OOLy48x4yX9jVDVBCRKNuizE2mrBqoRhHIoIW3V64GbNjOa5
bFY9NZXjBzFFwmAzMgg1GobLLGTiPpcunYCQy6BLNyxmiIJZOtKnkWCtCvdpqfkXUBWONOEUR3/m
TqR9jo/wu9scsxks+Siy4Zhjf/Wm3gLS7EiepB3qzOrp2T0GBIY9tP83rHe5qIkj03qsWdYPNTbA
buwDiXByWjidwlyOtx+3BKq1V4UrmxkOKC+WYFEv7Lq6LtxAQgz5yJvXBJnGRDmne6JZ5niN7Wc0
721J4JWb8dGlynAKV+sLRAxgW7GLTRtcNb9L4VoS0YhVT0mkeRrT4F5leKTyLKbcNWSv8Qb1IcHf
/XHntUQ7ouR46F0ayo4AUhP2wyK6vZeTaZ6M4l1nuf0rhCJl+jSuy1ok4mjLqcKYbquVjwAESLWf
0OIxDy/XKvCzPLONY4urASkLfSOhTZ63ZfV+6CSZxgAXehpgijQ1cAiFWHcGzyICNxo5DZGorI8f
1xvKpl+BVNZ4I+PXxIQXuCczedMzW4wDmJZk3fimR2DwPiYqzrokS8loUkSFKmpoKHIpQ7bu+2ZQ
dofK6UIISg85hiyOKi8yWh4tY3CC3N4vPP6gdLM7tFgXa9TlbgXnK+j2G6XnfGG1qkF4wKqUWX6F
Ao52eb2UBrfAEHJ7fjtgVHTOZLmTgQJccgpzVVdka9NdK8TgdYbG45D/DPgfbh+nie+nOupPPxRU
WyG1zmWmp9W/PuRghDw/JCiHwyfJg9+q0zPyfyA43VB2EclbVWqgTAUrcDWxJOpXKMtXf8QZDccF
t7qQeY+zInPHDNeZihxgaD3lxJqHdbaUqpGIdjpjnnMZ/aqKCelOS5+cuivma1b35S/Oy62CSMcr
EUaRJyYKW4fuFhb5WAv6rtMVq019NTZiUWt6Vh/aLwgbioxgKGIiCLvmpfsg4w4vDd85UzvE9o6g
tonsY3c7p+Kjn6rY8lMwhiCzQUM1MsVYUHtcuHFQ76Wb2qhd/XcZ44DZo30vbHd3R6IQngoQ00Dg
LjzTGnKyHEtwKWnQUu1OXt8Cd9+j99oLt14ew/YR6pAe1MfhrD+MiLZLVmXqk0qYIZJ28ULSSol/
XCfSolx0O19dxHvVKr+Lr1Ipt/9vP86bPo1bSbIE5lZLyrZkX3Uh7A73h4+NrQij1/w1MkFpt5/X
EgOdC0ICLX+HgTwiTbf53Axk/WrUGdCS/GukfUriQNppzbJa3e9XtiWGKR2UWEl8zYCSFjS1t/OI
mufkhs58X27WyZ430xeFMQqPUnqR0+U/J8qsH8+sUGEO3qSwhinn4ghnHghcvZdDvWl1j26hT7hi
mxzs/Ss2lymRSsEH147yXLH1Tevgq/WkSj4wiJQ936m0/Lateqm4nU1HCX3orEpbUUvH/OoE28gY
ye6Yk/bdvD8ZP3hvJi7oVhPx0554CxUVVVNDpIlUE8cmHerG7f1pxXFJO/oOGQvBEoe1nDzfzbEl
4TVzZMGaiIbw8oTm59tb63+FXnL2MGTpm0Ws6TiVd3xA6hELgobhFT02MLxEzgRKQ4viBqh9ihek
p1Ej8n/Bs63aqmiWlR3NGrQAhB2O0BZ7JrgLHizi1D4lBCVscbt+1dZXB86HbUekagMYEXT4VUBW
1drHoGkkhO9jkX+ezJ1E5S0tehpHeklXwetBV2RjOogKRdl/gNvW72EyP0mFdQjDDjBkSFNZKbLQ
oHr/UozjWM/K6dkM0+n+Tca+mtYnCzHrD4ozKJ1ZYDCQlpJtizIds+iX8mz+nQwpCf64v595daet
XH0pYFei5fRKbXoD6do0CEhY20GJil2q7sDLn/0P4cH/3f50MHurLeEOj8cXkOorNpW1T8lqBI3p
zHABm8TyKKgAQoEgHMazpOvK7EPwHIngYvhX2l3j2lQHkoj8vtpcBUgOJMzEh+7x/swehuJ7SeDT
xKmYCbxxgvFz8Z5lRCr4XZ9QYJAkTSeGfkwg1WvVTx6IvNxKj/umHcPSj54bIlr3WAzSn/gGfCrr
wSTYtOu7rXb2k+IznGHGaZGtXtDefDCXW3YzRrn7vAqyMmtOf0B8eDf+OpAajIcOQHQQWhtQDWTv
PJJ6jeaXykEM2PntM55k43FsikxfVQgSV+sy6Sv1F/av5RKXbvPH6S5xTb8r9n7USMp13KNZw9vp
2zFp4PrfQyI6DxcrFdH9pQ91HmNUOXNYJ7LFVW2E4mh/heg2OceJ5+vIRIw8Nu4z2K9dXZXiRrpN
jQnUEnKV0OlumY5fI7hQ7lorhDh+pnOZB2bl7I7sx+w4rMe0hATalNg9y5Wsasn25oD/Pv3TIJE9
cvos0I0M3JGdCYG5shHpGyI/ge2lMY2/38qVvvjEK9dlbKmhFDhA0vVtQlUBYRqskDwhwwGR4Qna
kw+3rEBhV0duE2RA3i0BKsikKCRHIO8RzEWcf/9ZXtXN22jFyKC33/KU6x5E8I3GSdmj9VOPSbbA
uKkY1IltmMaMIHAVkgylPbEDeznaq3JHJGNj1yV1ForxqmftTCRCKZvUgNR4Z2YQIuEebH55FQso
AS28mKWemYbHQsLWpi2gd9W5u2adB/dZLYxxuCidq6wwlPPSDPaprw2jZSdznswOSoW89l06Bzh/
X1H8S/p9QD+DnajybaP4qEoZCxLjlcrWptsr/ovxSMl9zBnXCi//rcZiTfA1+yy8RvpeflS1U8Lh
9uOm+FWFDc8dar6g2tKxE2Jh1d7xFiSrUR/9wSAPU40kcmEHOi8x/JBTkGIhsVaCEKg71BLL/TV4
sTTeGR0e+9zmL6n4MQXcW8pbd7/dlO8MhESgZXx+nSmmLBNXaJffoc8JpVvBDbLD4NnuVQ6FToeC
OzLjj8iWLgWn/j/blu4DO2xpmmJBH4gKPzx7TAF4L7airgud+BPqHcu+HxqOAh7kPSzjDtl08vIw
8swy5ZA9IPDkifprItC+jCzJ9UeGou6SXdJD1fIisAdwuIzEYPQB22a20w25lZWZ6ZQ+sCh/KzQi
jv/b10fbqHwvuvL9cilyFYZgzE49gx8WYq2mkX53EFi1GRWmrvSXHsq1JWO3FbmbomvLKjbGIR4o
wPTu/FHe5nC8A7Cz5s1U1dRmZWhoCpgMs8Z48EFwYoR8j5a91VRLIFVIzJK7779WEQg2j+6AxgP0
X83vvs0aVomb3yv4ezeusT8Bzo1nrFOagdRh+/OyGnCeXi4y528Luxa/gtD6O4JATWScXLwgxkAg
3haOU4EHo10G9fg+CCVM6a4S2N40X74wPsIgumpBfAXJcQKB+TNws7rRMXxs+P6MXmcUgLqPSTjJ
lBzIfIfG5mLYrDyguNTQStPNDhwhY8ybUJDT/fKuMSGhZZOr7ajqXmyLehb7hxBD4CIEfNPZfUoO
RnIuQt4GFlivIUdP5THnQmOnUsaKTOhDZ0dZwruBW1usx99Ap4UCK9GAsMfVJfME00n0x6NSUuIg
5EcVmPJNEekSVPLdsALCc7BwFkpZTUVjvWGbfRIv9GikLbDvldmYjFGYiIXLEgDVFqHOpH92f7sh
RBtDPwp8oaja11nJ1G7xx6imwOh6MAll89ri2hWWR6sxuWrtDpEO60+Ufj7yiqe1HlY2MyGlBmJ6
1TDVqv2ejJtw/lrWTjKnfxY9VBZ9xCvnh+CIlUFULJBN5Dn0eRfLS6YrTdZtppSN/3oIzfNHVcr4
qAFZttt5m6UFDwxDKNkFh+s8EG4UYr5R/RxhRB9KVTJ9x+1kRB60lmCD/065lWdkStwfPP3eyMyu
zy4LGnDm900Y7NIPMqaEn6PsK1CAhnbNG/jZ/z9o2pwB1g7/Cxibbz7XAEYleqxW9rOOXS3Y3Ure
cli/T5KZV+i/jXhfcTKpr/EeEvr6KqgsP104XdeZONU9+w2Q5m/Qes4atdfnVjr3C32tr01yDV1Z
bmnuSalzQIiX1zTzBiawLon7Xk5kVS+sanZZihlIq3D9RL22c0k+rsKsvJoqKAcucFbiGDWMQU3i
4xB7vr1+ciiYKflsB8bUz/RexU/QD2rtT9bs0eUcmL+KKz2cMcntLxrEvR+3pq9sprxWm1z+VdEo
fyY6AN8OCt0zQZ7+lY/fn9yBZaPSD0hLkHbjOLCIJ8XSwc3SzGFUCjZrPxX5zadQkRCgmFSJOCGR
rz6TEbbPziDoa1uKHU9hM3/98ZsMK5qgmhx5u9ED9c6ngEaVkpf4RY/ZHs0/2zgkINc57WWTKEDB
Eg2QdsUozPhBFTiTMeeA+oRg4iGO1dJDQWaWVteOLVmvLtB8KbdeVZa7fDHsOght5kMu7PrsltF/
5dy88hT0y3HhZjwiTCwnOcHv38ZX3wOKeup5F/d7Jbn1PwkuXhopTLiD31BF49UovrBMomMR0gnp
VXp3mZplGnPE0r9DwgYQ+fmrtRpcMq0PQcbXqL3xIkyMguBR3o1IjS7hDaq/zDD8A7ApyKWI0J94
EHsuQ6XUmOMiA5FtJwpKBR+14uWzT44ny5xTBn+prtwsj218pHglqg5i7bWK0niRLy5Y1huooclW
VQWbAouYoC8ucbGyunUlxENUCbj80d50sWMBzhAfdCzWyf0f+XucE1aB62VGz9fm0zLaszsewKal
GcPQzTHwAAtCGOc6v/mp0GlV0TvyFOzB3sLtP99ZaUlRz+OqWCgVWgxuMSXmD+5oxkz3lqvpqK21
qH+Uq6YODEN90TA7beeGPJIFZqKxSd9OGELUrAktABTPFJm9Y/dNPemt4MXsLeMUvoREHDlBQzDb
IsIkEPy4Pv97VglXXEZ0QDIAlKv66NZFnLNa7z79Gf4OtMyfDAKYA40xVGgrEeW4Cq2IrTLL9CHK
OqDjHLRcCZjptLDpARdj5By9SO0T2enmBsYdsnkjaao8oaxT3AKkstMpJHuEjvSd3acTTio06+g3
2Enj35G9WSqNj+bU0iN3PGFtzLD6go2Tw9F+PU4iUHne5p2RRPRQavBe30qP4KrFyf7dTwzqR1oa
3d7G5JP9D71a0DyYtXmEaydSRmPOJQtY0PQRww6yjrjxtPshW+SEH8wIG08OvsCnnFUVfxThbMvn
QVDzKQreFoRQM+pB/jAQwolopWV0khlnYvTTNUeD5niUzTRoetzt8q8NPJuQF8e7qJlVuMAdcgrb
jRIAb+ua1rwNaRXelMc3XAcVDlZ7b7hpOmfCAPcb7llztg4IZ4h4Heb+rHen5PrTneTN4TjPUr/Q
WeCLcMH7sti928dgc2yJNOGpJEgK232ggT+ehQToEFbhRS9a5LrqGvTOb6k9bfZv0FWP8Ut7FkVY
aa5DORExPm+5S2mmemcs2LyKuMovmp/G3A3iln9lmgu2aA2CXcQSbgEr5dO/zUM9PDHqZqBuk3YA
J/9KKpTNm5rYmvI54ImVX6yUoSSPplKCOKAUe3onVWwTmvFg853yLq/0p0139evANeyTxbBdla29
wZlvXMFiqNSpvn0QiL/4O/iv6GbL46mTpRobNrmYWXAouhdsR0ntFXdohR2hyeAc5Q2sOjg4SGT6
b5wws313JRzh2ycInzOaGI01ayeE3MAeCDbO6XWLMq+7A3bYDNAk9BCVHnW7goSkyyhCwVQ06mxE
6O633kTYxFeF0cDxoS0eLcx04FRQZO5PWidQH2ReYB52xK0e4qxKBAAWwL/Ngww53LR6k9PRHESC
DseTd4RBnAH4M/XiTubABRgQUKLHc3TKMunqDGSMELmRiKGFseWVvc8mgUXKX92KPPguhg9AVezl
FZ6TjUPZR7pBfoH306EV/FlvqX8d/KhEX0Sy5NHbg+gYg1GI1H5G3PKwKsAPECUqIQHqJUI+xeA0
nQUC3GnSMLvgPbliEhsyu2aTMAKRMGfPfWtDPXsVc4QOwFZjYqN4vajBZAL4gVnJ3cuA/s6uBghg
B1F7APILqeh9pd5CU04tNWDZwchsrtPp9mjt+hdnE4zoKFrT3vsXaEO5tnC7dunpSof6aQET8fyB
XLlWdBNKQf7ff3zyB1o6VKiqBgyZe7e2V4luIzteQ1aF8hI5lNscULDP5pUhDTG9fQhwQ9fRne+m
kGbR9g4LbXT0uS6M/tCc2X4y7Yur8oX81DGjj0lZd/K9RHrfPbomecd+9jTjXWYfpkQ/LQxnU4Fq
SeroKFrSHsgPrrWE2orM/zUg0iv6pXCAqsubXDKu7Yef9yLyRmQcgTFOZo0Scdj664xz27pvMM6G
OT4L53y7IfqzfZgO8/qn0OQVMy7qMmS4/SJ0sKBpxBYwC7z599IcayfZJ4iy82b6+9s1xC/E/DIl
r12zeatn5cxa+SCbaE6qLf84e7aVR29lrT7DtNIAkJdY74SDyJTgeNrQe0o9qONua+u4o9NeyDxJ
D9tZ1VhpebieyhTQHUl1Xnkcei2UDBczkrHZXfwX661J8ea4kakkf3YBPkuQD7MWP8EX/K+JkWMv
9yGtCwZU8SnBeufeSGP9hOY+/XGhDep+FbVQ96d5Qz17Ot3huKgWoFoea4xO6CH29XA+ccFzbhke
q3CSqRAJ+VkXI8zexA1r2odUTAmzYi6Y7NGRmLepSmJkhOp1nhDr3zwJ82h71ugdWbXflITy34AT
vQxJt6e4RcbP2bMIp+DVYHMGNK+dqG9VqfLST+rH2N4dwAqvBHGAGQRb9ewazc/w6P1/NpFXOYL9
B3FUetmz4bmRY88AB0OYqc1AFnmOBStDNbXdwkTynH9I98ptLNN97b5+He3rhh3LwHuChFj6zvUL
FzQKUKAY9BS+8KxsXrswLoZV7LYzcVRyJKmK0a6txseZXgBzG4ys4i4pI/vm02sOvdizUa3TpJbC
a5CRwEZGR/P3zFgj0forA+fqHjwxd9cc3krEGJ0schicPXvcbaQbxcLIqm9eKZdnttX5nXjNNLlC
LXFiSG7NxF2ziBM9SIPUyz2SayFJfi2wMwOShIHaLcRphP0WCC2/aLlrNVbMlwFd9VPNMr20C72G
OZQCVZBpXwt3xE/jd+SXzlY8tiMgdq7PKKThbxAae24UXhPizzwIi6PGLx0UGizWFaeobvY9OF8y
N9TrbQ/pYlR8Rit4ZgHXrL1Dqv0h55Wr33s0u9KxHNTF9t1uAhgZ/e2fbYcilDqYCGwgsuJ8J4OP
yXxhU6uf5zS2QPgjKw33dxKU9xvJhD6In+Uwse/MLUbPOKApCyu88s2oo1Qe0u4uKgpDIkWDWx4r
VMaVb1qk5NfN37Xl+DBkQedrbN7Bm5nvm4+YXrt4bYj9Bp54EMuEutLjv2l7LRb3MoLLFKDxJIlJ
gTfm32jpr/rq8ECsJkVSniphWbmMhMVGLFMF6jA+dDPiQ5+0jzEuenwCW55x2L4MaQw0F8vXop+9
W1qhEHgINDxqv6jQDYUEmZ1lUmViY2KhKS0T9v3L5BmzbPROOuTGKeuQLmNVfpjvrZ7udMMuy1wk
eRpxSAvIzwcBmFTSJ1W1axCnCa6ILyO53UbazKrnuPbvbJ81BGMOsN7jh7OYQVQlWpC7s4n+fDcb
YcTp+dJ5AIrr0De45lR4Ekuank4VpSA5HqLvsW0n6UcBQLIhYYuWhuyTBAsjifLufI+33J9jAd35
YGDlqZ52WGVrAycHeeYosG1k6mQ9R+DgSN7kn18/crzojhk4CmgxFQoLq6iCMguEPH1IfZ6BPtAr
rEh7WfQlAvLbVYwVRdN+xzRGi/UpqXFKh8hhdOeCkq7cj3Cg0yZyszNsvv69Kf+aCJBGXjIavOrR
LakvTnoX5pA7bz4PuVWK5rZ3tqzw6CMWonLpeoJd/HO6/8y/MS4f0l9wxMtLyZQYVzol21Z36O4Y
vBLh1IIUHykmfjxWSoHHAe4NjqRgSKlakOstzl4Pbf9ocSIeCY4ILnVmCTa8MmPCbJjdCo6H4txl
OnsH0badxPMR8X8+My1ZuaypCr0TXMFxdsrWlIjhCviPCbbRNdf3EVMBhfum94BFjYKuWv1RhA8N
BLYij/iNJE9Z4fhviLSAdCghGTHqEdDBOeM/f/QmzON2RJyVpGXfU765dSD2rBKvKaRvrYT+gLVl
/DGfptdjd+XC+BH5Ke0xMtVFcWwNVIplMwYOkdPH11YDv67wwsJRlPhVh1mZ7RYJmTYyObA4wILN
P77MUsy8uiyvPXC5j/U7KpuH3/VIIjmXji/hlI2FjhGKtELkdh/W0Ui0WJ+sLN8ej9A+CbEoKj0v
7IiQ60d1FmLam3Obfzy52vQnd/kRT1UhZ4q0A7z2prxUdkWSoEfUQTJU9D6oCWvtTWPJRgXwk4Hy
k6Br94juHSFlcj0GtkyOzcFTsRjCod5pKxU3ZjUS6WubQYLT8LhccgUtfL0xvi4wV6bz3rDrlTnf
vYwFu3+WMST/xM6kYIiW+IuG32Zt5mYfPv1H/FNVaRhtwRZKpvOB58OgbHyvCkZvTvBeVnzFhRZ/
YwXxBG3KQ40n2xsgzoWM6u7KJWaz3YVX5Y8ADUmJemESjKo0wwbv6GoeeUiBTTNHLWalPsJ4Ghgi
swqe6Y6Kg4E1FrvJAbJonwCYS3xgfUymCozHNpOX62ihy7PUUfHoAqhN9OhpXnF0QiCROfK2Rwzv
06eW9wMoVXh7TrWfpo8TosSQWhMdh3KHuF8dX6GhLbFUfGzXXSIiZU0SISwAyE4130mpi310A8yH
M6Ewe6Ge6ae8YjN9XS4WpQCKsq5SEG8Nz5G6E2VznddVeU2EFAQhNN72kLmMviD3z/Bjj53TDbPm
FehbbnmMwnMZDo3GJatHLFVcf+6YDOF5Wgt1BlIMCxLQwgtwO3IFwdO17kNhCt2WegN2S2aCRCoT
HKRfzid24KRyl4kxvmiPZKva3UX+o1irCX3I0S6ZiwfEacjMeN66lSThGu2ezPLWzVhGpAIRo3kP
/kxZZ72Rl+u9ruLy1o+M0/Sz+qXK+aolysLN1U3Nf1MEOIrk3a1Lffl9YFeO0qzSlVdfUSqAuMRA
23SA+kdRftxVLrMJ7pVHT4S8S6JOIpMoMONPMr/5ems4wMungznJ2OSIbGV1BBnrzLHijAKgmwiV
yiGne4EeA4ToRDwMl/tjePCGvcrKXrNW6ZC5VuF6MZkxb5XF6wli+Mr1s/cMYqQoUVOvoxUHeS1Z
dY/wyUhvxpb/BzMTzuSStTun18QPUZBvWwtyYeSUCQVRKeKXznjqDsZBx2hLRqx6jQqq3jRwqzEQ
gEQdwnTU0g1e4cCQc276rD23AEw59i0L6KsU1UrclJqW69SCUartDBB9ddDOPvnSOPDvNAxMJKHt
5LCq1jgfVtSbjpF2+btpd7FRB28mdHBEfdtlHwfNSpaHR+G3umqrprSNWfDkGh2CgZSwaPg12xTZ
a4LJ+ytCwKTzzOd41WAcNc/bmKpfRJ4AAPD1BcaL8pM6yra9JBq3g6hcrGmluBydy+aJj+GujKzY
iT/4GCBp+WMstfDRdMHXfLErTRXcso6XPrfw407HLk+3YEFR0HgNARqmr50WV/OhCHIkFuyGLxaH
h+cpHxBSjKrv//BOsMCj3mMnj1cFW4QD3Vxf2CN8NFJkraQPIZGB8Oml9U6rKD1cr2FhA1rxSvYt
vIoc+FcM4g8l/Wi2W7/ZGUCfog/O+a8ADTeu973Apu/0qNsttOzplM52SRviLU2++uq3dzj7OHQ4
UmHLRsBFlckDSs46xhwfbj5QkkFDadMe9atU//PwV3nF2xW7PkCa8zkd224QlAlfPv+a4N5XolEK
doKmKxe2Z4OwXpNYGgb6lyzDMGdwWpS3K+1ykoLOCcjPMZEuWmax2IyZZnmNTNyotO8T2neNYbcO
4mXJSdyvJ3SvtTBwneFnoxkosqzn9ThZ2+SvRxtwLqKC1ZNJUzxZuhkgodipe0nnf+ZRNKygTaIC
k9iJoa0Lim3z8xLBFS0+AHgVXR48xJJB71DpDX+iRwAnOKiZ+gYEICuIVtvkOb9HHNsKencLpCXc
WWAw0MRPGV3k0MyYapFPSdubgYu0YUIGOeWHsmh4CWxCdtgx0Sx3UGCdN+LxDuCy4zvok7L9xr75
cVjga6IEd6dBZNV8v1efX6hJ+97WCI/IaQfhuknCaJl3AnXIGlevKZ5/TDfEWvKepTKCddtGYIM0
6nZzzBTGy1vNSod+WZNk1B2VREqWD3IatAE2oOrV7Qj3tJyyQXh0xtKY8789TBy+qHSAXp8fMYsw
KyjmUc85Y+XVJg2/Ps6yE5olMrIZ6mHGXS+cN60kWNluJEBKX49kd3cMRVWdOQIWKLLkh+OjGzNb
nxG7Osle/7lJ18xXbmq0LSQTFFNvf9IMtNZVV+70wG2JmKtFJqqovHJleqv4wvvQcOlQ2ngDL63W
25L9/FuzaojpZD0zFMui9utboJLvu99R7KLD/R/DNmoVn4VeMS6I+BwxzuvkTraVDMdmaYUBMpQ2
nMA5BsNdNqzUhXpfLM/+MY0JLeck6AVBx6SJ0o9ZcawzgbOdAnxL9ZcYM2rIzD2lePZ2OrQ7IzZD
JtrnVMMRam1hm+IGYzga/1DlhTf7WyWRDlUQb/iTdpzC7ZUix8gRWC/Wh4v0G+gVvUP8ihJy6JqJ
F80m8zs2H1kyfqaMkq/pELca841uP53YSVCR5YX3tynLjRzs24GtCk0oysv2+79Ws4H1u1a0j0Cm
d8aNagM0yCcTfcqK2TRrkq51SFCsrDbeTjhBabcdoqew7dS02rpP0HBS86sfoe9x0HKvAEJxLAni
IorcSo0jGvhdfGed7DY+qChTx0nMP0ZeILPi0oSDzEgfgMT0lmMC6jyHEsCYs1odjswrKyajzv9i
ZR7N2o9qWx4q/DWTCjrmtpcjFfdtoImJGYudYfHxM1K6Xgsj5XrIlfLFB1IQB/vPOlOmjQ0B2ebA
6HOYMLKVqipDoTpAcIIy1VaU10ZmiyXh3XgBu9Llvh7mnF7/rlmpciTV4eozVlGjq70aomVD6BdW
J2wpCCgQQoxjaE8wwttzRGffLA40DB6T1JaC/qiqQkLhasMP6G66uOHYjhRv9uII2ksotAS90svd
5Vu7xgUVnc9EgZd7YiQIX/eSjAnB5QNmfQCVje4YbPIVHAfd4XbwoihBvYlweACj+yk5zZa03OxC
RFFmnAhIeoFdgsiPSUi5PyYsWcdRMzveLVUHC4YgAgZrNMx6KFWh50kDOJ5xMhqFktvtfBuVrCjR
vNZxVnqPa5qLoJeuG5bEaKTZVO1mzu42ovXESXAbOqFdHap/r4HZqCIraQ7svffYAcXJ7YudNn/r
YFZUANvbua3JMycQJ5K+rannKa+bsszV7re6UVWLhEGJYsFKy+RopmyAwIqmCgTqmqtHEU3x/r6u
2o95H3gGv0Hlq508yshjDuHGSmj3iRCGwQN401WAIywlforN4SttszjJ+gVoBhdmokg8fe8/9qra
wo53bCAAZcm9rCCSwwKTaw3o5/Ua+OHouxlzzsCNj4du5zdXTZGn3YdFmnUrC9GCP9lp34uuRc0f
J4NhhbR8tl93bm+QwPg5uZClI77jF7tXnb17sjvdE7pJw/U3m9T0dduoFCK6U7gcnZJReo2R3hdk
oTUxuTfa1DCv9QcwzkHr/IbRPTYEz2fXkbnQCYlr/uTnnmaM1/TL76LPRS+i7eu/X2RiKlTluQqV
A7r+JsJahbJZ6afRw0kobA/OPCERm9Qq/IFV5aB+5HA8OnfAzp2mmWfVdMleLUVnO4ylQQS9RQl3
0YV0x0s2DLZfi0IBSKEYwLks1H3FTy6BqX5GENssOKFq+/IGXzRJWvhxyfafWeMBZJA/MicIFi8Z
04V0LD4oQdgj+BkB8XZAQMYFWqxsuc9R8ZVT0F1q1mP09Z2wk8wO0vaa/JM5+RkydofYsjnsW0os
YaZ4HQUovAwOP4Xe+54lQM7uoVDGbs1nj3RfE5eSKgliBNWIZUQa62yMUeaBAgjGyfpVSBhGU1H0
Nqaa+hql1D9jfJ9Ve4T2PudHj8KrZsgxcWG+Vdvz7LW/uB/AkO8ZGwYndioqDOu7K2EQ5kgWKovj
FDm2jUu74m76gnasZ3gM1Po5elikMJSz6NjJvkx7z1qnWC/uL/p3e6UppaIqoQpH4ZWkK6ADByay
d/5npalQ1c9ouphsVbdVtqSTBxgvNbZ0HzLUwky6KJQOa6Bg3fvWd7o6txg3+2DYVolhpPp6dnw3
MYdxOoaC/6uVGKrSlif01RCwBpnd90S1nG5q9/80gzRwzG8nk2jbt6x69KTd4KGZrcT1U3FyxQDa
0DbJa8HyGsbk9jJrfazbqzwenh0sXzomWl7Ng3KDwpFMfZBLiEkDFebLtNVJtprLNXV1IhiwWmMz
Jkka3jQl8zwwDCxfLaUsvV60nt+j8+hkZIkrNuTto0daNl5Oq2XXZvz6FTPGORvk421zcr3BYgET
leGjF8nfoVygb7Mhs2jBHRGrvh53oBgIczMTnujWRbid4OKpkfUWQY21Cw5LL+h1JMHdcDxRC69K
gC0KsRztX8PZSwRFejhuXwSFI/OOg/mfIOSLHYlNnhooNIu5Ne78kTtgjbhkRIY1RWQ0IY0urSZV
L/9IO+zR7SbFuJI+oCiyd7+tVfJFtYM7GpSXeAAz1YVt0/BGxexRfzYvauxN3drLlP1EXh87BN4W
U24yk85MQqMWeKsnGG1mGZSHeOXNDW3pW79nOlx7CiNwBPOJWjHI16J4zaLjz6j3SlabLaCmYmpZ
mSNcOrBrZfcxeNQh2BU7eClTwbC2y4UAgwqO5FGkbzk0JJZ3oeypq+aWCKhCg+FQM8cL/SjQJbKK
J2ZR+iZKR7KoofOUO7b55Im8h4wIXVgMGCk6s/sX+kShVdkEMECLaeDD4dtYc7mhnYNWDJurws5t
PrHtKXTGYB/6fs1BQwwlGyHd/HbL1F+d5dOcpOTc7gCzXDV4ds9ezxdeOW3++edvSudmmSIc2Frd
4bXCGzcc6rJD/iD29rstW1Fou6r/xMJyiH8gF7SOnolgERe9pMgoQugQT+tcUp618387LFqwXt7Z
pmVRldS6ZyxS89HRydwE6UHQtp/iC7e+1yRGlOfNnVNQL+kSiolG4fEF+k9Y+EftXfczDJQXSY8E
Is7/caKZK5prrT6qmZhH3mPVbvZg8DC0U6XOJ5lX0+BdYmiHaWgVJW3q/AVmMF+10ijIUjM6nN6G
fXNnHdpndEU/p+dcZgqYeJzdXkJGrzO+vDgEnhzo+Um6tQFiSudZxp1ISzdA+Zq9S2exki/e+wJk
8RRj6/h2fnloTCXTJtmkgV6fwizwb63snXrSbsRR1J/8IT3rM7vV/9Tf6ymqUBjvR5OTGblF9MuZ
H6D7ji9KOP+p+qGw0He4f/+g4gdFaikW1MgdxSEkWabViPsL9kMSbTBvrMZhWwxHpMhp3M8Ez9cp
EEjc1iLYuL0RnfENvTLKc99xY5oM0ziXWcSpIT5W77dkicsbALdUff355E2H1wn/M6TUEELO8rKv
tCBcs44hcHuDX2G23DFW/u9Gbk5X0Mq84XwHo24K87zVT4piCa+nxd/orkYM7OOBfHtSHKGoRUsU
SR5ZQnX3SNVTJs5/ddlpzOvzDsdbFQNjJ6KtnuCrGRv61YNOm5NZb+nNQAh+M9G5CxLxZouLo8CO
mbnnEoNui0Kn8I9P2JBSaYULhIH4ZpyUayPm/wfmgwWciLFzvFReCclQU6EOv6P1jjcsgrq7LkPr
hktTmMzmXSwXPWJzp7qKcQV35sSWA4p5fbiE4oOL3o+Jey41eKgngOaopWmcK1GDTcKhRsrOfhjT
3m0JP/LX7B4FW85S2s+vxi5NQhdg+s/9ARte6NkACOMW4cm5cFAILTbHvywR5kPeP4Zts39/Fn3q
f2tRY7aePWiwCmAWyyX1Th0GPXetzL+6yOaV3jybpc+Lg5PcxOdUFrq/CRY2ytkDaZWluPQOJeqY
Ci9bZlZ8AcCg/bvO7Xbb9ovcdUSuf6pYNyZ4GrpJExJnM8ygB7HCoLoXWMgvKF90joCEhM4cpVwv
+y6iNDI97rpu+B8J4wf/J3kSdFEqj2qjL6mtK5PSIOuWgiiscNKkeHbqmfPmMnUnY3DS1QXJlWs6
XHnEt9uw63MtwFoFE+mWvVMr4mWGWiOsVif1pPU1jKHplu7RhqbJanfo4bBA2xFR4yRDeaoUiO7F
SJuHmTZSXhi1iRpTi7oc55/taCpQiZg+bGqEIIXZjy9mPcKTya+YRpxbh3h8CCRAqoAqqJTNHAeC
kCTzmLwoK4B3z9UCX5fqg8IH0Ff5kwBNsD4G+nnHL0slI1PjADUHBpJ6KiLtXvPiDH/D8Ne5k1Px
892AFB6G7yhdcJOf3EDF2sM1jMuf2d5wb2dp2h+nL+ruOBLCjfsXzIpXhi52Y9TT0WkNixXIkYA4
Ban0KZg4VgggVyllQ83GEJymqYVd8CH/YwOyABJ5wcnR1Vgc+6dCHTBggD3gbPlavHqr5MmoKmcX
GwcYB9TNbllYiJSWn7NBMnZlIbuIY2B5Yy6Hdof+NoO8DkJBaYJIr6GB3d59Jh/nk58axhqryrIM
oUB6kNk7xmtK69I6QPtnUKNMzN3ih0rsFKrsdJCQmQidEwPTdKWaUDd7gDd3Nmz5luvaIf1wbIie
WuAEb1c1On3LorM3iATRH6jEW1NFjr/gDT32qG57ZKYFK1L7cAqZpicZ5/0JUsspam/G2YVwhG9S
JPZ8N5zZyvAqSMM6VqEFBVzjPWLuM4+Ko1nn7G4YOBw6t8PSEeHJZjA7/Lz6YrUGqKiWev/wLBcG
WB6fmcFP1AQvwCP3Y2P4QdmZ7rebO3VOWrHn1LlzZHeJlub2d0fldP/qsXZq6VFQwq/+3SZsU7Ma
4cOoe3rSBsXzyn4MitJ8v7RxcsPLMdWxuRCFnHcZGsD1IyoATyrH47+GbI+akuIuywzpNffWdE7d
ldJ+Au97NMW5youLFqnygs4zjgw+iSn4sGQeLz1KqwNtvqNy2c3s3fwVTYgReCxNCZ/n0oaCUwal
Bwh7R24d2goNGso2m95P0oz2avlFo1YqG8VnDK/OoE+HYMfqHs+PVeuBrvVsWvfS9pxGMRy9QU/N
eGfDu4E+mHcOTNrt9gAvLF9BjnFBIWcObl1GDuvgquxZWaNIpeyBD8vmxNNZwZYTFkjLmPwzezLW
mKo6I6BRECjl3o63X5CjZgwIcmYXV0WECABr1xE9DExuWkEipQf6LCRPmPKjqDUA0wxn1h6i4VFk
MQok+XoBfgMCjdbCb/khF3/cAQbq+xg+QH2v0FHgmZvygNinqm/a9OtRe1NNCsiuXJRN5sZ1AhTC
e6w2hiE7+wzs2BiYWS0rnajtHdXpXs3Ydbndoc8ZnCF9NXnWEfuoVZgEYJ2WzzY777sXpPgr5JGw
rSZiTEFgK9LJd/giO1zcI3Djr8srESlBJ8ArDyhVOtGanmGucafDnprYuWiyIcBGqpDa+1MUpK+l
F6GeD25kkbfF1AKNR1GenRA5YW/3VR4h8gjAEvJP457NPdgM7fkdh4KYNcFC1APFXXP4P/TWicmR
G3xgj4fgtIs2E/vQj/vQ6j/W19ZSYeIT4Qf8xkeXvuI5QhN+d+QPIBNZpuXkCh/1xj3I2ovA1pA/
bovKgEFXRDH6uIMVaCOAISZNUoHV+wAMNIRt3suU1dJreebUtgpjpOxbabSARuReoh7eh/E1uGAm
FP/fLGrh3kVRE6o4q/mLDX4i6ZNwBbq5CVvlsafU80tb4FqrFddp33BzeLpdQ5VUikzIeokram/i
Q1WbrbeLq09o2sYYX4mslyYnu3YE0VIkdTJre0mGux4G4WeSplUF/wHpyXUU3Nd5sFIFHMF/t/0B
88UWCjJG+kHsk+GPcev7pMfoqRHqpEUFtB+eUcW5GRkyyV7jESRndlzdHXwyKjzQleAYaDke9Kwp
CkjRQMZV0/EaT8zS3INtQ9fKSoksf7JER9mI85wav3q2DWn5RjRPLW0kVJJa1Z+2DRhHzRBgkJxP
oo2/UlD4J0DpvIiqh8+LXqgRb7dj6xw1gYUYFieJ97TLsVGrdPq//b6YMmIxINcCA1VoUyF7DG67
qnA+SSRguElq1YQmRmoyG2VMl0obL6reOIp7aj7t0/lZzWYy3UFjsB1bYEK++uW4bkAaxqV0iWxQ
ZXz1F1ZMmuxPtIZ4jKJLQ7Ij73JoTfjaWPtyiUAe8BTiMHOHaxQAxOTnIJqhLcVEAv+B7JPmKE10
hxpWCZ7rQZDYWu1GTnS3hUZ1S+o4xAZ3MXfFdFD+ZTKA4Gj3KJwE4r0YpsJV9rVLvEQfJZ6NX61E
rBoAHicytaahhkdac0fuU/QgwdhRPe6mqhnZbMzn0IgPdmkxdo2qSlEGS4olrynyzLX2yFZ7Xm6t
7WcDIG7nMht8hrIa8GpqJ3iVzgWv7p921xNr66P5AYo0iiqMV3mahhKE/enf6o8Cy6aT4NSnSlS5
TaZC5EUa4884S9BVLVGgWMX3VFdZEwJju4p9JYqgDVxLoGD6i8BfMwheSRREcQ+SfGuHj+i2cwIG
09ukH1UxIdmI2dy5YyQ7NrJZCRViUqomQiD/wwf4LtO2btPARS62BHbVThb4uYCjrZe8mt7aePeQ
hbGAx2rx3pDbGaZe7mMl10g+/YrpW5Tr0gImBnPZdfo56E1dTKm7LgPSWdvjB0rv5PuKCleAHiyZ
a3xpkVVqkz0gBz+V/i0VlMAOg/cNEu81RYiCduflpmZwTlSgq9zEhQzvmq5nFx9GgR4BD0XGhBhU
0dAJlYQeQ7VxjYNB9k5l2vdDpa998r9MyCsP7UcB3YhT628U0Dd+yKQtEAWcSVx1Crsot/38OjwJ
9xBzt73oFLn7irWcs/Q2B+sGtPfIEoYZDubrlVT233jv34keU7DPcajUo3rwxYTXdwKwXT88c5Jf
yA4jGuov6xo1HkA/YGQbRJfjAZei9Y1sgpyeFEJHX9HlfP4dFnRWZ4WQCijplnDF37hFhF38sf9q
VgzFfNY84e9X7pj7wjxdmh0+fy6CjD8KERu/tY+zbLZLJW1gR7aoKgYJc2eCZUHw7a8cqqBe6cms
VitxAy1/y0yVZismeDrzWVlyRBXwJ894+3wnwdwki0GzQhZGF0ykPYBlWbvIkaoOEHUNEgwD34zO
5I6wWg7cvAnsMfe2rrX3c7lL7clcGlc6OctLrBAszQZYyDtAeAPcuZ0GLpOoevktobtaMl2f0kNP
KdFvx65nn13w0gY4iAGgBPew7+OJBo6JkhfO1lT1lNc/+O9ZzWrv5c3sSvyCwRAudX8Yq0VVmT8W
nXU4uEJ6+Y3S/dgALK9+bN3aF6VqANW08dV59wCmYTIqcbr8verUPGy88QIRPCKIrKl3Cnzj38a+
nREUOj2SQeWURuSfvfsjaFO3npZA64NfP3uUfh1jLf//cZipP2wUKSirFxDX4CVzxfwd1EzoSKuJ
7pOdCmXkjJeGTIXBGHB9ur00814xkNiHhPABA3GkJIvHXvBYPU+O4qLGc/dycK/cZ6MCZvCKGLAr
S/u0y3/+A2WO56MWY/CsG+tpxxeJLBjyZRgfvOgih3o70IjoWx0lIXINLdIm3b8VjS2eybIU5VDh
Z3Abz5S8Fd8+e7jtMVm9XRPfnYmjaBm4qwb2cVnb9ap9BestQhUVbidVtLkxIBC2dJshf7wcTX2l
Nlh35g4t8EJckRDLn9+Lc/1WPClyGeWUpKwz2hFMZnSxezq92hSj2Z7OIpkXBJ0/X0Liw8KjYRDm
3wz3iMu3vxRxIX/5SmAShjU6kmAmjtjhH6GSDGytP+R+aNE1sF8rC9t8yZl60b7Sw37YB/ru3Akr
bU8Hen2UXfGeFUDWwvd+vi85LGnKPdT8tHANfoikKAlMS+W5TcWHtk+HfXwWxzEfiCFteVhyObRN
dPovPeiCwK9rvL+K7CgnbLVkTyCumbFpDvVGUAmojUPbf4LR2WEup0LUm1BJJDrXaDqIdQdjL73b
t7ZmBbB7ZDqfmTZ7EQ4LcvCRh+RQ2K256z75Z14QbCZrp+CNs5OZ29Rr/zwmnAJ+33bQMQ8uDSM7
hTMQRnF9fx/854szHp7YtkHAn1+uds6NUl5SgQM2peEwmAhhg/zoUBkPXUqsOeauUzdeb664viQB
LVYwDzeJMmznYqtPzNV4tWkJppQ30KvyGZIbu7N0b5lGqXxeZmI6P4gzml2jfQBvNvLsZIBJUcER
39DyxyIRcoEzlDc15LF2iPhZ3VbZ1iiSLhJHQ3NPiO+zdTnOhRuYT+hWK8pLx5YZ/ucPcvkENNH5
L3X2rrM7h2tG9hrKJzgZM3osiXclfX7ixWKKajACMG+nIO3x1JEDqzSe/MQRhm7t41bisgotMLhK
qJ9eNlHHiNh/QrTUekoB2dQWanXVqWWoc1Jl0abVzz09xEaEjCXK3tZtJ9C9NmL3bhbTwPUXk1zL
b3OsdjhytMs0UUcFBk4W7uF0/7DoWGUMiw7ZMri93V7NxTMGEe4eY+dHnTDMxGWQrJAtHwlIxygw
9BugZbUNESdUPZdEzU7iLwhtVaD5R6bS9ZH+2JnKqKFI6R9TW04Z6t30xmv+DcyvFs00f8z/bTNu
AOl0sXntSCKQfK6A/07NQPESzQ+OKqkRc9wPxqku/VaOUx2B47GRXGlezDUmKMNbOEGs3DFYmSZU
pYnccQeZrJVVG6pwkH7PDrGY3Ww0v0Wwu4r9ENOCnkeoyYR6jN71ICnWzhkaqzytApsn2y1Hs6AS
ZH7JmH81+geqWj+HRYnla/oz3OKcFxv3nWN4ubklE/5HpWu7eZJTgHer3hxy7os5iAz+xaauA6So
K5nMja3E5QHbHl5HNgivAqRqli45b9sauV2Axkn/oVce6LjRJhpdYPMSCvFotAHhyQyqQfOwGuW5
TMMrhRJHpgeRRjAJsGY2xt6MuO84GgW8om+flNsY2SJdPYjquW5XPs86rD1djGwf2ebUCFmW6gr6
pkJkPc9+8pJUANNHawhe953HNbf1+pWZzPOQr7GPFho5nXLYbmEhFZpx8VCbMufAgpKPLjZiDjSi
r1dOy21Ru4mskbtvCAQzHxKfW/cFYiE87g5g4m5dO7XLpO+igknuYVBGZrsbdNYgRwZ0Q9OMq8uP
JOXC5rLpZqLek7/ovJSTBSQ1qzLR8tE+r+7FG1WYdHZpqmiBq2DQZgIdfgXWYWi3RaCmyPVzBvq/
YdtGzn39KLLcVw4mMkCQkYlNQnCEgKh3viFbR4gN3VDsMhEn6Vy2g+TZ9d6rDMO7YTSIDY7YgLuQ
jg3wYRETDpRCWMGDzn3aU5no4N/ZUogJA2oS7/kGUEjWmjkzRsXsm9AshrvHAQ5IAP+gqDf3+cAs
QvlFEAOeUPX1nuD9dk8mW0gvfzo70EjxrdLQQQI28OYkweY+TRjF58kkKe9XC4EGS1dhpH1vHODa
JjqxZYQo5zAvrNdOeyayNTVJU+7ClC/olht/gd5c6qUQoN2It0N/I1LYXfnjUGLi7UU6wavnirZR
hu8pFN1NGvkP0KCufGACUaqIhvqNlJHijUtAag/END8l80i35LQL/tCLp3GjKbM++qSqNlAqPOh7
UONKsP9bs4OX2sOIxcB2r1zYv7neapgAKshYiYqq8HuNPpIKJQ/+AzkQRwNcTCUcQ1CUpiHn8UC9
3854PtKW5kdLEkFpHSKNlZLu4lMB+gz8E2k6KWidNzvQ1LOikw7OqjoQVNbIHUUcSSWVXJqcKBcG
xvq6OhrIktJs3s21E2GJ4yIqcHsMun7nzPRDOgnaX4UxkOomDDRWBT9ISf2nNglWY8bj0mWpod8F
KWb8yLM/MoABKdJ5DeNngNkIQwleruVILi0OeH4GsGwzpwtOe2WFgXLUuYCRQDAv2oXgOp+jIKEO
VKJwYmu4TExcu4JCI2cXaIR6tH+A409I6QvTdHW7BDfODWHDM3DNyEAwf4NGB4UD2De+2qxxkAPD
+9oGBYr2nCjskh7OBYdoo0f8HMUufJ3gkw5i9qtlsuBwpzJsyBBZ4Rfnk5jCtlCp97TL4ltURuXe
XXLd9BZnm3B9l2TiwqwP7eNTcA3XvQwj0PpVgoUPcVhqCz8g+QSVTr4jMyaKxI865W0aJjOqKD9m
r80p6P0cyoU9Ks4ASs4h1oAKC6SaaLZkCsK4sp1nyBQR8PIB4aUOuuefhZSTQUA30N84PC8DQMKj
f04DPf3ag6wK3VEYeMbtfJyV0cMiYdWOPafk4M18JX0tUnRUyeKuolU/m2jBc/BZ47PXx1UWGzdB
kGOZaCrvVfdlNHe8uMAhqZUUfh0MuGsX+SnDgPW+XMTuq7CJNH1JssK6U7wcbgmU4pDSPo+gvHmX
yYpR8ArqtwTxVoojrKuXuIrd5RpR+Jn43bO1qNCj5pPloLD7IcBipIcDiu45dqi8nkmVOti6F21Z
/nNdBXZEg9vkkSE5lmmA9A8urhDhZp1TLyfspt+O9SbIveHt2dWWxTflKNlQT7q3SflNhPbbzNNs
VIS0vR40/c51f0335TjrMopyn9W4cNF1Fxygg8Nz7s5htqLmDD4wl1EvTEJuX5JohII1C233lhoR
Dn9kGu0LVQuqS2O/ZjwruYajNAhHa4NRt3IvtN9cuCSsoMkaZeZxB79zuuz0XnSc/kAXWit6KD8O
6swNX4Z9cQcyAxCSy2EOVeBH+7+o6toXjVFakjazz+Wwjbfa50T4mDpMxYRXECo4UHu794vcqr5V
C2oW28hraMesdvoCM1JwrdowlcfcQaHc2TFRyDHMMeeVg1v7BKvqCh3LeFy6xCxIqruyoFcsWxDL
293Od9HXR9zjtwfO+aWNJgGjnXwgdY3/8CP/Bcw7Em2bJBQAw0zpQKJTSPEiYR2M3/BGB/DlgfKJ
cS3F+R9snIRRjAUoKNbA8aDoI6hwHImCpzmsUjC7bDLexxrAGMSPzf3ghaF1phVYC2dfnndCviWk
QgDbi/fD3shvB1ipD9KoNeBJhzBoEa9XxFNfqPZihl4hY/Pdm+KhpQrEmD2JnuoNTszI6++Lzmn5
uiaKUsi4qB8hwNgBBflI2bmAedcSS3hTeX1jz1O5qd6PPvckTbrmuLB66c+C8kHQgzk9O4c3hlLJ
70Sj1v+mNWUaQCT3Cd8pnniIdzKfFVVwpbxHmH6h8UCqejDk3znzWl1ZnMbf4twhDdbjwiYPACr0
/MQtWvP+gCZp+t1Dr+nAm1BiDjZEx1zNlWZA1iq4OhO32wjeaJpVzb3O+TojubbypomKzCqj4RgF
2f9kJkvmBlXH4P0iNF4fstvoMNQpUrwA+ZOCq21VX0S4DX3VLPnPJ1DgSMeGMNtjoXHZa+lr8w9j
o2t7s/zMaV6RcYABQ++niusZUx/feIlw7Jy59qWM+ZtkhKR3JE7qlAsYgVbElDIYNEo/LX8wUvdr
cxmTciHMT5BcfmSWcXoOsem2zlUg75zOZuEvvovQadVhikuR19C0304BdRzEGXRQv1BkiS6vomRy
k+F2Zu4y7nEVgwf75+vGhZlFNFapfJhH6W7EldySNooA5VmICyOdVqj68nRvbFj5f3qT8mFn6Wec
nhAB4/KTbxQJUocbTOfWhCtqJABzCXMQfyy4aSaiXr6STh2uIZc1U9Ap4kbLyG3GpyW7YFR1SqAH
dLT9DQoB9xyNlSSj7H3IO+qSojSZzK6Y0gUDn6xUsM1mmyai8yrTZUODbyL1PiU5O7av1dPFbLdF
OCEcb4QzBANmWovENFLsXDHvFuf+0seyv+x8MKYRCAqkK1YnkPV7auDjRsCbiI3qasqHhvPd4uhk
Mbar5QdkCKidYZcjy6biSv3i8QqqhyEkMF+n34j2R4PXie88MEXNiZvsTJOfCxspB3S3OdHo88In
55fp0QM23zs28j4MvM8hCdreVqUr4iiSDC0BmDHs5YmCSpAX5rtzPq9hzq0gsGLgCczNtTuGRlYg
hSsWcjcGIp2s10v8RrN7h7MmbupwulC65mi4yE8hDuuzgfa0qrHaU2Kvn+fOQ5guHQCWsmTa82bl
+wSudjmlRV0Yyae4RfGgki2YvVVrj1uDf4Pyxlm0hBa6EZ1KcITJImS9DA1BKeGeC5W2FqxCuc9t
kBrrmIPLL5lOuuc7TTG+UTaOleFyJ4wKIp+aDhwwVU50HdoSv4Bna1J4+lU92dM1fhROtmPYOnmQ
KKWQ/1sE4QqQt7U1b1jh7TXJF8i4dg+OxnofeliUmn3xSJ7sF0G/pRnFDwxXSOslI5W6DnMTTUWd
U2FYt3/WkC1+NeI6fnd5cbvRj2O70HveDuoFuj6uOk97ge7ym3Sj9mrm/BoHrRZXT+yjPCkreHcs
z6pAWPzEXIRawdcnDq/KGw7aKKQ9VrPfRo6H7royqkzhfOssEM5gzZXU+BagnedTfo4KS/xdMpJf
o3QVjBGxEh8sOpCSy4/GcXXEcHV7VzgMxMhHv1KVXBUTsmma1A7abQeH2FRTUTLOjVjEHK7jXrRa
1zssKus+GrzPCc983U1a9LY2QVTMk8/TlrFDg4JMNtG9GAAzi4Rxq9yc0whtGzabo9qaIZ1l94q8
3ACb/fGDnqpZvsMizuwzJj8p2xvcPVEpwVF1j4JiQOl336ds/Sk4JDK/5RzWdxyaEOp3AH1trS8X
AV3RoXOg/GoWsM1TS4cHDUPiK1HEb17Sc6TfwusU07BhfFS4nMlgBUexZZXQDo/3oR2kswoNbIEi
9CI/2SCvWXBxswlcH3E84Ab+OI0ZBMFJjRFj8Y1MM7V2AHTN3L4acNIxbwmhwoVwQCPP4hrGGVF0
5bFwQH29UZKgxUn9iL107nRfeetsWEWko8Bh+sMnINw5dwm9x291K2rf+gY0YEkDhsFxgLstV6YC
jRf6mDPZSRYT/JOjtpufTb4w7Tbnxq1w7hrW2YTdpu/bV47cx3Dd5jWGEIx4AJ8WCFLb3pEkbpl6
+5juBny1D7X19iwF7Cpzqy797tP/5p7lDQZuJO0QsAwfpQEdjWbgpQrvMRifZOTaUgzhJpxBzWaw
ChLJ1P/0gcycrRMig4xuB4+P7n2kmmY7YRk/j+JYdD209XeaXpTXLPtw6PShmTBi8lbwH28qMYSH
qZYOKPrCiBdeuADpHjX/uMYoeDHbQgLo0EihM8uZdvbOR9C2nPNJHPMptcpoWa+S1scy3gxyZNSw
vTLnU+M4Z9hN/Ra5fHUI+h500I/vER+bsgqfLd20qfLcg2YxZfCqgP18h93jnM4hgvmaF0ed5KRL
91rJYoRY5pK9OLIeknmVLIAGlriUjYRlHfpGzX+DX6Gva3NdVz9kzL0GFBRuJwxUbNLSeSAAlKZf
msuFUzXN2jQ+MnyoHheKx29JWscX5DW6iAeA5z0Vtnopm6n+rgxqpfI+mAJ+5O7exq8Hu/YfMmnH
EP7ZKp6Vy1s4+5Z4TPpgqat0kHhVweD5QGAucUO93Ric20hf+2rONP+sIMKvQbA9o4qNddtuA9hN
dYRA5VmrF/dhYAd4I8clVqfBkyTuEKzPt9pNxmG8TtMcUsHwCi4D3MW0Z1LAS8/fCB9BMomAdec2
7XbHDMVSa/X1uRZhS4/b2Gd1jSSWH3VQH7a7xdlsYG4KCxw91bvk8Gt0eWtt/z1rIyawj5FJzTnZ
IcWLEjIatsoMI6VuGswCHyUV8iKt4qHJveIyW588rEZLLZt+5cHe2pnFVX5GnyIA/1q0WvFUbq3P
S3QkV9Q74aHFO3t3mPnLOMdfIKPWUTJ8y3Gka6QLl/jQF1gRcfumQxbiyPs/8MD4wqLStpxfhEB0
0hsGxRvXLRpmdUdZN521FFpgTw2HhiACrYazik/+oEIIB98bN6zMxmaI2iNBBUEYHipxWEN7zpuO
+I3MUi3Jt1NMUriNMMx4RWNYu+ZFAvPJ7sEtiewKo4JRXsKEJO+RhaM7uAYHJjAF4jS/uFjN5yaT
aWnC1o4KGQPoIKkilhojLPM/FeL7OBoZm+HFJhNy7o9Z2PD/VmLYHYYMD8LXNcaeF+hlSLBIbBjl
X34NL34RkLIcPRKv1RgJBPaERlCHlCrVrav4yf3liZafsV1blkDZgQCkVznMvqggVfd5VV36JmVU
Kdw7xTx5S8KPLkFasnxZq+kipkA1/cQFHXLDJt7hGAtcJKNq61CwdBKFNbj0zbNqGlvHxvGzEZOS
OPR9wa1JXjgaOy7YkREDZ9EbT4QDfCsTkG0kyYg2D/k9LtxxX9OT6IAHJGTnQnZr8Dgt7c8QVLJc
rgFu0QK6I+DmcHub1sxCk8VIMJtT+v7TZRR4Yi02cUmMKm49fnSDAUccuj4BRQmIdN+92W3shiD4
cgwNaWNS8moUf70QW8kZ+bOKTHG0BZMfdqLcYy+eokiH7tncjfU8Mlzxx0urgsD8zvOrEw1yV/s2
4s6VKjT5GnPdG3QjQ3eMw6fnPnABxT/kDAI0GHgJonTYY/BlEzWBYrYaHZjmASlX4ywWzfiE9b6l
WPxtmuY/eR+DSiAmFMAEPjucO57r1xPIx8gbrJDLGGoRwMnuEOjCS+He7TpgM41Ol13lP1lO71xK
aCDi+ZAe/zqsULF3QXHqzx7h7whSJRS/zQsLLuj14JfhmNZiOmbWuEv41SwVh4C3rCsx7NZntpTH
7Ma9hKKE4ey3+65hdn5FWeYAy0kaaGt6wWpKzPpFjDUBCUSuWgPt5h8pMvlj75vebU/W6bvGLXkC
a1wsuH00I211sF4Sw2nd7FpilYpnpkehpbC8+n9WE88vRwc2uVTjXYsRiOXYyY6KTE4fSkc0tFzI
G8p7vGDXJXyat7SJYh0YiIQAL/w11vL12dS7yo5PuKDsFkh4CSwjnh+b5grnNu1FF/s5ooxLqE7W
087bLIUwEp7TJ4mnSpJ/S5wa9YjkadPtkRPHQdOeBUOK+qNhUHlaXQRHseEWq+Pu2+CbhV2TIEBE
o2RrrTjcQ9zwGe2EDSLkypEARPxjXAY8KDDE1XiYT0CIVbNjQO7fkLFvmJB+rl6XIukP2zKu3ktM
NGVVBueLF4IuAQBRguQF+Rs10LaGiJggR28wKuKpmtIAozxUkjDW4TapwGDszvhH4KMID5bysPGP
nzTpCYjQp0GKvgJt6eOwkLtc9Vbo5aPGz63BcEVLWNjJmXPCRUdOxC59pdQJgksDXFeugZcEh7Cx
i2Pxp0DMeHXU5HodFXUZ4lGzHR1QT8KK1GRvB1JWVVCct9PiUPg7Z1Akfp6S8/h7a8d15/Z5QAkv
GqAgi7Q65UXnOJWHoWbzTlt0y7dJ6Et+y8iut7sdT6G8utzqMkeQWdeKxbm/UrCM3D1izBHq+PnA
/U6UOzpbJ042/2KYumO6c4kCJni0Pj+1PG9QAFBl5BtE3+JcWTh3c7fIkVUfxoVEmx4uZiVhLnjD
7A5Xkqlf/qpIC3zqLD1n+R4yFL2+oqi7RxnfDtD4kbFRPzZqZXNpiAncR0e5U0r2r5fAeqOQHCOu
Zp3Lf3xm5mzJycgLF5Gq6vRrENOAo8IN9R4w2Pz2z7OJ6+i9DSFQRMeXwz7sHE1v+K+J1hu/N9BU
h89vonYRdj9GMgwbgXeVscCe/NMYzddjGpRw/vPqSpCTCMbED6jMceY7ZXKkfa1foRqmPcFknfqv
XYnx8cAgKk3Ls1dNbEbyQUgN8lzMKnXYnJwx5CD2u5rx8EXWWKZ+ejrQyMcJ/FCR6cOhBXscUsDI
eBvsbTcF6pOLw9vLXFHNwI08dOK+7U6Vc2S7l3AgFUz9Epp+fRnIDSdav7DuuvJLi8tQYkEGW7FT
m/x7xxkfxvuG6Xkse7hMbtaI1o8+tJmJ19FKHZXcOTc93VREeLrbymNGMtHaVs9CtjJfG9P6Dt+M
wKn76XV413dod+w9joaRkdkiaWb3SSGhuXcdMprxi3chqbXk4LT1cvzx76e2/zgg01fYuKBGgPcp
3fJ2UEFTzE7Ha2kF8EBKV9GvYGMBN5foeHb8fe6LB4l2v6sIBfnKeiEjgYfBab3ELoNkVuyugAdL
y2omyAT43CAoCtbJ5bcqN0me6X1EvOnknScR9BlnnCCXE/cZ1EuurS7kC/BD0KKXxM6uoHbezI0G
lAzvtk2muclGLKoH3AXIEw+ZfiOkEo7Ks6/ga3i2mj73xJVGU+P6eifGZTSnjHzah+L84zHNKyuJ
mCL0CObGss/7QJ5M38zS4vkub8IJW/MoL117dnywPz8VeikE9DuDoRi9qg2oCD9KeNuLaWlIMb4r
PTcxTwglble4WVglgxD9OWELnAf82BnSZuttqsEaLnk/S7PuwBPHyx83rC4V/3zuntVGhdMdoP6Q
980jGSAIXmB9XAL+bwrvnBjC2kqSuU78LH3jR1AdZUSA5jYOppjxsC790u/Gb8GTckrLPnq48tPG
YPK/rZhDjM1UG6bX0jZXIMzPB+FHgvrWl7gHVGSVIkLZOxDGc/RbbrxD+IlXyHKT3nw1pg3DjuPg
ucp9NS9XiwVzTs9qHmH9sFnFVhyWfTvUwFJE6glELQcJwOh3XCg8J5KDlui6GEQn3cNYWx956BFD
XE5Xfr5T6GtZv0KlbeAXQBtUNotLFH5gsZMAUixZfG6IqEnH6Ngvv1wVDl2gTeE2Go5adjLUXg7t
Z4c3FB6OvEkSgj6IknPPItFZT3huTzpTDJ8niJM6HgfSJbJprwrPsQQZyluF8t7ZVe2mgzM5N6Ha
nL7N5qMNita5za4yYyfvK43KdxnkyF5V3FHu+0Hg/rjBRBMLqf5eicpOipd3+VeGRsNF7iWYnLM1
uP2fqgYRSJdAoO805+dNtfqPjx2bIok1NKKcse+Bfe7qoTPQXUMuM1uqPKOelaLhGjWeh4vXc2kf
TyHlhVSGMYZXjxpomfPvuC+BlQ/+F2UnMjcO5BS90gTkK3sfpVjsiuO+OA2UDdNrJsoe16wuOnNP
zHwGGjifu1sPapLqaXXAJcSvFbm949NGnBZxw5XnUAc7G2wiYuSfT+poClgcPDt2RravmmT1Vpd3
8Ywzinwxks9vume7+CPwLdBS7DQSrMJXUAkFxfHDouSOiUPzMTJo3VFQ9w02Rcx5uN87DHPQv96q
1IVmRZL5MjNnfP8jtoRuxBEwSu2MfwZ2Mxs6vRIsvTAKQT6HJgi5+J7EDLsYafOui4ZlcZhJjbtM
6nYmT8tRKdJR1jE1vCbzpJ5C8AT0vPwpRzcD+bhQCE8f0qqohP/FDvHAAQ2W6+mEoK2RWNlQ/eIF
/4NSPpfEPzTk/0diQm32vMKn8kEWcfv8EmP16qgLLIgxdqUxpZjyu9Q0DMSuIYX1303NoBKHdOcm
Q8OcmmRwWX3K3dC64OHfSqDkdML4r5cifKiAPZhief00by5bnZye8rNG0gNx7H6euHrWiYdCdfy3
4LGljRx0o745gmNlSCuvGyPmhcgSpJzAzQltsaE6k/T7LmRQh4mcMkPFqYI2JJLAkLL7lMBhLOsR
6rIy+7lxEjXKH3VFHqaOBz++AyTBdkrYDf/LK2EWTKhjIw1qmBfTCpQ7sSyb+N1DZR+7kTgB7CY1
5N8Mvxr4QpH0TJY5AK3LbFn5RPP2SwZq65AGgsglUDjcX/P1o3l3mZvGc8QYcCaO2Socl9uXo2pn
nPGdFafRjET1qtAwY1D1W7yj3AfCYgKBatSpZzV9nUttZWtK3pOrkRXTFnTVabA+VEkCCYePmUJw
sCJYlZQCQnuxKxQWryiUuwgDDGTdR7nsqjNwHeYn2PsGcKB0I+/5yJR//z+s0UGE+d/m8FE1WYTO
hNm90zizKMBlyTgUAKsg6QfZ8jSckdaLmHi04GKQtsGU/VyM9QMg/tz97H3DdiDPDXhq6yrnRdV8
O2mmWt8RClaRBb54l8hos3saCkrH8hn68+0HuNodsF77ybaJlvsA1hfXuqPtuyJ+ohqRVUD6dgxh
QOBmaiG/OCSMRZyE/730sJJoKcPGU5wvhyzkOa0bPbW2rTWv1seoTch4i4G2jrwoirLkn27wooSj
2lpNNIjoaHWK+0R1ZMHGr/ATYykdE/aSoqTw2pNQitNXJWEaic04gYGHhiAp2A/is1QhdPbLKg+K
Yko09A+aygGrDMenER4CMEqwrpnvnChcUJJkrm7i53TRdbc4OZwOMOA4pefnzGONdKNsXTQwYM29
xk87jOYpbP6zXXnKvlyfqRCaTu5oaRhB1Gt80TmDcVHBAnDdInn/UdaYEG98LANANbVlickLeTc5
Dxn5tbCj081NEBD16TMYJoIUKWPARESa/TXmA+lD3OSEy50yAC2DEt9U0YhQB/D7tzJmh9yDRJlD
sJlIz46fN3WSVj+02xwcnZq/O6HjjGmKETLEtd7G2Txtcn+ZOf+QFp00/Z5/ybMFTV+Qd87hJ+T9
5ENA7Vt0I7eoWe2UqKeBamCbZC9x0a+IR6XlLznOkPhV442+RjlyYuQZjQhV0qFW95zdcLjc30AJ
b3NhOmsLvNWK6qDxZw/lDJfsHNDXQEfPxooK7ZI3nHIK34S+k4XzmOFF0d8AmiRzhV6Od7mJla8M
FvyWXwp1mtonmlcQHN4ojcJPJKzoKr/g8E5e6cSyTf7eMiNpcHv6jmJ6+AxJuGVEiCqQMMiRN0Or
Ecz+UJtZBZk+NCQrnvi7+3DQnmYRoMvJ7ssQcLJ4pO0Kc4OihOYlaF9PDBa0OPL7FaKiMUwS0/KR
oQdRHRCN/rz7AAdqOr60YR89pWMPPor4UbXhVIMUCLOAGV/nPjuPrBszLHid1eRZZanmpL/clEYH
qrdMtOBF/4k+SL7ubvAg8NMhS3yKGyUzbtsEHp+X0iBXq7FTlR8FjCtovvClsm0ciYYLWm29duSz
yVBmzJ8pcsqqqzb42C7Etno1f8tgSM3siuXd9TvEmNPgmH+sgG5iWFGoDWqqqn4ACpCdovOaiyRj
VqFw0mGb58cXEfNrtreE7riNKv44F0JEk/ru3ejNvYPc1d/tGjdAiHSduhZcU3plindLTlYxNZbP
zssHLQgDEnbOVY80+HooBtGOykPEacLZm6C6njxrTIytm649PgH461RAW/8rBCamEhu8btNqJ1xJ
1jgJdcp5dmNtQuSfMoouZdByx2MbT8j/ejA6lf9DfaCDGiMxK6UpSUcqlLc8PrizX70TxrUP6Zim
l+oufc+IuhhhP/G4od0viBmLOgJpOdTcEgtRCBaFpWkXVOMjRryLeyT/f5A0B07rS40UFtNPSxEu
aWvjRt60mHr5Gx2rsKjowBJDfaSKcSjZ8n/s6fmhi2zD6TEVUgeCYTFISQ9qmR/Lj2axPNZNJ5pi
/q5A+s+A5aHkHdZQ5lVETqzaRKx8YmY0sg4Sme51cx2MuXrxDyLIK7+zGsFJwtfnzuYp6yESMmZC
tTnOOtW2EsOzAHiCXYBRMLZ+LmtwDH5kQ1v33F0ifWzGquKB9dYjgWmerU/8esniRpq4mQ2nWoTp
cq1TgqN1DW+MKSDZGpLPF0nkPqYloZvfb44KlPqGA/B4rV2RJQJF+5PARmY2NqZ3iF9Y0fYL1KJA
jh8lLThUfT2qgmGiHM5gGSBxKCbloI5k02ld8T3qJrgR/x+nyNIBD09bjRgc6F7FHX1ICn1Z2R/E
loU8qWznRnuYvHydHNEq666vR8m4Rewmot6KJf40F+8uysqvsgZB2Jt431A1q2bAaSVps+l3HCq/
ta66GgcBrXcwVTFGKlagfUk+bJmHO+ApGdiSzB2vRgfNsLtYKwAEyS75eK9sWvfDcCE/qJ1Zp7F6
A5+qolHLpj/N4gkieyib2bzDWX6YyGJwzc3rWK36Vf6FctRD7J74SMKQCsTe6I8k8BOCeCy9FZUu
7IVzJLNRAeRMWJn/WzpPQyYVs6ialr+OtBrKCoMhnvmL5uC3LNXLtRG2m4+bxt8p3FadaFwfH0Fx
NZHIMCofPxFamRwJGb9P/oAniTg9X7FFO1D+hG0dBoOGf96sACAqmdNlQTMSnGL/wbY2VtfvTHp5
fXf3JblagC0zYWKMgUWRm1npgqBi70VVcrPBNInP7fcdehmhIEyQ/sylTGP2bbxYidyIWCMS7Fv0
npcwgDNr+/TU0B/wYAU0YW5O2QT4DaSWv3a48hrv+RuYMyC+wFAnC5ApkRRi4Hze5nORjXrTl08f
2KQYW/WooWpET82UKoxlflQzXo0jlYX6bB8YQdYAYfO8Vcvm6xJWx/oOszVNkxvXpdo7uBTR2g+D
aCGNn1+KznBK0ZQPNEXUkxlBq+AjQ7J9u2POwHwxsBu9FeRAG7KNd0Tj0PutEN1Rl3lGgrMnsR7G
VjeKWDFbydibpB89b1xyMTGYILD8CfiOb5dOTbhlMREw4gLF+DFtQkP9GqLIe/0NvkxCIAUsgBMb
NVOxJwIn7tp4XYaBvzofCai8MMAmPALVLxeGo+UPsZFwBx9FwesMu/+LIw8eoB/2GjgEQBYjcxH8
+UGoarUGWE+tkPiFRM4f3lhOi/IRMfs/MmGsihlybTem8s2AjBENyUSEd6TdnWjog1uiL+QjBs+g
BFrHvSiGsPCV8U9ktv09NChDcZJ1hHP64rVyDY2PwYs2hkJuQvUqNyly/GUo8HHewMUsD3AFJWli
B9+6BLA2zgMIDpMD6f54rUOsiX3UlBou/kTotqUMmShhJldV6HiEWH/os/BTtDNDntNv1EAem4nm
C9MplXEaEuZoOYdFmZZj96McH7x6s62fFMva69aBZ4ZZMcETDZRXxxPfk67SLgxxugmLWKPX8+KP
r4YUjDcNy/5+9HH5LqXOxrLpRJdFPsIul5Nhsvcpv4KKN28KWE+BwihNchPuy9ulMPL47KpsY4+2
WOllIorXchmyjwWuUbc6BfmkhV/bgvjaeKRNTXQlhJFxpqqPzWnWWpDKCmGY7XcnLK9+2F1C0oHB
5ehBqIQOPl3/AJKjtnPttFUqJvTsGNU5M+6ADJVXZoq+k4nTOrFvUXphmzXBOlieKSNcit2cSCZu
9j2pA3iSjz4emmMzgxDY1c/MsPbWO2/4Bio+48KjR9TwGFirmxTOXx6CnjJK5xExr9VdKJoO2E53
CRs3IqIMe+XdgefPnrtcC+QNaLFxUQ7m6g8BfU0SIQsAjBpN+s25QHEtnIdZmb4U42raQfrrHdQi
KjE/fR3nsXx2mIFklTh0pj1E2vMzsjUN2FlVHT6aPYtQoQnfolpI1TJcH1byqEAv2LdUt4Cof67w
xlGtR1inIpRVo5C8FaKJ2L7MQct8nHW/zdXxCIWXs891t3ns0KgdWIF8Cz8e1Xm8i6UUguNyuAqA
4xi4YHlCO7xqMex8AyMkdvbQZaQFAGEgizhFFVB9buArLrFU3HR370yybtTwnK7iGfl+hjX/SnQs
7wRa541k83n5ef0T0mGaqqFv63mwYS+jjRj9IGlGdZPaJN3S0U3I6RvXmGj8wlt6A86cGVRHZfTu
PfN1uNkmuEwR9FPsAOTNweNy7OabuxAJcbuh+r+QibQa8bpgXA1m0V0IIF7oEo4NEq6b1khLD6JL
BKI2YYTaHnSp9t8JxfcGVvYOC0hQSyFDZA6eVErhswRQ57PmGVkxz5Modse++jqj0+RqVPG/fPbA
RBai3eG6X4+PO+Qew0oJqyUToYOnvrAzUpuOp0fK/fSYVzhn6bajjfK8CMw7xbiTXk+tO6Qh3QJB
asQI654ESHLvZJBThP6XrxcSfCvkjQOFAOxwK9CQWo5fojrh/ZdsDAHjcdfgS3ybKhkbCA1b5ucu
nTKVVebd/U3CztENAoxdk/re/DTe/TprGiFhaE78T1cEUwwSyqUOY46xVrXANJsWMw6+Xbcbj4/u
nYWgoMePDyTXS/h83Cii9xUd7d9uAJ6FZ7xvztQH+SHQWyZx+O3VQSB86IOFHWjO3/PJioS1YBOA
IFFUuthLut688lQrClU67yZ9Ahy02Wz5C4slNh+vLBx2fAup4wBfXW6g58y1iOuoeQXRQQYqOc+Z
c7bcMfxp1cD/jzpnsRfo/4FCHVNjma47ZlLVLDAa7HVeOAXc4rmeU3fqMQd6Bi0N35P6cqHEIznz
Brl0n82CKO9FJSIib82RsXdH/u9aVoNUoYTIlNjZ0ZyaBhtTelRh0LpD8Bumf2sZd2PazncFkDOw
9WIqUW4SX7vPKLfkrwSUgX8cENTCFXKdf7HJRQZQZd1ElqfFCGiY50TXMDOkuZMSNzfsTOORKx8T
gl1k0uUxvl7W+viXoVh3xySB74kupX0XadmJQwOIZHDDWbrRMINSFe7g2VZqwDaknROfaXMurfZa
43nOkj6r4hd67GvqWLNE+YgN2yroO4xAxspjx/wg9PjGqCGzx1yRBjCDS7RYG38QqVl/SXxQY35c
Pm0BJpqmF7gD2H6/uxEdn2oNn6Xu/+cTLBi1NlLyOR20SFD+yguEm7Zxes1TKN++k+E3e93E0tjL
bsQNIrHl9fPFjVk/FUuMr+S6DSNKGZLenxXcvUDU0sXZ8W07kczLPdfh2lj5gd8QoY4LLvpt5kHq
dh+q2uTP5n0Y1eLvjfluiWlak+UWgKAXmUJLyaAqLfeNOCX+n3kvGIFuwpMgGAepAE/9ntv95yRV
4uowu24/8QpVZW4PZr0OdVbj7QYG75Sue7ttKmKOz5X8M8sJJ8i+k0JTs3x/K6Q88pbMKCWOvk84
gUQOd0EkoidqGLK4blafjCa2nkeeVAi4EmixEZ+MT2syIQOYd4Vhfsn58T6Y4yQbb2G5xA9gphZU
qhmHYt7YRO+WCwpu0RN0SHUmH3kDRKYWbSy2DiuNNPT35uPFlQD5W0ZK09OAfH6oNQahx9LfKN8H
zpOE29rm8U0+dJ0JyvipyjZ5VEYZZSl6jVek9DYGoixjVcgUhpUJ5PGZetKS/IxVRGRGNM8oYqd/
/bHhR0jueMJzEuGwh0M3CrU/c6Xgss4oEgL9k2nAvL0kkRD6FYZJQ4G5ac43wuhWtLkn7mS+IrxT
yVTi5cPCekNt1ZDbtv3pHP6en3jb4Zg/eFAbQ7UcXxErXz6dVUZ2YZP7ptJ+kpWWCNWA3Ec7VKEC
s+t1bfR9K6uwEFdj8y9iyhKVCOx61XXgmM0jVjZv3ScX5VG2P6WGQK/xwbch8z0u76en2tENrklw
eBYXZwxvWzsMEXnTtcfrvHYgu7xbTM4t8iJHBeajv7Lv3H+b7yDA92wviRqWqqxs4EOh6L0fWZZF
XbvTMLElxMA9571Ltdn8Ob/WkX5c0O9/Gb+rGWvTkEPhldyh5Ql0Rg3CEaXiFE+uMBrKz+KYB8Kk
UYXfOO5Y6JAj1EQXa3h18Yj3adD0YpAeCqH8D5pZqcxtrLxqJMaxOtDLUTlL4SF0XsLv2/AEs45Q
7teCUM936bFeqWl1k6LPj+Kzzk1SmHTkfBVpGPL5UlRhoheJca3QQarjInQqPk8WPUZ1gwtB28CY
WptUbYQkN4FxYU4sRdr4DiditPfZQT2fOTTHj7ww0NHX2HQ/JjDrdWnor36HZEMK3htNnKrNsFP8
CfC7y+m+ZALJCMOmgnqbFKQ7uV8lhTlrzYCBJ3VIhj3wF06QUj90rZmtxsoWBVCWT343wHJfhlxY
3eSSHNyisqmJI9qF6YY58YRvNMkx4UgM3ipqVqniQ3EPO91CXIuBej4XeUmperPJnCD8K375TduS
HXZqphNB9lvBjlFvRueY4mD1kkeBg1MA909Fa+cizKdDnLxVuHKrSKY8hiLayFOWcW7kI1PVzH7I
tY4cLlfYbBGjoFWdB2O12nXiCsxho4LtNzLv5uEPJsj8jUs9iBPs0w0oVfhMcnBNtNnX20L9peZ6
wQG0MN8ktdN3GPBSGe1m9o/aJarNxjluc7MW7fxhsTXGBJkZsT3J59/G+C3W29s6EDfBcGtgRbFQ
Gy6BT7OlHLmvXB3PdztRtLJN0P3od2wag+LmqSUvPTsGVdGSUEtLmldLNuXqUrMg+Ggd/rxDZrEW
H9c006nMV1o/cHcr8TyVqFXRFhalWx5lEuZPG8AZOTdg1qYPu4RooyZzjsoxcpbVmkH7h6rDz7f8
wzc1fF1+h5FHQHNpMMYj4yjUZXT2uxnJtzRHzcROk0vSMQxXWg7GOZtltUtqISMenf1t4PsTzH2T
Llok/m40vB4W1zU86lDq1asWsiFIm6c2HGqvV72/WwUXvtODIx3sl7ntrGYoY4DZEfG/ayUFSMDR
Xt+ExjUwXhZ61WkBbnE+5r0e3uUOMgarOpan4fCa4RTPPwDA4jTVZUgsQZiV7HydMQSqdLzeATCY
ZI++mbVahuxpY9CHaw1F44fTqzupIaCxLLReQAb4NWJbAHIMWYD+DQGZGVEW1y/Y4c5uZydKMkOa
H+2GENZ8OQR7ck9tvkMIdm2Dwd6yeH5O4hRLmnnfb3xcc5hk9j7PeErShEOnQelGUEaH2B55VzmC
ad+1KLHpYUu6LxhNDg5LKhZOmZlfvMElMG7FHJtLab/zkJev8JkhIpxTQDC01IjHBSBiXHLLhnb5
aJ8tUnLGn6DLvmcV0R5ziHIrEJppmCwHqrUwSroTScyvFtya6DJ4qU7NBnZC+ySRjpqd70SAyLeL
9IFqDRM7zx/Hqml+B/vlCYuAqSAtrQD43Q1XhSQePd9Ff9ZG36inDg26UoEpPB/3IcQSKy0vyAhX
BuObKaZclNG1SkfzH8OLC6SaziY1TBDyyRvNxKbM82X/k2AKNOF9P1CICRYDQ9ks4506eByZWq6d
a0qGOGKjowb1rZ6qQWNTL5njdJMexwEkNrkYFYAoZoPxGm7jbPS2EwyFVU3Z+X6AK2TSk5AYUBo6
axwJ2x8GZa4xMN8WsgPJprvq/8ViaVPIUCs7Fz/B/PrHtBwDBokxFufBbO2TJ/bY0vDlxi3/Gvuc
a7mrxXQp1xAB91tezm5SQDEwrdYypQeqBh0KSF/xN8AeyUvUKAVOYHTWcOU4iJr4IrkvRMv9Ly6I
fGk6pNj8TqNf8X28qr1Jxl2AogPmOEU0MKbcGqsuTRFqSGJgCvPk2OPlSXRe3sOh0idAue+fz5xS
h+Z338CL+hWGSUueSfqZjhiVqitzH9t2SST+ThkdYlc+f3xykgXgRaV/VvRqQsnw4d5CeUcSeTIi
/Vgq/ylsk2/ZrMWfl8MdFqVkcciy+tChZeiJi5Q6b2SqQ/Nfgr/VTSgKgsWsG9cQ2kh5oYH3MPfw
RROqAgCOHkgF6zDiqe73xKkJrxniGlQSvfP7ld2rJJIYuZ7RssJe4VZxay8JqEtXbfc5ol+IYbgR
UJYXvQ1skReM98ldNmLkW1d1nABV/7/Nb07x9pfdjfewHlNKVVIWUM9ARqg22Hqxo3oQWqn2JlJt
tS0SZ4T+vNtch7gDkedk7vNSRVem30yGIvw+6Oq+VvI3KtmgVjiMkn5iKXcJLg7Vl6Zw04mKIksT
D1ubg96+Nxo/7UcELqNJpv6GMFTnKv6mwwRTBFn02HM6P2S7cEHGlV7fvLTtEXq3QxjCGScARH1B
29HpsJBarfZ1YPJqCv0oVYj3NnSDmM/pkQtnChTEn/pzcvWqCbo0TzBBvGMVFIm66fmMVlA7QeUc
k1hdjhZF2mBfTdz3egRxo3/XtZ7HfUrehU41rhHg/V0TufLtEHZmOzpNxtI18NK4QUqqm2/YMwgS
tGYDM/BWwlNR50FzTV1V6dfx834FxGk6pUcDWbuTspGkCVEW2SaNH+lGbN8Bk7UoVsNyPYPejicW
PdCIkhk2SnMt4ZcBnQ3jqsiT2XzyLIo7J4Os918w9PeTGCVHevK2gCf/dXjiXiG+Qq3iPQjPfQxC
twpTY8DxPsHVPi8CUPcIF7xEYJIJzPXW4hN17TPqEohg4u32BIM52PrASEdWveEK0KvZsh6uIo3a
Z0+3xxsIGrv5f9Z+fkRoH/0ZT/y8SDfly2d8xV/wFlwx9HELwojdQs9vc9YrK9whsyBpISm1TPQC
yPuyEHfBwi3FyNuzZm4Qcv0gP30TZdpLip8JvVzjEOxe+c+gFp+6efAFoLoSKK19bBUFUbWEugtT
ZLCOEN/7M05rqq0WyQrVjJ2Pt2QZxVbnTQYljxkG0lNe1pmRSp0Xt0tWF5pNoiv7aNtFwP9EmDus
sSprtCsKW0Gm5f2NfGe2ZiqnSeOlBpA3g7J1ZJAPJ3W8OIb5ZG0H2k+sBqSo9yPVvSPhiKPZ7axW
NuvBWqKUEiJDEDS91+U/37DdfFX5L+3a7+jPB9qTr4kEAMaaWshAWwU5DIv+AwhE8keR953Bd5+h
Pzgy9tj1kA0aHA70KVUJqrPxiZ7j9PrX98YG9/PG0scFD4+k3p21Isd5/qgIamDjddpQMGSeGTgj
mUbci2x1w1dkdaSLI+GdtvATimvPUtVLeGDKpUypnQwRPjCCL4fSbybvr/P2i/zuRahG2VnkCoTp
mkdIoo7jfhYoqu7cstR1u787sj230ZDKnJlAl+KPxGfyANcJD82clLg5X+nx6NktVGaSNJt+/UKJ
aM4VREqYwcq9pDEIYoFsMn1thaz1DAOUrM/Mb/XHYFswphvmklVAFQ5ooJRLCjc1SRC9UIUPEFWP
OqNrgj0Y5+tNmEUd9yQRrPkYNfYUh+T2bWSbc2YqAhRkZ62KFb6EI6ethlmyvua2Awt74PrvEtdL
N217maIyv/49A/3oDRi57mvoCwhI7n7icaYk9AFGPsum4WB4Z+Tx0lHhs+dIboCr1XBREPpGl1/d
3kk10p20KMxQcuO4FyFM0Jyqvndsm6970FcXGh8Etjhda0nUhJuVlm6oM1yVYDxNwvwG6gAOiCOp
2mT1uKDqAlN5CKtT/5TGJ1aMKBl+zUFFe99OGy0ta8bJOVQhiY+TK80Av27qvGIuImA60cz9uOEi
CyJnqNvd9MnWpk7zvLFUYtZ+DzFaFLoWodnMi7nYuo08n1rQRh6Xvm1f6vRlm40kO3I3o/ct2b0f
TPOp8UTeP1dK8IWYgokV+cub5TjFUGWTLYGe3ldz2n8IrAjY1Z/jWlVqurH+K+x2DIHVw0Z03Jvs
vJ8kFU5JkkLdXSUmAT8EQm6rl9eu4CkjleSWfYGy0UonMEWGrE8YKxxskh20AfnX7kt7XJWm9iK+
+ZJquUC2St7L9lsZ2CyNuqjl0FAKAUmWjC1aJ65Kx0O+ZoTKfxrdgXactJq3TxnHwQXpc1eXm4fX
w/20xCLI+GC+atyt9rMLWFg05wcZnEM+pNB7eodjd8W3h1OTJ2qkurlFsfEICRoghnqKtSL5b543
KjQ5BPBqPvLtL72sG3OaCDLVwL41+m7g3B5ws2BEFmp9liARxSWyrEWJ1JvON0Fc1fryYNlUBg+e
qirjLQ/9MMjiCGVb4/spXwZaLzUfbhO9hPAUy3KF2bDR8LEccFjfkRuTPgq812lhDeD+MFsXKv17
snFDA2qbzLgkrMeFTdEjKD5gICgJW9NUT/t7u2AkcwEzTAJnSRFPAHChnSf79IbJawcZtw6IqHzW
EyfuCSX+l9NolnROEf5irkvedffLFlvzCrirkF+fkoxiaZSaCVf1d2JtW+K6yTzCaCJlFBSvqPzw
kGGuFCNL/jZUU6TPj0MQqrTt4vkrX1GZfEniu7D0ctimKUu+sxRkXx2fOT19ZmnqIyLj3yBpd3VK
2V0flAp/IcoUNVjw3ngq5L1cvmZN5xWNEbJTUJSnijzgc7GFPEd0O4udBihtHwlkoMlxDz4aVeSY
CoG5LhXWgTqFxPgdafbKnsT03RwlExVMiqtVGGT3+TWCllkOBVM/GT2tt14m11O4Gopx5grzxAm+
dMpH8CqRF9WB6qB1dDtLD2GZnZSS0f9e9wVgswcoDUF9RoCVPjFLeSmR4z+ccm8oumdMLcFjNWSW
Q2ALNfyeIBs+4O3tz9FMJ1vKQWTbTbOgSP5KLmH+fhWX5zlx/TGKM5wxjRbdtuz+oDq5eip3Z3pW
oLEOqw8PCmjA46yXWY249vLUnltUgM+Kq5l13eCdA/5K88DHQZqBOs1L6CxfDDNcPc6F1K94KETJ
09HEyuF8fVUVVYhqAVYpEtcrd49ztf90asBjlMCzbnDnYNN/Dq7NPplMj6oIn4DrKEbxswP0lq9k
9ZDdX7iTpwrAX9psoNLlFpBNXSQolGm4UBdEa8KACdQkAC8L/NZCbGLnDwyj3CbJ2lg3Tmo04y1f
wNlZ3EuRL7XoYpAiKW02d8gnTIFRonWxE3oRJfXtKaujEJtfgvsmpOZSlFy+EjNT/Fcb7j/gODIk
hDg+GSS9BbLFX2DEViBBvSKhrIM9+8vlzd5RC57iZyFgashKGSOCP+fqKSKEQi3FZtvBvAWbkSCF
OuGsNlayGLeCh1HYe3CQeuV4MUQehNx5NAk3r7kSdrqA0t1yRwk3hDdwcYuSNMHWMLcQBW6Wz8+Q
kjMFrEa6OENcAmSrAo3wxsWqxLL9yEovCjGrsJ8qodfUiIuN2FHzct5b31JUY9WbluICjKCmChpW
dAn5+cHyqZzpWFjHId8gqq35Nu5kttKpyS4aMIyw3GweK5uKCsBHL1sCKPrQ/u7Q2zC0OmWU8d+e
/lQ8jZ2K4clajm/7LbxpdbNJZrVeMdNu1xayE8DmELL9fziTzY7iJqvl8+K03LzoviIyXY8xICXM
9EVbRlXp3+C2cSWP2t39vPxfJJoSlXrPOLV9JztAWMJQgBtELxHV201/uetMC6/d/hIQ/5BR3enU
69Srrh972By/WhRgwsX/g5mHASv6uJcc9DwuB44P0pKzHTIufXJIqcLVc4KHh4Rl56wRiUI9ytsV
pzNvliKcuOSKuAvLC9XzaIaBWB6EtvMgbpj+v1O7kGDQIWayGkF6DFZmnJblBC1XEfkXZgdatB5K
jvM0oUuSfIWd32EqIOVsEAlKgGtitD3HwLEuqbxk6ms/hF5EsRPs76azw62cvYYyTJueZj+TZGZH
2LWeDsRs3mxH+CpqqBWlr5EH0DAY/zbmDAXMWYsAPd5FkTanCD6nLIOziixXGvP6sk5OlZ4T+GZH
Td6k+ZxGVDkzOwQMehGnNIoZvg5iyf4DSxPRjxXV/dwwWQz7wMUuu3R2l3i4xMff8ASjsLffIRJH
nHfFEgnWdwPZydMbXb7M/7e+LG4t2abzaduTYqwdKo4KY1Jd5wraHeezYEPBS08lVQ39q5n3qz+k
Vk6ntXJN1WlznF9yfs/507y2fZCxjNGouKyWtxVraFY7/6eiVUqtrZN6d03iTnfUGJhbWOKgN1zO
AdVPJWvh55xCFVtCXbjxhXAYj+GXIVufKA6CJ0cvFwDznACbCUnA97xSjZaP4lO8kuNBJOux0w9w
9ScF8aVZMhrZsV2XpUaw3c61RCHbJpOu3yeNPV4/fgYg2iEpvl4HgI2vFCM1xX1eVgGuSgBK8KP3
obQ9QuyguJic27i2orJ9VDyz9CkEWv/CcpS9B7KWAw13Krn+KRIzBUON8e7UZirbrJIWBUptDv3D
Ek4ikqq2pP26oSZm6PjsR4atWcXMxQZafasL1BKXnHJlPaxOaT+9yPKZp2/x8WH/BAHq8RgXxfcN
le6ugo6VvdW5hJt63sYzU6/QA7RuEQn+6lFKbz6mUwWzceHzDHOgzgeVDIZbCog4DAUfh9iG1Mbp
8ziaomF67ajizF+40xw8Ag/GrF+LSAmduWlEch02LYBK7scuKMZfvA1MUR4Kyw8EJMGCeq5cezds
NYDczq1ktly66Z2JlbClZMPGMEgl/kKLnAM7fZpZgDkl6A/vfdt5h1+7EE87w8GqDZZYa2PWrkGe
R15Vd2Q5ZfU1UN82lysqg6UCdzKK2tlx0Ya0kJ16kD0opZLqL0NGaE2a0JSJ+ngR5LFc5zlsWGAP
VDZEKFSSEhqJNqg6SQnx4IqfHKl3xaJBHinM1sWuPPydD1mok5NEPiQkzfV4xqlsUTCNwxHPvn2v
+LbUa9uuZC8grU8zwh6kCWSGI6yue8HDm8w1lMDzoJQFb0mNtKzte53DVDjZytIn67ekz+pH0NAQ
j4l/UyRmXySQ+ORVnZu1T4X+SRSRvSRB6rBtWS7yRahK77/nWqZ5oSl8sgCZBHw2MGlMaxqpIBoV
+sYp4zN9ykrs5K5Wbx3KeZd3ykthwaqNScFrVcBMqJ9n+WA4JYyXJskBY4bO1+rzq+ejz2YR5tnU
ij1O3Lypqq1XTL7Lokr+yhghesUWBIuh2WJphJAODR7T6yapKfMnawe5RlagscZlxotYtSC5KrWX
nGHESm9RbvVwpUFyM/U98l/zZx3+qivYb267xohk0u/OzHGpkheUIUKs8X85pcN2ThcVO7P1Y8Lm
slitz555D73gQOxDhPG0xSw83OzqA2E/qcaMTRakeYeqjkJc79yD3qB6Ek2GlBmTMF4Qh4bfkRif
gtSiQ2wK0i61NzJdNpEkQF3IR2h9fswQuknLj8BEO0vSk56/hnycHGH9MgfnyRU8ekAWIRIyOzkU
S1MFHk2tu83skmw5CyLN+4xgM8pOy+BY4UOz+fgcxmEilLrhxnVLBO+KsPdZJb/SAMU91FhhBNwC
ZQ+i8uXDm6qjT2MNp5A4yro5ckQLdd3i5zHMHBQbSx9t2gUqoWWzQnPDUIJPrTghyOFnNbqfTRCY
hsHVQjVIHS523GXIZj36wTfhJ3xTIB901Iotk+wr3zZaRU86BRAslHYHNSFkbIXXImxJzmIYH4Eg
1/2CVzy+C6esqq7zxnTGstUure2cPBIYNYWd0cFEnt/pMfCQ30OHVa+XrAADXOIvI3nHCYn7LwcD
mNXIl4cwAqqHHs/nA4PJXU3H7CuILiCgJwPp73BL6D6ggOHpfpHgGTqEN6n0zMHk9I6rrFcIEWJf
A49I6iLwmJzt7qLkZ05nOrITWkAd120zNSqQOnwADYjY7Nk1BeSesVDpUVT3KzaMK3OQi7sKLwT5
sM8Ck70KTlfrW8yOIlYU8b3eP+N8VbhkxefFiTc4cqQyeCE+2k9dyUBmIHq8ck98K5+7l/SKmpAf
OWsSnQ+B+HkVB4n1I3XQ4OaBT1NpZajXPxehc5jZYDSRDKFuFlNwtzsM6cHzRnXDs8IKfb/+Ag2s
8eWC8BK6bszTXyBsgVMXsOaw+jM37EhD103Ue8n4ObAz4mybWxeF3bzxnVDmN7kecqbbI/p2Iki6
uYONfeq9A+mTABRIg8gj69bhB2lp9+Ic0QyE+VXqzZtSu5g9/dmjKKVdrkjBQ06quKgHv00aEnAD
QxKUyyno47IdHdg+sGbQHeotg15u0KwOGG/PIm9Fz9RpiwmBBLQMziZ2l6Z4dHf2PUD2uOYKqrcW
701OZOOffWC8q1wsB4jGfb7ff6IlqlEkjAnBTiHD902/UpsOCheyRfWU6KpdBSVyXwzwEB3IiFaI
efoK/g1nPPsoNLjptgNVZkVotpKcC9Z1jLfggaNZW12G8Ve2AG5BmxdgedtkvBqsWhhufas/BGkz
kvpK84fDPoUz38ajwwtRpfeJLxMVaGLyGYsuGc9S4McSQi1AZwSaobGXLP1VnZOyqO5httZ0oJ49
last3QWrSUC7xAD5oucuMnLtmf2YwlK+Xfth1Od/DURvLl/BR6lLVpN5s6fhcSy/4CjMIW4TQD+t
03HxvbHBBOOtigv7a7zhhyPRE9FPleXlcFouDN6a0RtSiLhipWHFR2Dnbdeb+mJ1FCZypE6039Ev
OoSM4/BONcZlevPZFjhiX7+d/0KTqTLN55ILoVECHg1uHZWZaKZzLKMzaV1zw3jHwqrMeqD7o7f7
L1XSo/btSztUx/FSgBU8F/Y2xwVz8Qgq5rqgNRYwgk4j1Qdi+cMf0Yb0jrh3xfVOJnP1rokbIgKG
bLSTDH4iD+0MWST5oX1aW6yH5/bUVytlniHeIZYX6YujSdqOWYuMNR4H24TPPE5jzSeCtAxBiTMG
0+EYdgoDee5W2bpo5e8Dmh13SPgC5bJ11xuSagPiSqEJgjmu9up3y0Ab4eOVprJjKelRUMA7EZ8a
li5yb7uYompaLne7ABOgQymkOFLdxasGLadzBe0m8ScA4O5kLA3tJFB+PkwJVTwUkFnouDLkCkc5
tKdtmKKWlByCfwVqS+ZbIq9oyG76elgeznmUuS/wbvWdBr91WAjPpTOFoY/A5Ao8ClB0NhqPc1pi
viTxDLaXqzWKzOzEvse16hsmZh9vq/Px4K2CDI1vx+b/vfTDm0+HstvcIlLvmEeDHuP2lid3SLXv
zA2oPlPT4Af1jApSlNRyanZVSDJamuZAelEwjDUvIxRgYQ0/OOtVgmdQhjyawCqHgn7FWGUMWFlY
U/RFpnSSl0tSvVvptdEN4Wfqkd4xtUDAzWpvAbnmoZ59pRFctQaY/Rfs20D/AVuC/1fjM5313L0O
oy2xuexJBzmsr9z2poaxZBNENKJBUV8whifcrGX5R1PKOy0ERzKQArID1k+D8+stoI81hp0/QZ3m
3R/2Oid+nnpTIUBXjpJY9tUhqPhnoR047TvY/1U5doFYqCFXKbtW5QMAAKDhU7cho8crDst3db/n
5HRewJnN0SB7VpJ2+cachJO+f5qoPvhYnaUOL9L19PBPIX6x3CYZe28/CoPmUXpd0vZ7hF3GOWhk
vpVMpm4oShRHuET11Yrl5KMfZ+GRhE8NYicrAcJ4hh7x2r9HuwvEcUYdI2xfgeK12jNIJLowbHVq
21n2LAB81HAtLufJSU3WfRl0zYrjVw6krlRHOIM/hjV3y5UjDNCgUTgY/GCJmPG7W4KHDlY1rqrp
p/K0mzrVYFcw2TCw3m9uFuFtiW0PRKhhtUGHsC7eb6SJkqXIjgi6oBHXSSLsZ798/TmsXF4hY3X7
TUi0HBDswLn6BniqPy193/e1pxC88juXM6rAVnHS4e73Hoo3unaYrVrBF3rnfY+yI0QS8/CSmrG/
biC7yL6zG3aG6QR0aDVPOLUv3ISB12+A5YWQbeivuQcOn6CX5st7BPLTGjH/4qebN94Sl+m7/xrd
8yO891sPYL4SHhFUsuFJSn4Cm5Y3z9MRmTFFsTmyVJhb/XIDDyYEUhlcOWhc+FlwQCH+DldxKjcG
q8AnhnEV4e4jDuT88V2RFxUykkc3raup0GXkdCInQaD3BsysXQ3Kx6bRQknyJ5MOh9FaSwV1kVzH
0haVgpn174Vjc9G1PDG8oChLC/otmiwccW++rf6yXg/Bdhxuku9j0cmxHj4CZOLBF9TJDBYGROG/
Ko2iFkWJqYUPfcnJgQYhoLs2PhFER8bbyu/AvagOqi4FxrXRBtH9KgVbkpPRGMiSCSRGgj2fY2fU
SLOjYijVba2WLg2vTm3dv9j9Zftn70xLM03lVcXJqVXLbaaw32d5QKkcdf1Pny4G7DDXQj0GpenG
kKWi//JBgqUs0Qnm2094qtBEk4+IJwy4ojy7Gx8Nuuxig5m8RaTXSRjf8LeqdpPXYdTFFaH7u8yq
7Jgw4rHbI9eOueMNFBJZ9sq8i2gI65Kq4YV3TJXtzjlX2krj8VkIHJH2Ylzzrp64PdG42vP9vrOH
mRE0bA0UiHysLEe/i/RTOkYFKg+3vc6/eRg0NftvLuYWkVkWHZma0qSelpyvzdgJjDe1Uv14b5SU
vYouIpX5yFHNVjyZhf4g1WV9VcEIep/zMPlOdPY+l2EDJpUIC/N/y213o1//b4d0XdZPXQnk8/Gm
o7cTvJEQBtz/09rzFdvigkJtYRumr9+o8WW5DnyyTYTngPjJFZLMLEcIoe3BokiNC/Lib8bKbhrV
u0y37sTS2iqMoyRIC9eogRELEDRQvi9sQpprXqibqNxj1q0Jo6HnYVbuIej/ppZOchPHw6FS8qTm
5z4013jnZZw/hbnZcWhTFyZnNyYz4pL31LTjU5C6uinUYK6BuvIJNzFQ03ncQT8Bj5k71h/SePMx
bQAVkaXRs/qctSQ40mP8B6EuMQTeyToURB8aCJq1vNjEbnngmeXxagBzwJwdI7COJ/729EAKCa3i
bIECL9vhKUQmXTyExsPfDZhIKC+C266kW6b8geKsRDph4w5WLonXzOBxEVaZESg3kMyR8G4DKQm0
baVSeuxJhhcGjNqaqosayRjzalPc3GxBlbb1NQQU5WNqPQI+odPCw24O9q7oYqlnVct2+G1nQLIs
PC12hH0okwsq0X3BRoQwkpUX9+xjDQuH5vxLPxVo1BxZcUdkIp+Op8g8FpjjkEUVy/XqvbZ21o8f
fSkpHTFkmi7DdckkTitla/WeI0j76QYk6arqK1KcVaw3Ut+X63ftXpi+dK/+WoV0/ZcaWAVtLWJr
Ay60l7XsmLtC4zrber3QE5lyAARfZCUJq8nCipsN3u9bB7z5ZoBiUEXpH+gGisOqktFXPkr+uRFa
2xT5wIlIGEVnUg3j4070oCu8BfNwXAc7Zg3BMy9bQI8LIiORUGGIL3ZzAvEbD0KgwMdbKjI/Nr6f
VqjCY6qMzJtfThMI30SMvFqM4XngRqoEkTGpUFg5t+Dnt7CV2Mj6YAnIG1tWcs2DCVLBPs31fDaG
zgXqWspFLf8sJe/p3/XleNXBuDOyvMWAv/J1sRz/Ekrs6hRmsZiQI2r5/qh0/Ntx5jCLxqsyoLVR
3qQeUqIUrVOTU6k70RrLTdEZxgJos/dZXn1m4tSNp0uK1L0gcxtUC5ab6+lNJkA+QlsiIu0sALBw
jgP5uDs7bETxEgWbxImAEPuVVf4wdsaqWDGdQXu0DkPPBG+vO+mqfmQXHfapLpy37A/vqMCYlX8X
wNCiyPuy+pssNejbZufHwdaA7wGM0eCI9Lg0x9dR5979UFISArwLGaRkXhj+PE3JIW7hsw0KfRY8
w5VSWiSP3SLh4d4FTtIDK1NRpPdxD++qpXHDw7SyP9M6qXDHvwoRmPI/jDp0oOGxcPvEqcvIfA6U
16hZqQn3+ltTcvk9xPF+wb6KsPykjsQGjFhK0XnpXupNtsTdHhSO3BaWYKYmCgYXqKAHA3ntsnbF
Fqd9QGEi3ZLtBk8FFzMu+awyA0bOXz9G2k5500AWUKjXcZjWJqAtOrSZ0e2O4a0GdiELZZuCj64e
OMXDACPiPqf3aWzGYoIIN6QH0tyhDuBQP2M1yQMtuX9oVO6cQSTijn7QsJQfSJczYghd03MttzCX
Yj3Lgjtp7oUqcq2W8tKuCPAEsVX4MP/kyOr9ekhMZaA+xVGudLHYQSYLzyhFhmS2pKqVh3L4HnKN
ZSadbtEHwWV+KQ9al0OEdR6+cUOYzr9BP7THfoMHkKgLyBfZgOTk5EHNKP1tsSWWrb40AFgR0MNp
nO3i49iZ18DTUYtmAz26nJi+iCgWTZFwrI/mRZfNI8AlyxMNnBlotbnJEGovCox5VRlVP5OHK3Ig
eKq0agdyadveyXjbZKmLyxSm+ptqmM0JL7oiCLj+Cxori8Yhh12JtRy2mQYgorH0ISRWEldmivvv
oP30S2m3yEScmyuj9UbVuZjd+t8bxidInxx0TE7dTd1qN8trDeNo+Y7GbSyGqYoJNwFykbKmn0r0
Lpikbz5AA7VThnAf290ch2AzfZMKjH2i4po6ZE+TcTvT5FzZGP+MOlfDGhC/yf8/akcpUPapujd5
+lBqV8yeQlfU2seIe/d8rptldvspGqo1zCJllRpjExCfAlhbBuIxr2+FwrDIG9tl/BxJL4qNPbFN
nvtgtV/EBulXHmSor+F8wqI5vd3UGNTOt2oKEuxGs7gbnRjwM9k4obujAhp2wvynQ6OcLSlUWJUP
5T+ojRrgFLi9kv2NQDgF+YdE3+jCH63jm38wtpf/sDqDOHfTQLJq29hIY+eZVK+UsSmbWTlnUFqh
ufLOsyarUehsnWYbPVuPpGxqtzugSBL09EbCiEFM9MB1LOELEcCl+x/bftf4jmEGe+MvVdUXdq7j
qJIk05+rlXmkDh5sJjH19sVcr4hmwVmAXTbk1y37IB4IkahIjDOuWlpPzVjvpXkHwqset80ldJV7
8KVqMM8KbW9u1ry2W8IrgJjATHzVR5Ll1/AO5YPuoit+zfMjDtGehDE9zPZdalvAFTfkvNnJNUxU
NpdLvdFb49lOJ79P49jPhL21fq2GJzEJG07Duv/XJOnKHOeEMtVzcHnc8RVwUJzk1+lh6H5yJUol
zYW8FkTATuliKVS7V9+z0g53Jcx2qU+LZh2etG/1UBOeZX510YZ7k++QNiN0PfZJf3nwVvB1rUt4
FD85xOXHCYmGvsLUY8fpMIy/snDJvODW+Ie+yIY3Qkz7c0ooRaXIu1zdegC6NYxI9PJtQwdAScwE
d0SCwIDKEpssZmVp3HLCOIf+UeXofbdpA3rUAwvcMPlh8WVAvaRnEs2717U+hgjuiijQoUZtJqB4
6PfUJ8NLgT4TVavO6AYGIiCwFa/8CwPk8tM4fnNkYFRPYIONOHancjiU6eNC7MxyDbk41wwxDurH
E/UQ3FKC+5OjwDi8UX9AoW7Y/xLVyf9DWfwBtDchknM6P07ptsWEOFccxMh//K4X7fHQ8aKyyTSh
dhO3AkGhWKVvuR8qnq2YMHR1C4IG5T4EDuyNXULf37rm5mcwIhz7cqBdTwrlJ2rrYkwuFaibm7fD
lwDJtThRt0gjulNX4kIm0ISGLmVEOq45MLRwyZIYB3txnk1K8HE8M8Z2LU99dirO0w29NF7+AqfN
Edn4wpXvIlPD+s77qYhX7Ex/jxZDgvIQ6HCXrqWJf97DzObDrsU6WGPyFux2WiE9pr+l1AC4nN3V
RI4GlvMzXupbOiBZ0ePbIjTUyXgYokULoFTO9O76rImaKMtwfF6zgi+wyqgsl9tXW6JBk8f2b0i3
kOIHUrBzq+f98UwdioaLZRgWzowm8o4GwyFezqiIZcoPHOCzQsklCQeNBBNlcbbpA7bM97z67VkF
sXA/t6RvaKaG7LcBZOHmUdh0ni8sX9VFiGgQitWeuuUUc9AAVO+RSJAHox1grWIpBcu1c/W3WKnj
HY4ebNQpBnl+L/GsLXRMz1bY2upkVX4xV1GX9BzyIdri90WF1rtcTWu09Kyp44Sy3vJKp6GYxPIU
U26GLrUH04ccNNqpmF8dgKd7P0EjomsDtjAez0bQ+LNtfOGDwURWfbtD4ZEgV0JykPL1S9aOVXKk
5JioNbey6OEJL9V9QBc0XdOmNQQuzgZ+jzLVfF8nD6OlthFpn1wtcrZfWC8UH1k1nC7Ezp+3iFPy
j9+qE4++CEcqbW95X8XI18aL5QmBnyWrqUepWUgpZxoDjil3ZmzPgniyihHOEw1Po0Kw+pv7Qu1g
VuhSoiDcA8gElS/cM651l0tiYZoLKA7BJwYVEXL36oOdxfh7nRLpll0WE49OJuh9vCiUcfAt5e1t
96q/kIzonfpxQNOOsix5CDFrCXpyJmwaILyP4JKl6yIiJtYqF3L3rP8SmQ6/Cu5nZRW9xRP7kK5V
G+9YVdM8RBTKub8XgHQ+qHPYbUORZOq3Ks5Iu+5WWyfDO4qta9cGGh3IS2JZd2eMJELyW3Jx2YGu
KG+HTOH6zh6LDS+/p1pvFddFE5C0uhCTsLasAbjSE6B0kNVVj/OmS0EgN7lsR2pOKTv25RsPQoCN
M/qV8mIiumSWMo7DYkqHvJeh5zOD6nrZv5YqRdJnEZ1eZjGCPuLlB41RPEmHfY9VzVkQMbKhy+hU
7TXAqdBloJr70fqtwvwC3hd68r+Zi0TSAOybPcdEwVdKUyMci0M1Ct0ouAhnPz4TiHXqm2COxVfJ
NU0XVAZEFPNDiS9Kr0bB927/UlB4Z5xM9eaiyxBX/GR/GceOGExvtgeBnsmb/W45WH1rri58ro42
PJa2MXXUi/b9PAOHYYMN2QYpXlpdDhr065G7x7xa0diegPIbQSmtekdzEEeQynlj1tLv+jdVJMEt
eWI3AnBYIEoLrk6zXieDLrZprkxlTZhPCgGFvlaT656I/BRWASjUnUBKzlSx3rzK/fhJgJXMg/kX
qL8SZX/C07r56uHt48E9mK4q3vU5wtkxFMcPxhqwMgHpvBTruG9R06yKQHAEaVS15jiLmdq705YW
YiByBOYLrXvqSx/9af8hvEMWEG48f63RKVjQK1PsyuBDtrTkrJYKyIQpH2zqQqroQCqEBZR7SeY1
FjbJR6y4RCp9OIgvubtqVxVZDhA72xiMEBnbPmP2MOLQ9po1zuyg1fZfEgmYGGoWUL2fc9+OoDFy
6cZNZXpFD4JAy3MG0lEIy/qerGNNYDvgEoO1No7XlX0nH8enUcEtJ9qS7Pt9kR2thete7Ogok/Xu
lkL1ExssMg6tYPl2pk61eXfT+XN859oWluA+SVc3h/Kn+jXwsFLx0bGnv7cBHMocozMp/0EPWM0s
hHlD+db3h0KQfexzQmDSmtdlCmnIGgLKuseQvrfcYugHsJk7olefNBqY7lcNhF3ycCM3Kmv0p7UY
GvXpYczuKjJKHO1yUOoWySF2qY3TtLNDLrwXaT1spXONe30FUX6wjjpLSmotqXscb5tQ1nIlWeeJ
hKVoCK31NZZpfej4tY4atJydObJlcw2sqNVisuv+bqXjYJtu6cv9SQ8B3/YWWRj1ThRjEcySsdhW
E15oxQlpjsBRrPRydxXvG2lbzmx88WY++Uxh8+GRjyKaQ2hzOQhEdv7gTmWU+i+6K6Y+oziK1bOU
T0DtYHyupFcra3pPfMfJUo/SCm3MSfjVyl/ZCUWrExPkIlPoetG/1LECwBnDkS8W17UWboU4TFHs
eEWTcoCbDKEcZc4wuK9CRKHIDZqLX41/TvoXRfTwO6vOL8GUefOG3GpiOnLXj0kdPvkYcwqLYcAc
RYiro9zOxMNHtWUK/G1gC0tbAPKOKZ3pwBp2JnLW66rQw2fYf5noNgIJO5+vhBaihulGWYGk/Onj
9nFx4DiqLWyX8vXEupkz7oJJTrYOiquNJBpiAaI8FmuMelxZ0XZBPznkG9sU3Jk1Ttd1RDgbtjal
PGGutR6el+seRG9Fhi8LdOvYy8P1bJaR9trNIo9sagJILj09LGx9owaaBGXSAEszCWOo9P76Oi13
5X+rVJ7IpK21iBv85TRevtELm21kIIZJnfUj6w/WmeHlero8Z3MbD4og2HHL4G/Sxp3+830+8Yuu
jeqJxh+S4yMbCZ/0dKItJkdjyViIk3CiyeSKfFUSjs2xYx/kX2YnTcl/IhbHrTPOfmC1MTdZxrck
jxQ+oejPWuMX+JoH8OtnBZGQc7P08RhIOG5pj51krO/neVfQzj04QIBWktd2y1LH2lLumqM2kBui
mGe6xzjRpVHbWOoYkxhdyLGy/MnLeE6vdnkdKwoocca0YOHR+yCGFHAwXnPU/AUxUtD6F0ZbHhHi
BEKMgynMg82OXt/Ux47gqX9gUZd7sGy0Qg2j+6WD3ZdsJVuHL74k7c/XNw5dxcuJl/FutXkb+Yy5
rT6NupRXOS4pA+Kzx9DEak11Ti4VPBmo4feYH3F5KZlJ9OVoM6tTdMDEkDLsdf6y6MwIvAuTCfyn
5uoqLk19YdUrRDDKHYgCTo8ujXktM6vTmX74DamiVW+JO98z+iYFJ6aJWQigywD+V5ZYquCu1aw3
jhzuPbd8C/Sfcsecmt+8/AMw0Gx80XMo1PkXwYSqe5GMs9nRG/XGCKnIdfo5h++bQJt3OBivAg4w
DEUpJu80sbDvIEv/1wbsatIzs44+hrimRVMlsHGNOjrcVurxFMMhuOlZ+ARkoiROf3ND/cxDg/f8
BRc4sz2LH9asZLTXVciGKPnej2Dcl40HtwfSTKVrWWKYQHuQBY/zQ3mG0Y0+fZqPyhPEKR3Zbap6
aQbHFKAvFjHXtrKWXx1al58t4SQOHA9Kc/tlHRnGT4EqE8rr872Gw0ZObrMpFs7po2e0hp52c7p2
F45d/mKA2v221PjmmIcl6TMQPBmVivBfjFzz7jLh1sMFOBsNqg8C/EGkJ1uNRjw4QSDV5JPEW1vV
4xh+z122CVf/dpWJqkbezlvRY69RbWiJ+OxSS0y/zo/5uHdfx9p+ofwUewO3nUD69Vuc/qNsvO70
pAd2gT8vPHV05SZ1oUcwIotcGCW8nfeKGer/Cjr5Ad86UFKeY3BYBYsIV8jq/cC2YFNBGFZE2MK1
syEXUhMX1Scf6vvGEmbuhMMRz8CgdsTSqFuLFgR5PkknZ2bN1UirFZHxRseJFU6GOtLuQqKN40uB
WqWWJMPjiHz3nI9J2ED/c97c31GjWJNl9x8Vhox/nX/921IWFQqAXyulRwwuARCdJGaX6QeADSUO
adRr8N8wKvczKBPyk8AjdmHFBDMYnC3NjibknWF85zg7aFyhzbZ8X6KGq3Qe7bshY5zOpD3Avh6d
WfuhIVEmdJ32aBx+rMPlKL2usqLODVN7u9btMuwqJVtHKnBp/QKx6KTYB/bepgWRHjJcEcLA8YpH
xqEzhbgeyh37mSKUu+keDQXVG1mjAmeGC6GO2Djo52HYUp7MM7wmEFqXfe33+v28dD5DkNcEIZTA
KZHnEolcX54T3zEBmuNBmPN3Rap/kH84dEtwKn4vW1gWDyOiHSuCqbnbrfN2vO/1AgKQCcAu2vmQ
SS3+bVkXbNxUjdTl/+i/uKvTyQna6qBEExsPzSFaxCK6SWKttmaIwxjZW1YJWn/Jrn+n458t+hUb
63CJNnxY86rNklXJyhKeMA0MOisf4oDBcHpRMRHS+/sRJwI0V0UVBpBx0MIj4QmgHa7kb4NX/PZC
N0XqXwF93DcFpPRW/Ds2V98HnPH4znsQdgMQFg6dKS9RagRyCNew4dfubwGOvxduxpmw2oUrpD00
FO8aUELFT/Smyzs30LY2mqwm4CFhFqSL5qgiZmTip9PQ9WPW4/LuMORnL6WQpskWoRPeTmW7F1wy
imvrbNtERXUzPAwJ68r5AuGCKD3WLOC16FouUUYdcCelHPj1ipiGoa80ZdtFex75bUXMAJxo++gd
iDAv9OZY6HIAUCa1GaCLz43yzl12KZYkRP0KLRWtoC7INpYTLhxGyUITsWPgp9I85NnZ1CnLs018
+DU5d3Gt7OkReLap4Sa84i9SpJmLDZbI4/ft20B+MIk1FRaYvGgSaEpFhVnGTyB4mf9EOyyKSi9k
9kg1eideoWQI0zHTzSrdIIPyNHRQbq86iask7hlHgGLUM0b8X5ZYm23CL7ncbItTytc4e+0VaqjZ
J47RrSqXnoF837/QO8SCDT2zCLJ6K/rs2RHgbjeU3L8qj1EiAxEA/y4vTtrmX1ZnQD+WMOYDFExo
OLGt6twsKFLEBLz//dFR7BL1t1j1FTDl3fWlgPBx0MKIkzD2hfy8nNZcaDdEEChZQCJJxlA34+0O
PI+ODH0mnItQRYvZDgQhVLnKMJaCc4eR5WEcJSAC6cZB8848hqTYH3/gex0W4uFmzaCJDyGE+GRf
mc6agQAUZBH8zl2iqM4V0sK2XrVSGTkasQN3zZGnNES3C09jCQTSWPguDg9M5LSbiysjL0SPqcmm
QSy9NakwxgQKJRWjfLvjS3NadLa4rIxzYO52nX2sU2Gnx33ULRgj/h6+ldKc0oWTKiVQmlunogHT
FScN6cD9FQitbOcBlgx5Fk9BXjhSuOcEqbSPzkY8NDAsRxThm8FbStiECdPjM5Jdj7BeB6iUjhZe
McoJXsJsNvxF3UTJOnxBkPE1dZWqX3Pdm7htlkPlcAa74FgUTg95Zy6ABoReVVYuprfKAKv+6iea
0mWRFKEhgJipcqCaq+X/YOLNRXGWqtRnyOZFSL0BV3DDOY3eFSgofWfLbdYTMI1f7r5DQUcWRhIV
fJWE2RkRjochoNp5iiUDSHpUhLaoeG1IIjuHMTK9jR6wlfP4kR/li9UuXUNPQWvNeSQe+bryZ7Yd
P4GjGQ96Z1T3MUJButI9iOilwy3EPYRT8frDJ9a/fnKBVnEAYIZyGE0RTI+Zs8ba6yNR5l6Jyd1V
iOO7FZQH1/Vsb8YMi47iXdF9CLm+ubKsgd1l4rVhL/f/qnOtPlN0AmzvrBmhfJ3BMdPJLX/FTsNB
shdNcuf+4YtbI86SsBlExEI5CC2AT4YXHioajc3KtJrcfGQkEe9X2EJi47XykrFhqBchzYj/l+mA
wEk0qVG48ZmBh7vLO3jwPEUlYPYAegacOtJnUMypfdK++EqcmeIZPkbSm0ClFo5SRiJoGqAaKIbt
5WK6eDefIWPe96hCERZiRV0upmGaFg/JbIIjlKN8HPbA+b0yIRTHti9nvku0ntlt1NCqK0QwJyVG
8odCHNui3ibpd4f4osjQM+Hopcsp9LhLY/55QZ0H7TvG6KcJAYPynkEHV+7+Kd37oQpRivEmDcrm
xcL9OFHZAX9CNe2KbE9r02XWmueK0zQhHacdai0w3t/xNG5eEt6rVuZ4fWMYdwHzDEbW4Sk9xNqJ
dBFwSgIiqbG5IAG22cKh/JERP0M5e65TgIk5dgnuuk+HK2s8GLbIAY46kdjZWkP+/B4iRo6ZmRXH
58rgoS/27P2EVfVHTBBCqz1p3BCD3RZx7W1pE9tHgBfwc2RZnd62PHIMUFPlJv5EloAkg4YhbpEj
W0m8UwBYbZ55m8TUJxJ81AlDHpCJXzz4SY1Y+u4LTelB0+j49EXLjCM7geDVsxX4MR+q9jmwANCH
Hk31ORT97QpLeCXhKtote5U3N26wA6voNf2nVK25st//f3YHd+hbD4NVzWTfe1YI6NKqvVZ3aVLl
NORdst0stFjzJdcbCR7WslmYvF0QyfAM8n4GhXdA6UQHD3zob4e7bll4lcOmFlAoiWSWsSfKJ1Nk
Epi9BQIbt+8oTTtSfSZJ/CMgDMBz5vUAJCeTZexBlCSKWgBCr4BP3mKUP1oaw4iDakL3Ref7oyGn
nhxWi3Wp0s3d4IxLSafzWX5YimTS1Pt+5nTauCqKT2Ygk2wpJY34BsVpB3XXLJ13M2ZC+EfxELGG
PHtxnY+3HXRssihdXdNzZDG5pbNVnz9JVaTFUhb+P9wDM+glaavridkxBaej+bHSwhP0Z9D9cdXA
EXHKayssWurcJGugmcnQ1mLpDKYFN3AgjPObyzs/LPFJ6xJugtMaH09WuBfS7foOrW4QvjrN/Q/Y
zS04tJYB48TJa4pFtqZFiqbNT+y8MuxPFUjdykv/oky96SoVPZKBj64CMOsOSZV7gmH406VIvuPi
BfEo7lJYBTseQABLRlL4XzZ1NgxwaK1PziWPzkIL13wPbjFwHxUMpP37pCqrDN5z0GemrAAUaMwp
PGy1eLBbZyPDcHWpqZMgPgW6HW7tClzYfD+zKofST3M0TcAt0qI7VZzJxTtWdJEJtfdHXXzQBKfL
anSWUdfSc6HB+/v5YBX/LyQiSupHZproKuepeQ6Q5EHqlIhuOesXvkIPl0CIGy3IQICohBQLboHp
0JK0XhhbkPdxa2oYiSB6smvmWYtpdijd7HwiHT1r+T7ts8Y+jbbNy+oHu+3NKixA9b5qxbE7+M6h
/RQd197Ad7vo+/eK2zYae3hY4tKwHO6x4HN6t9G7xXFFgNV8GyxYPa3P24qtGEtqWTm4+iPvuOvT
Svcv7y2DjMUWHhVDQd2gCc81/T1hjrgRKrEQQjdNkjh33k7I9UsbvdHQpRbqkBDCAaGYj/jp13FS
rOnqqmVT9Qn6PLemJbwqhnS3YaC7FBnw033MjAz8FVhb2LgUhuyVK6ioUGl/20u68zkoSllQWUfo
hqWMWsSU4ykBhQGoO9214ApGzAYou1FyLGXQkS4sDNvgRECcFCMbOH8E0K/o4nFq3MkH8iXJrgmU
mtnVznDZVQXf58zL97Pau2k8gVFV4EMhsqS6rGm3RijBV7uwJlYd3O+sVDIBV6DphzhIvOCuQPEJ
vXLokrH4WguLBis86Z4i2piTJ4VMbGzWP93a0MJ6k6c1qW2TnUFaxt3hGFC/8jetbBwdNKSR1qtz
PhtDHmtrYO+HEd6WwPefbaNrjljf/xq9DSgiuEN425nIcI3MH/jOKF5X++EJ8hGTNriyId43IK8b
Ol45umnm8jQgD0IoaOvjdw5wYEfhBP+r2P3wDP0aWMCyMHeFQVMCe7FNgthd6ckMhhhVGmkBqHvW
sl8aunFCdS5M+8ZqWkHrWGtbYjeuCoXvvJiFrLaQm0V6KiDDm0qELYWmjuCsbLXiOj7tjkhwi+3b
2+/ewF29fPJIBYycn97+OBmd5xvPm2Nne60QOAsftLFrrZ+tOWOqR/qgH2TVwIVz4SrGKXJkUdZ7
yCzkRbAPBzctX4KAj/jEWg5YTUfwEDVu7Wjv81TAIu5c/GXV8Bj6//czW1MpL4xqtSZ7HjZ6ODXv
HiYvi5naky2FYMjLGoGIUqM1FA3iqISq6y8RtBbSY4wNhfMxqMSFJCjhNfuLIusq7aVkLQYrDBtG
qok3SLU8vvuRfvKZQvznaIuM2oyMpBIjHUWgsZoUPMW0ybNwlLaAg754Q6FwXxmfIGOeRDBxRH6O
DG88KCVFbJ4+jiSFJlWAZzocqFD+jCmjzAPHaNG7nqfneEUGL82KoaVcg0RgjUWF50ehTC1RZo3O
HFekskhI03SvYj1nsHvgvjdspCwQ0h8SNtP88QelRPjc55neBHn2yvFHXJgz4JNHqBfyXecJlPux
F5PlAYoSKwDPp2EjRGU976CmOUVZ/xzG0OVsVaZKsUicWep+Tug91g80MzlcIEy+T36RdseSXo8v
KmymklHoM+Fgv3K8523MFjOYMbPM1yfIMjQeOnhyCf/OtKrDdMZ2c7KtnNp04elCT+mUcbVckAH1
/1qDcnr1TIPoN/FkrWM/LGc6W8BGVvB2zEqBfzWJKSdaIAH0CijeddmyusDUouK8M+Xw6WF4nbOs
eZdHTMVQKNvZ6JfkVwvVIK0HUTz/tQxkiSrHCTNL0xu6vnCK16r67uLoSvgCkzLkfeW198kcAEa4
XhZ3Ajuz0s2Q5U1ArE5QDcv1puUTXmTc5Dsd//IAPlU8MVAMsteEDzxRT/96DKQH5RSWqZV3TEGo
H/B+24/R00UmEf+kESQoRXwDTQjZe1lV1+EL2Pa5IeDEyIpPtbOHG43ODPaF4SWyjMmRPxp3DSPO
Zyai0dMHzZjqNa2bO0rLyQSXNd5N7U7iWgVOouHONO2QowuUcXSU4MjpusZ872LyY6GWXT9Hv2Lj
XNTd0HjANPkZNm3kYzv5v1wY3MfdsxjH1MjwnASwX2H5wVJZ7OyvSM4KbVm3TsjrFjxWItsCtkOO
qzW/8dzp2NHFe5qRdD5L4G2GnzBk302nvpdtgCT8jMP0PQ8qsQ85jBUnzaSe+4pnM/qO39E6WGKo
6IUPHdUnNV10f/5TKiWLLr5r1Qqj9Oc96O5RB3CPQew1+xUZ8rt783TSmCOwG2ZNTQr6+mCVLSfj
to7TwRJp0+s6tp6YrqFq6RJM28pdsM9wIlTYgy27YYyWIOez+WbEok0Ox+OwHfEyaRFf8hvVAU9r
g9g7erxr/ZiXwYL44t9ms6LBZwrlgH9LwYsiWGUSN60UNwxbeGn/k1bW7ggAuM+CSyd5K1LbqTof
CJrWt5AQe1ZoTaUEYilrycVC+NJnG4yPyDZpC7qHVfLiaYLGoqRSP9/qaikxUh1jjKVY/yXXT0n2
jnEKtYyciIzdK2OPxdDOi8qHLDBur51ijgn6hGAhcO0Ki2ktuNz1xwA6rhW0c3PLOrdPHApeq8fh
tvJ2KMgacaKbTDe05ngS/K8pTXGm7nVpIRTl1Pm5NiZ365To4fUnaRt6K/b7SblalJwQwHmMw5qh
6Y87+tzKk4AyonrMLTUypEZNN7oG4zfu/y+owNuhkwiDed/zFx+v3ByiF66ZKfxqcnwijs6rG1Tf
q728qMYhhbQX2gVhJ4WPrNno83sj53EYN3yBnxqf6k0XSKrJV17CfKOz8kOAYsCw6B/EQGBR6ztm
20C3hcyf8v0yJAesNTowmNRtR4IkUoBJRjRW0kB4mKs0bPummVxii9cY5rsZeCEmtbCnkOQ8dZ8g
W+7FaSvmoPVz+/YW8z76M9mmnS0uEBPbpPlrvrVrAh6bMSltI4t0L+xasSRsTU31nZ44M+sHACjh
d2H6UbIOqYYay40V2sV+yVrbSfvVztLM2qJ3YySqO3AGbf4CWi+hN3Gnvc6MJHzPmWjBBsSccyTR
s8aZX2OMeSovNpwvuDx2f+8+u0kiajebHurYWALW48Su/TTLBuXtMA06kJ+EYDij9g0Eyle0i1Yb
+sbohs4mT7iU1kYv2pvDZUn0jqXitM37kG3zyXN4TtQ3PWX5q05tzEZOK2So98xd4kAHgimc8jDw
kzEABjQrEYNbRP7AbLyqOWL6jMVbgrgNwj/ZoooqX39aNio6rtKh5fxTgBrq2aHKBQT0iJtci8ZX
+oWH9TpvnkuxZS85jU4baiPqexzGW05qacfWJnB4nKF+E/xTDnqHU9lYRteGlxPaUr6h6bK6dkAd
2+fM/DmuTmxMy/jI+azCcP053DVE0pPTbKxBlscj6Wc0Q7hZXh4p8Q/rdqmGmq7RFcSH7zj/aGic
pf3c1m0/UDaA8wqXYHNH4ozDa5Kl3YB8hBn9ComMAdTGsopPVqKs2KNFejufyEaE3sjG9PBV7COq
YTtzP96PCx4p1nhD2PjS9d1A3u2879B/3VhYZyaAzExLgVuEd/+M7yAK4GBhJUvYyTgAanFWjM+y
L2ElzCJh50ZH7Tyu9zT/Yhxfd3NDmPNtPp2v7XaOLvaO74sG30XWz4o+XgvNn0miXHXTt04RUtsn
QRAyDnAQv/tyzpAEkEElMlM9beGOP0vjhqXDymVV7TJ9pLV2CM1s5MKChzGUUDXKo2G90SUmVVeH
XFAdpKuSb1xhdMnaG5dLIVhjFnaLw7f9/zM/mkNgBny7gtGG/MCWGMcjHZhmBiuQCfsoNP8ZkB8r
2Ih8S9jfG+TGtCU7abeKoLGXW3eHqsxVUGjU/X/FAEf5Mg0ag5CcjiTq0GHaL5HkM5Ku9D11MoFl
MiBrgkOcFAuKjk4ZkSTsRiG25NymCb0rD4oMVgn0KBlifhYKFmc+W9OzFqhOOVMqnRaKQvodd9/v
IlmKd4Bh/23/p3ruVN5m85EhI3baoF6DRIOlI4eE/o4NYKRXNHBnY8tR7RlndzVvacgp88SYJCyw
od5T55AccLeg3xG3/0QY+H9fyJdcA/4v/vta6U0Gva4VdgxAxtdvcghYc8CkR1iqUemc9M2rsu+/
yc9Q7mukV7TbgwVDaxGCu+JJGhN+istXIpnVfznnG1Nrz7wXlQedsxRTXQTX64MtRSWaSgZcb9bc
3eXOcNUdVZ9rQnYBaHrkXRbCkKDy/cIeDTMB4S8JtG5p2s3AAQCQ8d7VuunaCbgpmMsJD8jBZC4k
i271Exu7lA7ZC7pABZYqCK79fKqYYd5k1iT+ykNeAgv5QhDnFAv3xaDaMTI/uNF3rV8SOiwlwBQP
a7eDmzU60r0Mgl0aFUdy/fEGxfDxWlGTgo1sYMJIMEyxCJoyWUY5StyzTfg+urt5ujmmE2qpocfl
9jfR3wBwWf1NWBwyyXHcOrLXs+5ys3npGlPTbNdOcRKfCUH1IGuvzlW9G41H2QxWwxh/+mz8lq4+
61Z+v3JZ8wgTPEkpcVu0is4/fJW8zDvYLbF5Cm4GBfX4AoPFvXaVl51fff8MN7seBwJqou4BUzme
U/EicIh330NMjKCD9ZRO8Yt56ooTsc8yOb2heFdzAuyooWjahBfKl/Gayk8qjSDxMxVeOuFP40sx
lxkg2AW91l1knzC7AmUIr/4nlhBnHr+oZTBqTpjDWJCa/fQ+kzWA3OjJzj45+lk1tv70iEapuTha
oA8QRa9CzHHutCDso6TC1adxGUPD4UOzAwJ788cLy5ltzqYKHA9r7faGq7+iXmPKzDEV9kNxMWxa
CAsLt1HoRdWyPCXA7Z7S2fpCx25jcu/2z+OG/p45QR6ywWImWIiwYr1TxfmrzsSEvkmbGoHY23dz
YwDvmDjRBJIaDYI4Bw982/H2YA6sgovEYd0XJMQb4Z/wF38a3GfjO3EKtnbJ65Mx0DXBuSBN8Y38
+ZdoVsdquNcs2IyOA9hD3K9TUvOFNvmKci/8EsGr9LgkOzYBNyOInxwG+yXj9fHXAgGOU+ZyU2Ws
XWSzWj3SGKLoFCwfxfeihAZk8CAyFI1JGsT0RPFLz6efGafQklkokoJCwxTHc1m3Rv3SnBrXAGgc
34RnXwmu/mStoMtHzaAZ6Q25mnf7NuhGbJFdl1ioulXQjiTm+ohyrsRQRRVXy2E7flB9q4trlqoW
GN/PFKlEi+q2viLRLRuI4Rvww5jY+4ett/tpWuibscXFQOhWJtg+89QHk/+ynAuSJPqDduw6TNSV
C4NUC+DY0ZDxIe6Tm5DGt5yDKmNj/ffehodwrpRQebu8ieq8KFz3pNEuPw9HaBn7G3P4qnOjltmx
MYFhOyYjvMgoeNxCc9Ax3mBp60HwgrbSNnWWxUFlt7/n2nhwEKuNFje/baMJSzF6PfhJ7zaGSsLK
ijijcDCj92x7oRgVXZ3LDeEVVS6CMcO/ndq/y7z2GzabI0dWu2FMPzdY1qW1jxffzHxTU9y7QnDn
+mmySOsJxT8kHFZ74xxPqRwAPEY6OGwIlSrshaROtNOfm9GhHVugoFcCTYmq4lMj6A2nmpORQACR
qLK23uRv5M5KsGL67Aq5iUlp7cgWCiC1S57QmVcc6zQwzGv2yKHFkPnjG2iiSp8dd9ItHx9w+iRZ
spU0SJHZKgzOp5Az/aMsOSZDbwlKQRZLHyL7DYR0Bj9fYyB9E2vEs0KUN+ghqAbVgM6lap4FktqX
VPeCPaTlrCyR1VLE6nje3c2/keppFZDfS9igGfNbISG/QXGTkuHqxqxMMB9EyJG3FoUsu84vtl0o
l8u/Ng8lOmrxM6ZM9ipveMV1Fsl9eQoVrwxzEpcgVudRUQfE0wNmvJTiPuM/uRfXNUvPV6/j1MDt
wkjC45QtWK2lcy9VGji58KRONsUX9b0Vubwdwoa1o2/oSGYq5zVO9mWGsP8/53FflXQzJvyeVEj2
Kr3DX2JlwuI4x+hPOsPlxmFBI1naMbo+XysMZXD3PvRw1hJeCwqUVZCzjwoChDcLyjSiajNDpO2r
1u9xKr4sACICB3l+WmpXHWQ2NCYwDGA8/WOe6W4qIHs0UB3igBqhqL9Zc3CjYX+EUtqHZ6UdxGDJ
B5XUkdrBB0ZGkqMg9r0tOLlxfaWhQDJPBUJQ82EY9FsG+0JxKjKHFTsa1VQrrK1h0aB45GPQMX8C
lBm1vBpm/Bu6oBQfa4+XASzirdBP6rxUsm2Rpi+VJd8heuKgu6vhzd9abCVthLrPLg2Id9r+zCDu
LLp4P+yjNFcnIWSejJoJwvfwBQL9/lK6Va6HmhEFPLo5x9o8Uw4loPaiwHCNATzbNtIBQ29c1FcC
Tzt3yVR4RLJNXj8fNrxRdR7l4F3c30Lv4Fn/Ywxo66MR3ENu4HpP+6mtDG+VuDPUUmJxtvZkJuL/
bMGu7lRWC5eHGpWuz9IWefS33w9ua4NEHiUGavgyITSEm1Kgpwe/WTG4/92cgTvXOQVGktHz6xw2
qGrFL4Z3ESbXwE8BIQhLvVA3QKicL9iepoRFXmZbuytWuaX7plZmK0/kh/EEPyamz3xS3dV3kUV1
vjvzmYCdi7rIjC33IbTpJkhBEo/2q3E9LFNgNzTuGflzD7SccksnxS73ZmQyxB8JHyQ59qfiOlqH
IWQo9SWFKe4b3/cKwiOTo4gWR6QsJFPoZg+5RVmCBcUdOQGP3ukk8DVgYFrYfmT5651Fb7RoGXwS
pasxQeZRKA9gqSn+Vd7JOAI2Dia5S1+XTEgyYlC34R8KcaxhVQiMbMpkuKHBm9Ty0ZErpYJF8Fuz
vjdw1ruLQ0FPGcHtoQiw8M4j2endSBl8rbSW7n9gRFj0KoM27JsY7FWAEkuP6aWJRhX2AvQwJ3tk
cYq8KP0jd5m0J3cS2dJcEnsSTpQ8ZjS6EyfxYaoAv/nzrtuAJh5w6GpCwuC76hgjdQBZ0C3A2rxd
PwTgZdXYjpykVfNU1paIKs8L8ERvyhc7tajjUOgvrMmHXe1Ghp5q/wHs9FTJ9kvmr8raoBwDPyQk
KXj1HUY85q5pAP7ZxMD7rHOxv9ZDh7Rc3RihMvPSIJfh+A5FjN+7p0ov7zrFKt5EhhvVTRbQ/BY7
IWwoSGR0iekIW5VOf4jPYXqyYhEifE24a6yLsc7MDKi2//2JzKOK3nd/scsKsvantYvu0redZrDq
DEhf6Lw2A+RYjEUw8HxxlsMz9SMMJtroyylJGmQxCWk6vxAAI2D7whDqpZvsff5Lmq/p4EuDCBLd
R5tOGLG/tfL/yhXJzCgsjOJxOi118nwGecw8kKfTPLBrz7kwUKTbI9kG8aP/yMKRqI7at8OLiHFo
k1dH7BUnkIZMueG6uGJnrEpdFKNB7GUjh7/zKsBFyVhR0B7WcYzaajirFlZ4jAEUIYWlgMsJQJ+j
1KMppm0bL1xhlp/oRkh9b9doNz1Xl38Q1vqCgUnPpN3puYXI7CLEtLqUvpgpm+c1vyUJ5Gsy3SAy
Y48pH4loJMUj0QjElYIINdHqOuAI0jSrnedJKhXgf2gjp4NZTjhvq+yXZjpXr9XpIf6273ULV/ar
0+bi2YQ40UJKQ6/12JkgrSpFPkxWKk0zhwyIB4R7vKDW0v4GjIxiv4NaNfOUlSvNuUzuW6IS3POl
TeQWJkhQ/oSApgapzBEFPAJgXKTGwhSDnIngz2mhG17KDjZ1F7PT8xEfOyG5+xzta0lKdJmoqZVn
XpCBTQiIBYANffwh8KNlVArxGN0D3qWDk8Sa3iMi9gP5RS7EQXjL1nig6D99gaKFoOwOlsBkHSZv
78KN6lKKeL6ZtUOzMP+wYf+x8duY5jEE1ZkOSIhkVhbX+BfmDIGGIxq4XncTU06JFCOj0VLHvACn
60XjriuTY3Gq32xzXoSxft7YvoGCZF+dXWqaeeBP5RvuzQg50RPZ/ZhLxpDFaqzPGFfkc+KIUczk
/mJkHN2Hije41qrIX0TF5GdxzcGdLk172VWgPmSDAySZiik6FkGbx304L+JmmvPjZoV2gTHTGEJf
/SBD9QS9d+lrrpUAGRUVN1YiHJCa4yn49FVYwkCfbkWGV3qbQVp8AryOCqCamk3DdDDiG0/l85vY
mkobaDbPfeBaMyQspFJr8Zl5mK9uhHDddHUeR2K7uPPgN84DCNcPKlMp7Fts0bFsNPE5JDNF4+UM
1O5oR/EEmfoPp2ZD4MLZA2IOqSZACjng3jLq2g46z6ofkvxiI8orOOb32nBSMg9FfNl+yfWEfDiU
OVCv0yYmOdyxLOZQmFDtBwNNvM0gromj7wp1YffpmJ5WWLNarQ9LaTbVtJiGNygtC/PHL7wn8Rxf
m3GmRXYFlOZSIth+ZAryudHL0bVmqqKCaxTV1kVrpQdBRf6OZqC7lTILqkk/DAYAdFakXkW39BYt
mTDDiGoiIwKhmZlQK9uD1oJvL2JdvOnOOl/6XB9RGt12Nij8SLIK0nyt/9Llfs0buUl7bR5pFpQ2
oJjm+c+ahKZEvr3MuJtvvIz2dk/D2NqNnWFykU42P5HPmU8ce2DkD1DUMUxwzApjaPoMgWxNCkJb
ignG6Y+3oifra4uOH95j9VRJlN0hx1xtyRX+zmWbReVAOJz8uB2sj5kFX7yZTD8r88MjhozpdosY
osPyWC8KtYuZaDpVh02a1CftrJLcQXHE+gVyj3qZtmEwFnE9f5kYZKcruoxP7KRxUY9A9YMolCld
PaFfog/6cUqi0mEnztVFMamwV0Ya7CFPFkNM1wknCFkfpitQHMGuqUdusfhg2G7+gzcVseMpBn4Y
0BmNr6/pGVe4cIljO2ZxlRlo6An3pjOH9T4Yh75dMIMsEwvRlQ7jtkKumvXrNvvfFhvwuZr9ABx7
hAOeC/SQSyTbaHSo5o4iNvknM5ugIn3t6mgZozsH8n4R7KdtRyY7uGD440HpnK9py1PpBNbKq8CY
qKnntqC5UvV7W6miD3EGat+Bu/NB97GnAInCcgJ8+uJ9J3tnlt5+GrEC2KsutePxmYiKUD9OxdLi
570mKQ9iR6fpVAWWSNXOy/PkHEZmz5BoTAliEFYZtubGW+p3UGnBOFASp9fDCiUMs1jULFFSssyS
ZJRmEjpFxsh9MH4YUmCdVyeCN1WJucKyg3cxn7Iu/Yu4bOwBqoq2o79Yr5lHRHEJFzlfJqHO8js5
OLDvN9SyB8tiAjCo2p5+UBIg/f5SZ95PwqZk0jUuGZHYVReCbPGOboj4OxBL/v18U28rx684mvh/
03jw6LcsBy9ZqTjE7Liytcdg37bnLWBbjWssWN4ktXobCb7VcunNnGCnRenxPNy91UX9iIwFyFVg
WFdenTc6gwLVPnpXRqquz6nNc05sBXVrBteLHsfxtrawTmZHpg7vw5CRVwKUjD6Lz2cbNYddyDhi
G4Z7Dl0E4ukQ8cHflE9obk7wXm2ENNTtFf/qhbKXy/5Lt07zwOgdU/ql3S2hCORcALYSpHnDhFyQ
mkVdamGiSbSfgeC30GJJuvqlJKIjSBDphnuE+lzkltKZ727XVY1lIpBsZzPAjnwi+w5IoJwJvcxF
/jve2DzGOwVRP9GsZCSk5TT6/amGeime8bs0tnZwZuDkOQMPP5ta+lx2ufysOmFw6RI9Xevtfhzn
lKAAuH4fy7oGsVak2d3TpCoSKai8gmXhiwm3QJ1mYOSwLMeBxX+E3WA+U58bCC6ia44zeEeObKbX
TRcV1LHMut/z+dtyR3y5q/shgCJWdV7Y6Gh9QS9yEdZqvGx4G0ZxTUI9G/BSjoJRvq587fvwpAYu
KN2K4dU3OCQ9rqAWuDEzgX5zXYSt28EipGAgxImlrv551hz9vEwm9pVQX+Cd2KwWiYGBUNhWmVXI
LzKXljGPly3MOk3h5/ABlwXS5+IxRQ+Sn7spHyg63CW5zbznlXcIS+ENH/1jOzDdqPnRIYdJk0s+
DwCa9Xo9GetPf5Z2ztEuJu5NHzWk+1FGor+Wom28/pGjg3B74cGtfGby0h3EKc4qpALA1YqY1PNe
i871FN0N+PpFp8UGBoVwjZm7NUhw8gj+GzB1JhEh8LMXWpUsPd4Eacq6ij836S5mgVDm8LdJRMph
NC5OQacF3HWXPE7GP/XkH1cMmSDdx/lIiGKfix/d5FUfBLwBH+Ke2t+Kp3ZW4umqWIwKY2UU2nGj
/X9zWc7CtTaWoYLImZaYd4FgdGM0Mtmqy/n73BzZJp7zWAxJ2nGbuvrgPSbXSv8u55fYNg8HZKOD
RyZdMslV3DBZzwXOUnOFUxgyqrh3ZLjmZFnk+XD6AfCCjRfNkVbhvjsfOJPij1p9Y6ZrcB2Z/hWq
CU0HRLXs7BwyjzDW6vrl3S5fjM7CdS/AE8gRM99gvj/NZOsIUaypkey3EuJnvlh/Bg2IdwzxMgDi
ga/pyvXgkokkikoLQ2cYqqhEgQvc+qhq74BAUsVQNh3altmBbKH0p7PIwuzAsTkv9ltRaMEa1qQh
NKl9lKz4uHLyas+34qAqBZ+O3QHuZSsumB5+e0hyC9/2cdcKjaS8PhkQaTU3I3iW3aQBWVp+vrEY
YmFx102Mwhty+oT+sAUGvyF9VyPKVS3cpNwd4YQ9K0wsPmHCQCtGV1BTAR3q9GVhFxXT9TLSry7m
Xeh21ph9FXbdihVyCHEq0kLKwkUKBQL3J4WMUD/bjChDo71aQGXf6lmquJDyBU/YEbwRr2XKAmaN
UT0jyUCa6fLnttvafVMHWSA5EakMKXtgL6xK1X0rPJqJqv5c9luztTUpjvxNf3GRBLAHbNIhQ42y
+aHwWE6fQuxOY+xZA9ZnKT2bbBF9GGAFtQiYABj8NaZew33wmwv2ykBoMPI2QjZNCMH1Kcx4ecdB
EDvmNm8y4EFQfQADVo0skC6u82Quu+Z763BYNZ4+K2IXRe+/8RKIlWkKa9zKeIZOklusK7XZHaC0
bXdB8l6oQpvx/g+giJuQHlAini79EHrtt3Be1wFLP62YrdeO9K/+dYi0+3TKl5mxa5iQQOBBGZcW
ZWT4J3e5XGXQ5UfNjlmYbXPhxUMyin694jgsC/uPsn0I0Q7X4Hvlw5cJEab4S12+HZ+Lw+gy2jsc
hlWa8WMQ0onEObxcE9iiCv2BU7AJA55LmhqMDHMsbLs+A7lgn5xucG9OWMMlubiE2jdRiw3JTE08
p4C0bTdXPO7fMwYspcbOvcBGfiMs9LtcQy24jsf/wRujWtgPQ59oPi5Qehi3FOHv72QjMAUVu246
Ssl87nEBc9jEfH+mwvg+DDfDmJv/y9rFUsaf6DU+MH4vRDbPvhD28BM5CzNVAI+8+L63hKXhrI+V
W1UK90scJVPSHi5Fohfqnt3ZiPnsyYyK48ruhf4UB3ypifluJXfNMsUmDDJbzDIM8W92Art7Sr0P
g+ZMqU3xL1Qh3EX0RCzkRzWEHsNUwE4hDuzGeJbJrB1YM4CPTg/jI18YVByX/q+MUBMSk8TDTYUt
j5QtcYhcjmmxtLGHThgqETlOqa4vIQ+XiZrzf6spWT1IYZD+mqG653bvUvKzB8sg+z8qdLUDj7SI
dSm8bBv6cmNTApZzyp9jfn9ajctH9IwDcK336q1Bt3dfEjRy3JtyDv9LaaS5KM0li2q5dwPaOLKz
GDFUQRftHVYGw1Us2hHXt7eisi4lmvRULfL0MWxJ0wXwNMO5prm4AMleQUP2vQACdnTgP0PJhOrL
/PRan24xTsHknYYNHgtP/G+YAtaVvAFT2Fck3e1BEyqbP0htx7B/vdKnkgAdOTcm1B6FyOBB8DEQ
A0GsAw7Y6IpxqrMWMS6VMjJHha4qjjnCI1bk59ZGkpGEVR3kMt+bFE+7NJCdmqdmtnz7m26+g0tZ
Smk6EcCd+vIN1EmhZEOnU5ZcSBCq6+T9NdGVJqWFGm5FUpjOK7+SOHWT79cch9eXL/WSqh0L8BvS
YCPE/mr/cyYfxkyyFciVKLtnU8K2d3VLMCwfoFFyLdZFKkzRmK+mfqkox2eOhghnMPiGHE2rDYud
Ljm/nnCboY+aCekJqI2fUaKf1QiUgAPBEafZlk7wLB4xj8fw0EEVXyDNwqcciHvF76hyQRnx47wT
kM01TfXn8Lse34pRvdAbDujO0idxtOumKVbluTpzuUflmg83Gc9vVJin2JIwbzvOhLWkciT69Qpe
mION3AlIg3YM55GIyOMtF7KpbKVv3F5+2WM7AYZLyBQPvNnN3sm3ryAITuQK+lf44dzewaAhs1sz
crQnhoH8tO+jxTzooBbFujMRBzq196kcYxiXfuWc/q5C/rKNK+M3/xY3NEqoYxF+o4mV70MP7NGK
cTv/B3ScV9Sa86SbHScotsxTNW+6KKeWr0h36Oh+PuDbgUi/QaYaKbuh1snuSSmBpliTIjjxd2yx
uxr8NBXnb6J80gXUwRTNdYJLXwJtdGxPqoWE2/Vemr4TVtQy+LEFJeui3wbNMbZiIW8OLMfUhjk7
QnNyhQ20DFHKDSNlBB9soakGqrBEhA4WTnQvMzjrCcucsHUdatiUgE6ms5yz6vkG9ZybDyTIDqkB
/1qZjHgHjOtNsECAiYZQO52r/w+2ih7uI0oZFeKAdpLr7uwm+N3etmsx1pehPdmm2Fd0ABPZsiKf
VClpMYleQH3wZM9dR2rTDpQuf6gUKxkl7tC4uYOln1oX3pFVTuC4ee3Xor1mD4JtNvKsvR4UgIUh
W2p1pow4wjGvWfrNVAeUTS2R8hG/qqMZnHyb7uAZypfAcuNmRDU2HpXRJ8ynUV5wktSruZi5QFq7
y0LldTXGcb3gek8OuVBjEsKZKA5834DIT7iQSjEDCSjb3Sbk/3BegbS3uncDYVyUEu598dmwIhs2
yCs36H81fCRC0De7SOxO99NDNkguebenekkVhROjH6sgYxPCY3n2Wp0x6mtKVVUdE1lmuhOhVjXe
VrgkVIwGzN5xnO20Vq2cCdxzOsdAlsBws/ILCbMh5jKpKch51zRCmijTMVMY6+eTDM4P6gPAKv3D
I5yOC8XApYdOFcxwnGyXDP3e0rgtZjFT3K2SrgUK4OZ7Ss2ZAU+WtEfZYVv61BGINObKZnRniCWW
rygBgJVDW5nvYUeyohisZay2/H45aNajTHk0EOFuqWLRhWlbCY1ChUxoXE/HzP4YMaoVRubsOce7
QRJDuodnGQj1xITd7bIsyw31/msPye7gD/AV2gOd3bQDXDOPg7shFCGrAyJMwB4pJhlbmBmRRlpM
y8J3s97gsb3xRHWm6h7GwiU6w+354UNKamaXaxmbTS3OwnIZePjPs2nTpvbyPq9apaGQzM4hT5Xn
oUBKTKF22M4bT2HHYX0+UCwAjDar5XTYnNSZltlPDhhTLW954mxsFsXbdO/yU5B49Ww/bWDwqem2
uvcKnPaDYoPqBCJBAnL6aziwrYvfcP0eh1H4SkWAcphb57gqr8QjryUZG/vJTFx/cd7xzRa6ChHj
pJPk3uqLCrRaoJEDtMJFWtfnnIrX2eixJNbHMp5vOFgFXCrebTLbf47dBmBMJT7vrReDaQ2/nCgd
a/nWn1IYVShKEukFi/g2+H+Vr6Xfx8Bzf2eLL7WNbPXEqhlpc/BFDNbfnWKhv+GkXum8u4SL/gUY
XHnOO2kTjlEvlAziCx6dUiUj22E6qSokhqiCQ5uwsNHYwEUDuHr82oJDh/zMG+4gjTUGoRNA6uQW
Uibv6DkcOg2lnED6+B5w/m4hwijHySzO7WOkrA0wU5dgl/1ddwxOBdOmdjItMr4Q5J/L60Qwhl5t
5zDMvy+5Ub7UMquyNmm69qX/5oKX+/Wh/SpmPbRBDPgRNhMniytAq+CRdrQrZmeerciVFE0VnofW
kXKUOwarVQSUD2AF6hI1xkKLARMmu5P53BhxkbSjxFnPv4l3Xd2BLuUnrLTL+eKvQVZeI3WV7emD
FnuboeGoidI72oCiuM7SdA3SB/wxWiu4R36CQppe+n/3u8Ei0YiZKMZZ2pH0uI6y3ZYnp2T02xpS
QLOmD7bMSPGW0nDdrcJCirw9NZqvaCHyQoHUVJcRjMFbJd1JTGRVaqcsSG+ipC8Zv7j+wyrK2ZJT
6y1Z5Qk3e/SPVtSgcb7wycfC6bVZJi/n1veK+SSP6ZGazV5SLRwl5DqkFRpuZBik4E9M4xFi4jK2
cO8JNbcK8470LBHR6DIE5Qt4vHA1D2GqPHAuoJkZRYBibyEmNiShr9hFf028L43gHQ2rmWo0QhJS
SEsYg4Fromj41UPV+G0lXke9h7F6z0CReTamWyMRelau0zPuWvcYrdeBuycTXkuosZV1nYsGP62R
j5SgJAvmeHmHvfl8/uPhnev04IF08aXoO3xzetL1cx/JUcuir7wMmJ60KxALzbXnPkR5WYuNHzNw
1A1E+8htF3p+kGMzFv6B30JFA2Vsz88Z/dw+M5xf/zhmhYMvX/Eevwjq+tKgyx75Q2a7OSfK6xIT
6SE6yGNHQbjI3s+WEvocTcOjg72f3P99TdeKb1pD/L0vhMnkoDOITuuehGFw6dwBNWqjPQv7CRrI
SdDTqdkEEC7yss0BLFGvGruN6H7Y+qtKEAcFCFLVwyN3KCfdX3VPcXVpbXlFktNhO87/FX/74ReF
kpYE0BwhgFHFWAj1wLc+nf+pE1Q0PzF16XcuT4BUfjey5CQnbkWyHnTrEjlZeEo8CISTxiWkxI1y
9kIiMPm7ffMi0k2oomUFiro3Tx+iJPsHS4sCgLk1gFOG5e8DmTmBUYiP6nTCSU2x5OT9o8OFzpxG
uYeZs9pWMv9k/7FrstLUQPIWGIZtb0N/esKbWjt/SO4Ql6/px4jyryKo5jDDlIdXYJzjRIKPepOY
M6kRlKPVzN+HzQ74qZbEUzUA5zjcwFpfBMbVwcCfWyUuHSGlRiLzFzuhlPTTKPYmMbbF8eiCa71b
knLtNJl6VHhwqohGnVBeBgSuJbu4oC1WoCE8MXVq7y+QHEifxafXoFXrn9qwtZYaezmDFpGV6O9Y
EQVx8ChqpKcLAjYy95L6p1YsT/k0xXnLiJV3xZkAqa2NuA6QgMuq81I5X/LGQVkumdnd0V90Y2bR
oMpBdZJDl9rUxQfigkVPeAoMODwtq3+/3dF2dOm4j4Zvb397YS38fQnPooUSbuSCUVEIAiYCfe8i
vtua1lLpfclm3q0j+5gjLyeJgD7ODFd2JJHbP12ZOaQmCXvlsBgaJVpUS6RTRqxNgjcgxdzVcdLX
X1fQlwzxHByiYz4RGc0DahcL5FmBvgpTSgmtC0HhWKme8wyiD6P38Uu4fORaEvmPY4HXCX/gtwkv
Fl6nnHknzVUEy/InFGK8MVbteVW9NOXV8/CnjFkqPWoLK/1JU6ggT+pPqubdsOQy67j+z2/kfp+A
/q8uZPuEywQNMAYh7kywT59QSbNRweLcX1ARuWqFBYHsAHsUxkG4fcJD+3+Ssgd3PNdiVepMIy04
gk10s2XKzCJGVmfGAVhVtD8KEA6IiYJJ0XtRgrS8oAs1zxul2nPrVdswWsS3aZtvFjpOWMb9esCG
bHrV1Bs1c9izN8AiqPfxjCY2xYZhc/Eit8N93r/hOCSF/EmaJJ93CcMBmnLwhRLRewBV3qIuwT5W
oV2FZdilrT4Ul33fpr0P+H/1FT1JFXbLfDEz0SHg3dSwRQpmIiCgWX6Z8FjX0VWBAQ11XvZEce36
foARcVPTC7vdwqWQxX/j5m3U8pbuLdxav+LgTqFh840OjQe8WwhQ7zwyOceEkvTkgfvEXKR8W8t6
AY4qnj9gIyhBmg0d+pnn/M76Z2msAD1XR2lbtmTdrbV97HWxL+q1mRndisMX83AeES+mvwIJQwd9
GMMwPTOWZkJGqBDplQ2dUaCA7IRNuRNdhn0ebqUp0RFFeonubJPyv1O+ugEz+HC5q/QIuOUA4cQo
KQM5mOcqHTkcyZZiVv+1vrIDMjkWVQdivuMoCjcCj1tW+7KKFc4cW38A0HObrfmF7xNwz25Cx8Kh
XtANL0di5zr9mEEb0Cho4nb2Blg6xc4RFdp4hOAIkX5JmfuaJVjHlC4Nbxvu+GFOCqatfPMviHVi
es7jr6DdL0H/QgEt60CkqheDQJSL9mnbzJ0H3SfLGlN5LWtyPWIRmZaj5JwYwzavnhSoehhw7rop
tjiKoDLKAaBY+x09ECsvwxiXieBKsEZ9LqMEzn+V0Hoqi43FQ4Ocn8BF5mD564SaveTQeQKvTORk
Ok3RwwQoFSf/E05O9XnQJB7mChWlU362Rl4/BP5NKS+0n8ONWZd871LootqqgXuwWVeTwN8EJo+/
ii+F3PVw2AoLhMi/GigDkGneApcummt8qOi3/SByqS5I+V0/KWLTssobO/LKNJ9+aXezNWIEH1a1
ScpkbNKyCrXmUVV3rMvNpwJCOGd4SC+NhdDppHoUhU1nQt2i19XvUMPrB8W/vd9UTFJhE0TV78vq
w5MdbQBbSf1Meqafb7IPEdhqNRAo7ZnVgOFCOYhxBwf1PRNhbQvx9QZLTDWxVZ1Q0lDKa4U+c9pV
jdPB44l/sY1XCTuDpa++WZ4ZDumjGe552WVEyTYLJTFhLS7k2KFWU57mMxmBeFbAewX36ABLFLW/
xp76W2u9baK33veOFpm5YDMVG8d0u3bzDb9216DZOdL2IYe4teiKhJgOIK92wZf1iIqFXS5NQtWl
bjDoyacb2Ygus2G8LrHigbReHDjFu1zKcqmbkBWFvqhDbCssHoTejhPAhlQ38Gs7RPTc/hn9B73a
/UMC5CxsKG0od+lzwRZiCiOzoMSvCzXPZxrLTf6Sbfsvm735w75mY2tjjP4v8q9yrpsWeMWLvr1k
dXqMcg6MGTgcLvNysJ/eRSG+pBAOqU3yy1iIBqf9dQYzrb1CNbSv96+nSFsViRJfYWaIw5Lr9Uz3
1wxTt3NihWobjOWyPhBu0/CM9nrunuonDOQls6p9PsQs2ZBLVrbi3gt5kGI9kkqDIwuMF2GLMIJj
xTgBhywDTAduKzkAa/AxfWlTXf2QHGm40rCzWLZ+oalJGMWFinadnxV4NzqIiTsfoXMPySiTe48p
v5VOThd7QQsplINwCJeYtrxTb1yb8dH+rkz1AR0/nUrOfXgyKqmzXUg3ntQEDfMFKHxfij6ppw1Z
mUt9chRNa6P41uXk4nVh3HZAmqD9RuT8/FAlyIv3YKnW9HXta2pc/f0Bujv1fqTIMihfQYpzR2ut
lVflxuAO2InjrF/ps471wjrXNZK0DsKGPKkjEJyV2HQbJz9NUV4gpnSZzVKX8y98tomjVJc2G62f
wqT0TE22aupQkgGPdIzxk6UwkBr56rFSFVpQ9zzecaRiKDmUjR1XFTLd0wnPX1KQ1iFofjcWgZsK
u5Wq3tBJNm/FjTQJImKBee78p3K5B8gmHS/sxbYC1zuNJ99fuDl+aG9ourDM1TlTfw3cq+S9Y56x
toUZ8guUXWakRpG/Fm2OSMkDikLT76SKFbyb739Byr1fR3VloHe1l/+FA9U2h7bc5j3hzhqWYDWP
hR9kbhWUIR+QTXSzDHGqvNzj5Hd/5RS7TQp6U5TMp5ALJMFXLCLR+xgn35Qwinq1rROEzlo1O2gD
2LgJf+kvyp4E7qmZn8+BqJcCKa7AeyYf+H0Eu6B/NFygWZy8qr8jU0BA+sRAMZwZbWC0bDwmB9gq
cuDekPQJY4LTqJoruzjGf1/zNNTDP8scOkolzg0bC0cLxcQk4SnYA+aiiLh4BiIAEr5SavqGFnJ4
33es2y/QyY9IX0t8HOShEF5lOONBPzmRadLps3c8awRnzc5zmEMJWJ041D29wKvfFdZx50TGdA9U
sbvbiLGoKC/tksvopHkhWA2cTPgaVen2L2r9jgzJC3D9Ggywj8Gm8GbeoRhPnHG389pEYZT1ZJs1
lmnNQhq51nsz6CAUgK86uyL759WjJ2+7TU6dig1cRPoo+0sC7PfkwBj2iWlHi/mZnEkhbziFzs0+
QowmJbXzG35q9XQnKMFp96Uif9C3ILZvF5Y1Qqg+Zqm9fco8zMSuLl2hcFGVVi+9amze5izLTwXj
lapWbsk9WRnyMu13+oWy1doY6lYhwt6QO/ucQdfKwzMRBwSWA2HPX0wELsu1JjPfS4D81Ew1ZCPS
L9s3uElYk/5M5aVNzrTKTmp9awwehLSz8IzjIhXgW9w/BEC9UwB31y8hRDCcCep9PGSXI03K7idW
Rf6D9Pyb1NJf/9gA0jBWR5wSuUohu8MwYlJs//OWXbmkivlVs91yks+ulqBkxI8OsmxsSYSa/9JH
0nvLFJaUXUr2yRQ9HiliKAH8336p6cXjcrnjWX6gHiNCn1PfiJHsXlwA3SBAj+aeBsajaiXRrg0A
4PURu8IXKRrNC4ogscF5Sw13Kw63lidiDredEmuYhTImZShYFImgyv8BJQoO4K9fGTZJqTyOvhGw
ISebe/i/jfhpZXAjl7BkQ7H4ejN9lsfvHzJOteCEGDrDF33x/o6Ue3jH6Di0BlCMaw/8KowWNfMn
874ty6ur8/GUcP85QPfg5GoYbTpERL7cP6pOSDdhD9R9++n6uF6Qy7gVt7BxVCIL+yu9oEKox2TB
hXs8RdlCYpI8JHhtB/16JGs9gHnICTDeCEyJ+KYRhmwwBfDUIiW613WGWZV5nQz7AQTXo2bkX/dC
7In9BxYEu6G8dLfI5hgke4eNgdgR7xPnpZ14nBhRokDtSw9NaNtoZhv6ZRQq6R2qTiLmqLGqKgiC
BNi44feKfeGOFkoE8dxeoGhLsjBRIHsfaItz7p/Np/N1fM9LMohr3AsuoauQ8qPT9xgNuW1OxDW8
ApUbu9jdtPi2/TU+Frx1JAxvGy/8vlL4al89mfxwlgJfqdCIDL/3L6UhuO4NgVmkQ+g1LvBD2AaY
aqCWBjKu8AlyPP1r3tMyfnxVBhNe+hQmsqMrtCtCaDGSZpiYvv1SASgO/R/kVg84lKuPjMFyAFlc
wAq35SpFSZC/bMPnAr9Ig/wJKrS8UFKYxY9ZKzMoTu9AtH95FdZms1vnPhvsFFSwUcValCWwGM5a
rADgDx/RgtBas07t2aXOHPxfGoHWJq8hnEMpqX7DsFV7sTw3swwog4OfV8jyUraey3pl0Zg17IQy
/iJJJcf8XCd1JucVYTGNZa2OzeSUCsgbGwhjjAnxryLn8DAQ6U2jQIA6+pTYzcd1mfR4I2f9PvD5
clDnwGKJfrx5oUngJA2kYtsnF0TB5G8p9MXpqdmZeGJsSo0W1rBr3T958R2sgh8Mi67GRVpiB1xI
xoJrn03zvwiA2nzHsg9Qm5DQ6jdCQArWdr7Umm1Bk/AGPjSc+mlQNCpF+VT+n52M06fb9VZgYbwP
XinqYkQLD84Md2lxVRf3rFI2NY3zRCVLYdYBvyPSldyNlVFh1MLtncv8lxuGpbBF1Y6Jso7nvquY
vNIJh20m4Hb+Nu1egxSFVgEL9pRnlHNKAMWPFwsKd9cMu7LMG1VIf2lkwsf9X30Sn/LXPFFxTjt0
fk4avcUJ1NQiXNEyn4VsMnnvFlbtbCoMR5BPB9JGpe8na1npaboxB/GB1uSdSIguTyKX/67Se3SO
zUNJKc6qR9wIllOIrOWSMBaLbzfhVaQo1aUwn9DiVwDlcV0/e6LwrZXwlYVKfg307p8XeB4UQJio
QTAGYjGv4eJ/nqwtawojpQfIF2tkHE9mkSgM+G4RtCD/uZy73pwp3Wv4Q6vxzIo1/aVR8r+Nuswp
op79mjhXo9LZr8Y5YyE4r4TgAxBP01ewH3bkpB2SSJV3mIJhohLTjgvDU7ji+cM3GrDhVBEWdy5r
mmJZtF9rZDmZ8dfRw2B+J9jS1flOHfMrrtHuw7xwoLBYA6XlBiDve0fqGsQcvT/N0Q67DGHND7pG
Lk5lEkEgVSuIHOw+1v+c55HBIKqsKKFrXE9blZGRNrj2s/2+fpCqSoZsXJAnEPosY0kjyzm41Pzq
2Hw+Twi8bovu0vhuoJlvUd7mpuu851aIf6crpvLKQWLxPEmiPQC16r9cHVOnGzfb6H9z15V+AQjD
nzgbm5KcvG+a4iJ7XP6oMAY8VF3fpusec8BRq+2OIHcmFEUbVgPHXKMgFknSKYIs4SrWqMwe0jqk
loUFalS7jC9lk3hm6Rff5aDAuzBBbb+qgQ5elfdeLZpAgBsrUxcYz2JfwCePd8NN1stARbS2MV2G
J85ijiEl0kG4rFLUFznbrYtYImlIX3H1g1ELoSDNCiXciN6m4nyMLoypc8E+chfUTra1suQV3Ia3
rnmW8NVE9C2Ij3xClcJFZcNSNSAQUysnOJ8k40qvfT2jEX+RzGj3DgLeblDpZ6GPHi6IKdNMJB96
SD7kc1jg5alhAhbeHM9w713Pvl+HIWuBfyLkdr7tYQDieH8vOrxgI1f2FpZmqB5kQyiXNus1Djlk
hTPba8yLlE3SkNw2FX8UvW1syXiRyZik2Mjwu6pGlysnmaUgkjuutOL4fXNZgkM4Hqx6Q+f33KjX
sMjoaT/zABfd/n/2cb7ntJKMtjccwOWtuOv4ANpIoSL1Q/P4B4tfpn1Gc+ANOhIbAqDaIfbRulW0
THnwVEUHgC1xdWaZNgTqoHF8BV5rAnY5s9NG+AnZfDvqSLRSjP0X74j7wZBeZVCbZyUPhOe0FGej
BG49qqp+QH9bvZ1JZEL9t17iGPGuRCyPciy+XVNI4tDyzpFuAtG+W13V1tzNf0got2oJOCmcPfz3
UmLePxia6GhCCT7VnnSvu9QryQ83JGKs43O6mPWquf7aWTxs3GozmKZlCHPvxtkpwONPZLa1umLe
Zu9pU7FBdPyzMbIvdZTjagzcAdZjWlwNJLqs5VYTB6s2HXOy1huR6KasGVPNXZW6Bg84XtMFokZP
fKAG9Aw5DqewHSwJ8QlJ9kyFq5PSSvZRbBYOZe2NiWi+etEazNheGh/LU7GzAY22eBZbuh1lRkUz
T9gj7s4P2SSN1aLvGjfGCnJnA36hsuOuBwckJ/CDqRDFemuvKhjCT+Hlydj5LJOxUrxX/EU0gSSh
iEaegsthBTDegPsItUKP68NKL0jY65JUtQ47rml0exLOScmPxTlIDcYEt0n1JUWZIC4Ikg81o1j1
ccuGVAlNzcRGF4lVW3ZouXumHMlrNu0UcfZChbuh1zNpagonzk4dyz7B+n4Wamc1w5gfzWySx7Td
toOynLaRoreSnF7+pPAsVZIwjRguBh5PPbGL2rwA2zu9sRpbt8cJhIxcPsAJmWHaX+bq+Sfhdkut
m/2a0Ga9pqUgSvoh2MYGQUULo7hxNP61BD+2plaPRa9vzfGHrE3TnB12cUu0vd5iMC7JwyMZ7egf
ax1xOTZ3Tz9qNN/J0AkQlxlPAnrF/Mgv211lxz/KAHRKLqj1Cb5glOK5NOyuZzrtRaW6xO1q2YoJ
gZggMeU48OXcx2l+RvOPepG3XNHZi6JXXWFl1qZ7u9zb2dUO2Ku63473zzNlxn/SkVFsYrz9zvLd
nk45YpfTdUSZLl6XS1fmGpGrVTmS5oPRZDNXZiXmYEVOWt+Tt741qK1zUi2QxhcwNiiuABzp+P//
dg9EO9Y7QUSuQnJr2Xgay6lZ7IL8AAao9f8CTzdAoszK2avpr8gD95md3JvI04PsYmrJjvBNIi8I
EgvJXeLLu1ENgY/UM3DdlBFOmFS0HZWSjsB8RNps78JSFyElRkHe6IpTwBKFn3ECBRe9G89PSrR3
KIMWdkrTeDWB+g9mzYi1Ht4QnS0/AdfN1OHUmL46xR7+ENU6qbnKG+ZU9pAq+gFzx1tjDVpyXXUG
uxB5UW4A+8wgLY68YtSpjVJZog9O+rcBTb5Dx5vTBzkP9YeI02plG+ayk7QJ2b2MjuF8OdAVU8UV
LmuMdjfRR10t4oC/zMRO38IXo9VpEizHpRDfxor2TjCaJX5kQCXDywhNOujKB6p5U7ptav9P5YrS
aalSPbrl+zPfoZQNy/h/taUpY22vrLqeEAIM/ISa7eOnKrYU4mTA3FIt0H9tGZ2zbOOiTDOozoF5
NhomCbTQ1mUVShNsAWb3j8zvpVz9AMzgnefOBASES/bRrPjIS8F3v/2gmUqgBa+GBJzYC9Jhr4in
CgaKJWJfMa6Shh6TB04Aq4Ye8e574mtYYZjZ6lv4NDNW5gOKUPL3lPwj0g819u94S81OBKYJ0Uti
yj6q42vf7Seuv+mX/TrWC7DuccwlxYRJb4NdelDvw3tB/3SMy6lj9tFBlgWCvAkSvKOTDDWbOWfa
R69W+qYUSujJ493egTYRTIj6vuTub9vcDmqDHVVu7JfjJMBs7J/OfVttkaHLhkPgmlo+oSEu9FrI
OW1Gein4fDDmVdnS7e4WzDdNlblxZO02tFy3JbpTDWKSUrbIwPHASJzGcUXKe1ZeX3xETmjWw/59
gx8DJrI9slHPy3JH00kIhv713TW4CMLiLN3Y/JDnKML1N0TWHPBLuPcfyWsma1EbN+JVVcffekdd
8DVm4jK0f4Ar77A5i4zDLkz8VIVAF9IlwPpujU7gCT8PzBxAECXuOPFD/plpp7Yd1R78W1kQDLRl
YD+IofJcxxjrQ28cnrievjElddjnPbqoR6k5JtgeSkw5qeeXN0WXMlvJ6sNuKmMGFB9Ju8uPq9RJ
aY8Ri/6EALiPc4X9KpV/bLeWbTCHdjgyCTH9EloDB/4VHlappSfXLYVC4M8X8ihea4uN26cwfRAu
gsmHJWJonvwIcpvOoqmeHQhOp1DVI3mQp59uN468h2eqPkKzCFfzBHGbZ63ltJJ1BoRR5s9Ci4AH
uRKf7RrRL8iI+u/2XFpvzCA+P6MkMTfKv69bGHvbV53f8RfxzAvt7LIqgFfrWzBoGnhZ0mykzDNM
+rGLQzcNwH4z9PBH6QZN4FT81pkVXHAT/JxDo+b4L3DsTmhiSB+85AFtHW7F2ojeyjX4Cs3Ggl8n
ca9i9G0HPNzWo6Q7CKeBUFbdd8VTx07yJMIar/wOkpv3iVEbG1R/iEKxX6BRcdUCiMhXBVaXXrlV
9Oeh8CSTZVv8eKJPFxmJunzAqjpOq9IJtVSbrqWPPfe2uVx9NeNGgVsjqKbm9ed4pV6aa4pNrHTx
xYvSG6mi7TySwXb8Wvnq8d4CtIKATYLKxpH8Q4L8bNB3Qpdpfe9fU7zXJuSkZLQdA0/yGeC7YfMO
I8V5OGvm4L6hDFrsp3zMbgD1FS/dl/p+Y4CmV/WaXChlicXYYfGFZwRPwBdLAZ5MfcWlI8Q7esRG
d/n/A+WsTNB0Yn2YPWDzm3ic5h3+mUeQ0aT5idGGnsFvlK7O8oYXP6AbQqO5Z6JJ+k0pjaVN/j9f
c8MPL3XJ3rKepAtVd5j7D9RZTKk+zQKiEanvY69O1K07lL17yxEM2te0im5h1/04yic63JBADQ6w
wn2mWeyYk4mYGZLli+jtPDua2HacPB97AOIvqoxmL9g+XsvM4XCu3WsFyXNISITovHq6yRIYRbtA
WHY2uNFWl45+Y4ikPNfgG6sQa7Sb3VoiqIAp5qDlux9VlRVkbnpC9nASshE7UvHrgmlK1HX95/xf
9SkrV2HmNaTdWMbnWtIZ9to9v9lVRHwxocFeSv/GxV+9SKecykTQK6RLDOvBN/UOXXYx89tJzy5C
tHjvzfTL+Dgq0PtGXSddpwXqhO5wCfFTTVJ2M0VXDCzKsq3cQg/8ueOTKTDCfipZ6h1krPXhERBU
b87cKZj127RsqhsUw+Blp2HpNA8cxaGlTA1RWIRcfD+QXnS0E1v3bABuqrICT5GRxM6zl9a5y1PU
RKSCjeAZHgKxZKzaVxIn/EbZ/rCAXzPUYXcVhUKZjp9J0x7WynEecYoDPcia2tCasP7EsCO6FJGO
R/2UdRqqRPBhCllxirkcV+z/5BozebBuYgKZkTxuw02P3lnG0aeYupKfSQutRCSY1s4QtME1/YSO
A2qY4TmJMF0F1283JJZVgiE8W2i8c9X7Vj1MOwTvBCuSjSQcTCvehJPCED9KxYC8ES71E69GYLNG
mV5wi+tIbiaqxsUaTucVwSfqlNczwrw1wbuT5HudsqmUCnVbWbvAEz16263iGdFJuMqnvP4kV4+c
nLrws5fpi5uvQi5tlMPA4xnE+6eBNt04H8hwmm85U9FtinOWnVyOzO90SeeqCEj1EsRk6deYcrJQ
/f41HUNkO5w2tBIckKdEDy9luz+HBYA/vGEpjhZlTmu45Khc2UPigTu1oOk/5dYXhX6wQ/63p8S6
JQaQarBDY5YmZ2dYR3qaafoGnFffEi6LehVSzasEefuJlOMXVGXaWnZU8n2AN1vrbIiP2tZx1ZUf
Q60HNFdRE0rDwnxaF9ZEnVLuGCWHNAopyADcVAEyik24i4tgw1Zxpf45w8gOcxI7a3caV6lf31Us
ewQVJ3QqAbOMzH8siWcw8UHIPWykhT9jx4gHXG+5QvYNbLR8zpJ4nDFT6bZ+fYI4RWSIED5N0i1j
u1Mx6xsJRyHprpPc/lvP3GaprKuBeie4gpWQfB6acN4cwGI99Q42adN5Bhtj+W8VMWgS74LjUvr+
0VHYtL2B0Im+M2TwLjppg/Am1rptvbhknTR2jtia6k8DSdggAbNktwtWgLM6LU43RhpSA2ws+7N4
OFtbvce7PkkTTkgmDBCXejjxQGCsfMZXtbb7NRsxbj06NmRHBwKal+53WkKhQ8dYP3wQVTcLDoQr
dSl5jFCvX5POiZBE2/ozyLmgOK/udHox3xkPZKWp88rLnnYBOX/AJlzlntrLgARUTwnxcSener4V
+5SvqhmANFCZBV3KjLaoBs2rB4jCrx83CtjAePKvPTGMdiYQ0gpf5Rw7orm3ZKbQSZ4F3wgCwaYq
m/e+TkGPYOOYp4kSx5Pcc3CLZ7eZchKSZbdDaLNT+xadfQAkkI4D8dvOKA/WUBz5a5valU5AuYGs
JMqGzMBEoJzAkwTgpbNG1EsnfABRWHZLMHVjwRfSUz3qg9cOuAEFUCTwrkOm6VpnEehDGzffpUAv
nIauZbBvOst7rS+RkyX2XQ8tJOvHNAE/hHVw7gXdWrXP6N8jRU1wAFDAFfo3RBJ0xvXSO7ukgdh7
i0bY6uigacVqg0fr2hIvJ4rIJMtn+08jbVC6Oa3Yz2lB3kzpXzjOfR0P+qJYAdgifY5St8JlkdwW
LSdiFMZBxrguakkO6t7+BihZ73XEpHuIwB9zXCs52mvgC5WFEZzivAshQeXhNkQuVoYlmcLnTZfM
KYMvNbCVmiiYbqDqlEGgIj0IjYsYO1+7WIGvdIXde5AkeVY+ct3WzO64W4oQM/IJd55CaA/r7Q+c
6RF46gHYCoWwYuRfCMB5nA2IqAe12ksjKU95XA54BKbu5Mqsa6Mo30+67JUyswyOxwSOlC0GXd6r
0V3Tall+SmQJ/6Yj55L+PbC2IbQyrdch+nrPi1tn4SJ/3ZucY/oklfSOmrP7m+48k8UlkzjC7dXT
rrSbH3+HgmVB+bgJF7dqkyzucgdMun5rquQPq6RAAjohBw6ZPJ+lihyjCwWtUYUEBmcnt/epHH7c
pT8mfow0za+ii55PYQOQtgvMcpIsZTawr0red7SNGEPvRTCROqbA7GxdK6w+VEjxdSJ4TY/RdfTQ
//mWAR0CvHFIz5NWy5I1Rlu84MbobT/ptOfdunR+exekQ//rIWpJNutLpDhmrWtczqiitkJwrLuI
3tPxvP3OmsjAjMZROEm/r5qF1PG1c5hYZVSrzAa2NyYk7ENoRC1tIew2m5JOliMlz76RhGAAlZZ2
ItraxZkg7HiTTNPa8S8u4YQJIODGLiIooXpgfdHZdHbzAQ6Wsacv2VG5ZvuN17ipnCw/eewTzqHi
qAOCVoT4Jt3WN2o025oy5aqSrLB9dR9hodOxqkqGE0RfLZ+PO666lm6K07ZKM8VkRTeFK7XEay04
6PLbIOeuRjoREu0UWLinS41U8TAJ6Il51H/iBGbOrR62AatNkQKIEzRhtzYLLJ3cvYhbKWihHAIn
JtyM7MCDfWF4hMDNn02u7VtIWHp4z3TLLCDxYFlQ+zTK3PAn6IIFdmBnVArKUvwWXEgt349BwIom
gkQvFnOhCfz3UxuBz9xvkGPDgTIxuhaIhw0vSunUNVoMPAgztn+qJ9bFKG6d4AA8E+iDR9ZTPVWE
ASLAZuZ2rQ9I+9/tvq5intRlBn8gidvi2hUFUfuyKJg3M8QGqMaTsm+ZfIWP1JMZTKVW5P2gWETi
6V3Ypzze0c6G+K/YJ7GmQua3VYTf5rcNWWP8XrJ6sVYAdJH1hIGAcalFc7bgaq7QYq9axsJj0d+V
tGB/mmYi5TTMEZ5Uap7vMI+MyeJ9DWETiC8uiiRXXZn4xXViGFJSepSl+p6S1/a2sgJ7evQI54Ix
OarxP2zXx33/z/+rkVlNl8wYPjvnxm5tGIIf61pe7LLU7SAKGWOWmLteBIZgRJFilJlKzGVRM0na
j0mBuwb0XhwsM7gjIpDc8j1DbAZV88zD7bfFrpcYIJzeN/5ke1OK9JB3y5Cms/Ad8IFLzo6H7/ml
s4l6XFGduSrVZnl13EWaxXrUwW1ywA4Ckp7zX6WEscCrIiWQeOzfXYt8Mb+Z0k4jlq8rppOEVAia
DSVlxcvSaAuZjuE1BuCyZxyYayNl5IgYL4an9CYOPREflXl6Mn+ipUKsA/PusOcd1fHZYlxVY4G3
8kcf9X6jd5RXhdEqqEBIlWzUl9T3O5KGSjfSkzxNvTfMpq+FjXr+BKIQtmfBtT7ObGErE8YnuTwf
/b3LbculsPD+VeUkjte2Vwh/nSsOZx5iYArzuFVn/iTa0gyYIP6JQwIa8X5ousIFZJs5sqMgSU9n
iuDlgn339lAoKVMvH19lwi75p5yWBzOPrya81QhUS4SvIoLcWxspsoHGlOZkk6SHzkex9V7Za+aL
NIUN9g5HogYIzzzACBnlC6+WivWquAGDYEw940ZzxEAM/AXA9FKjVjajbV/FSdAFuQbKeloOEmoJ
iH77285sXToakUxvKHH2V4oQFdFTVdTiOhjcg2FaoKKGJRVpeQW+1aDhLlNk9FBmm+zJWNok02OS
/oaLDFhQnzKwp/ZHNk37Nr01/4D5coz2JCVfI12tt/hWI+KOhlpuulssPIdnhhJGmTokq0DYZnrA
YxhumfDZTrpEEUWWrTCxoXf6LCgMtJx6XwAcv+shKOJVb0AVkxKf+moYvAP18x4C5w8Zpn6UG2J/
kD29F9GbaveeNEzYbe3YZyUKuuQTubvycmcJBaIQwdUIIZQrN8hac350YxiIM5xlPhWcVwQT7fkl
ON7X/dnhJmfrXcYj1rreT/5g6W9Qtlf9rW39A8pHAbldlp3QId0xdLgTxB0DrZHhtMwzpeB6kxYq
2iXmh0C9jcNmGDIx4+U+YwjIqyU95aFlAwHPG4bQCxUcW4b4LAvalbIOYCCeYm4zoc81NSbY9EMx
4bmRVHKs5zRrqdDMklQH1Ltpucd/s8VWCnybecTRJBrL/jv51PRh7h+142KPVbjE60AmfbroDJ/1
5qL7Z/9wbRa+zG5ARmFz9YC2V+UYGg4RSW9eJrrEnS+1w0fMCxijBVp604Stusm2AtyE+EwXuRdw
knxmKhFc63NrBtt3g9v+4Nbjg0p5hz6YAxbeL91QmVkbLnj//hN3t81F5cQIVMRbGMsDjrSl7lJ9
6FrdiijP9hgoemnH4yTH15jGb6Ub3uKQTpGDku4hQbFE5Lf3qGpBdgIkkG5MTphQ95U82zqLDH44
5a6WKDajdZhTS3+TiYUC9MYEP12rDGas8aCI+Q2PB/EyQYAyML+V2JRg4jDXg3pSxj+S7ifCJTUD
1jxb8RrBi3J7PBRP/aTzSOxUiFwsJRyc1ZSGvQs/cpIGLy93GeFzeKac8U3hnNJm5qfFQg+7nXYu
wpWpNJ9IyDBS/opy+Hh5RxuJ+xHUU8jqBbtzU75Az9dPAZrRv83ToSy2xIAovjJLRJMEiT3DZo6e
jB9RqyGi9gRbKDHVnM/C17OCFUzaSDmhX+8hA4M5RGWfNsuL6JN80q3LDRhMDDouHWu/L7elZfsz
UfKph4EwufWYcAYf7P3E8YAN0B34+ZPZKmoYBLTMpl/7k8HtzcbahCjZBegxtzW46UGvoasfdJ8l
2WWGS3UrLyFU8YOAJ8qOHEgR4cxDzMUCDbSK6KvDShCkV5aXHPYOe5idPi4ib5k4z01XVFNIrDMS
7uvUaIRb0ZTpQMTlwwqqTOqmJ+u3LRdeVw/gDytx29SLZU4UTkFyIBI98qcRK+gZN3+5rADZ+Y9h
ScRSo5exbihvU1bjK+STcnm/rwHnO7+84F6cFN6/jPQuTq4f8pcj979jx3J9S4S4n0Qt6chWsgn/
xlPIKIDz4/v0I4nsZn3NdqD2gg3AyYgB34QWr65fe9pnB641JnXHnk/O/zjJCCqwKrjcg1oYVdYm
p9lhiGyoSvKLU3XpHNWtcBrwrQwJpB1FVEr7Lr+qMedcslHSJqs/TwvKO2g5r6W0ZwKj5kq23MOk
+nxjtrKhoI1HWzi8Nh38dUz9KTSc8WufJCrt1I/3RvkJiwUH097idd/GpXMpMyfmrVuWUx4PRF+A
MFmtImYdNsL0IBawvsloIyFlvF986VL2/GDECnySIq6/zcSxj/loEgtIb7N12vCUEsJ1cPJb+16t
5iiQeIO5umsGjSQvnXebVjDbpIPLc3GiThCM2BYROSS7iFlpNDMaoDx+u5kW1+atsDcZ0Q7JrYN7
X73nJd+Gypv4R4cqKj0sSzHar1EtKEWgk25eW1iVvG00ABEF2lM6+xE5WY6UPx7vwuJmEauPVmsg
pXM0U/MNUIfwARotasFZc17ucB3g2NomIQsLO/7E4hhQNUrdxTAU8N82j+0kzs4wd/AdtHL9xXQV
69c2jHMKmyhyluGiTWe3yoFyfK/oWXaBZLHNELq5B+5wf9eTkfvnHGI6Ximmbs0XNDxL2Q9ky10y
w9UvpoClVtzgMuUkbl6uUth2HhjEkJZEW2vc75Dl4RrcseZvw0IxrA4R+9gCkPnmQ5MgMYprguY8
iDg+I8174mRuc0MTtUJFCrJXBxvHKwnyi8FrOisT7ZvJgPxq8AISyALC9n+MIfg0o26Fe9smq7Zx
VVYu8hzv9d1OTFWgMX0yu7/hEw8EP3dS+WSMDZp8rt/I+ME0vW+urXj7LikuHtVKMcFNWyYMI4je
Dpdxoi5J5/LHseIZFgzrVtsDEaOpDPm10ii5vozCttIR/Zr7XgLGINl2TH/83L7/jb9U4CcY6SnK
XO7DgP4NaQjN/x762imLUAetdBpAe3PHLi8vUgZ4XWM9bIgQVAlPDN0SYMSt6A2mp4MxczyAbG7Q
+zL37HWbP+9JDo59uSGQvGEGK2Gu6bE9FY0vtAcJaY1W0kU4zl209tIhI7IUqkpxGEMjEwmR/r0l
KEwbexT0ydIjDcpTp6GzreUBMQGP2id73de3tDh8PunD9aK8drO+TYgvG0/gJ3pBMgheGWj3PTvx
QPKsa/Z9YbjiBF1e25nArhzdwV9AzI5CuO1kunG9JTOEAH+wpRhR/+mckmxF5IcZkbtigALs6e5a
HosKVL1i02388317wXBHwKUogMsFtRLj9Ji4sk4MxGR4AF9+jlN21r4Kl8D5y5rvlL9hkHIUE2j9
KJOFd9U+S19D2vWYELd1A1kbIWZ9Ub76dHMzbuWNPqKKghlp1n8Uv1EYqYvuqXRMVel9S1gOEym6
Br0PGw5wN588bEmyCXMlG0IpzJOzda6za7prSnk+8xRwepUGFQ3YD8WSHjKGMiB5DAqhjCGuyx6h
KJVzsSgrKwBBCpOUCYF83ZV2FGmClisLX37o/TSR1KwQNZNpk2ANoqhurdoBuknuw7uH4uVMyL08
TC+bYUNyJc/SRzfi/sCRKmD78IzJODTQXTZNxnvgv8Zxz4Nn2VbjLm5L0ROtzQ9DMdFwS87oGhUF
iZaS+kOKEWHCAjrPcxwNu08Ae4KCKnKaZMX60bFTmmZoYVCWADl2NpvkLtOWmzFncUvB3WcHE4Ga
8RIxPGW/L6gS/+Qn2JW4L34g+ayM9sDle7FAA7ppSF0Na29q+lEc/c3ilgjxW9xN37i0NgocV8a6
dG94j6REhab4xICF/g0NUaK8Dl6C0c7y0lOFngt6cT8DO9aEjdsfnrk5PfAD1xDU1VSTOMBr60kT
n3AmLyRGawqy3Lfrk1wdxwD+Gh+LX3OY74R8lj9TZFXz57yqnGuDEwjR1PRkswgnWqSwBPOHPY2C
R3GT+FqF58ZmAyMEuP+DC4ujS/ve5griD2MWqLfcoFpmtEa6GrYQwak6/FOy52/ZfjfZVvhkj2l6
WytXvYiRmX7AfT7e9+Upevgn/5gXcnId4Ap5PDCInfwN4QOM9pdz/cfwJA5/7XtPmHQ943GN2t+K
n21FYWf2y0Ischg/K0P32SuuCbFTBJZpbzSxqOpZuJiRZ7WSYFYmMzFem2jSlhsVupYDzVKHBMdw
FzZV+3ruC4Mh2PLYEd6nJKjs85zjR3/lvCnQRHkzXL4iZZhFwXqoEpQOGZGQdk77ZydwX3pRhwXP
RCtzBLTCCR+rjwswZV03U0Uws0+g/DxppOR25ZFgSvEKi5Osq4hJMIQ3c8XvRM6lo5hgKbgVi0Gr
j3Wl+60eG0ukL3Vso6sYQYshhOAI0aR1HFrvss8MpiLN/WhBJ8CRJYd2SPOcb/HG/LFflN8ci/D7
BeG9/sqCQitemPgehDTK28nC2sHT0HJNxoZXT3JraGS4a5WKWflJvDOFxzjEs2L7OtqrR+EnqRu9
o5WrA9MnGq56hf4bKUkqUD5VeVZW8ZEuBpQbUKB6KOlMCpxixS/sd/owq5ZT02aEriJdZKTeDvDm
LRkhWq1TeL6v3T9HUjM1gM0JkGNSlewjnpkRkHpwV7xqfg4iEsI/jvUGY6WlxOkGKjiHIXJBXQS9
15x37SEP6NODsLy4cxjylcuZ26FE1e/hLizXwL5uNbsOrrfr+ue1DjfPFVoYCPZVO2NS2x1lq5x6
1O4AioYEYxPnNodS3EClg+ev/zR+3MeMmWCuHXLcNJJ1UiOM4ntI6sMcvxf3kbuGg9N4mr7Dpd3G
Y6WADnCnKGqLxfrVBQMA5XaThqTxUh5+z+Dj8ELvqeKaRszTqlq9JAwltZ9BI5cioa8NfrqQ0dIw
ZqbnMkNOBR6/w1ha3UBtcP9I3KRj9Zt3RgC6jCNy2O7fE6LIaqKX+D8Plw7sujGpi3WjfPdrFzVB
zTLmqiFng92Y6PMewg9UZvdoR5IYu2uVybEhMkX7aW/tRdcC7Xl3gB2Wydq3IlcQE43veZ5INfv+
3HV/mQhRtszhztfJVSx6LUAixjbB6JEUt0FrrogaucQ9SKWokBWjypm98GwOEUAo7aoHRyydo1jc
kDoc8jyhxrByFdNDjuWCcgZAGNK+Rc+bPGIG9HLWCoYopVq2alJSF0LtUqWckF53xTB26u9fTuqT
nWCr2xleshxyKZ0cFDN5PdZMcoVSgfQXBY31k9/4jEZl4dpCo2WpDKNe+DLudKW5u9A2dhADqQWT
qiGT3/oDMAsyYI+ZgrxKc4FWqo9KZl55tGXzPfcrRaQMgCvuIEZZcpaZJYqUwgoeQYFaY/SLxZop
4cF/M1IBsJ4A0R2Ga67nboelAia0CGxGdvTz5G9MV2wdglyZKLrUWzBtjqIsVnKwIhQVb10N48o/
7yn/hp5wfd45jazRaUCmIxI/O9hjQq9L3fHXAtMgNt7Fjgd6RNthQLgSsrLCJH115xwPnaUtnqmj
sBvFsbc+XFIAA8IrQOJdm9kVRbwH0ZahreFqyQosPqTpJqUWOLqgH+W55sEisYwMjq0wSNmLpjw1
oCcEjvAD2A573ny9PbrVpHMTxiXb3LNaqazC0hM/sMgOXFYOJwQEvNYzm39rLrsX+jIShmfASbSZ
BmAex0vJ3UmmC14wROd0BaQyd0cQGLGxiPdKL/6Ra/WihG2qOLW0ALg3HHrMrjMad3wedUhM+3KA
O60C1bYcxS/5r9pJaMXddZ6cx+4W9kjraVGJN9aZaFWizs8kS10Nsf2tFZRAaiNMbScAbBTCg8J1
TQDhuCu8VHFP8rqoUtQOCwY3nIZBVORsQmxpz9Txq1AM5EiAqnTR2txsmZO0fDyMNPbqgJqwTPeW
EhA0kkWMJQClX5Aiq3/6sBzcCEfzsrVptTtUwlHgTD6Xp0JuV5bS3vYiot2K7yw9i52s6gajR/nI
0/TSbzZB6kRY5ixuEYjxyGTxhWhmyMuP/yhJVa5yhYYmc16cu8dCI3fPr8viktHaVE3KKtTvccxU
l7GVpaW5xwNqhqxwSEsEpkN0lHclsGtEF0c7HA5zu1BB/xBWIRl6k3rr34mAQxog3jI9HabIVRW9
p1bcQjNE5Jg6QjAyZj0VjwoMqceLS94Z46Hz4yp8zERkiWqoJiYFqYdJDDUrZfGltRrOmcL2w9ty
VIfgHS/t4hZqWlpllqHxjTjX0LyXYEe4QkZpuTiE0ORQODzyY9kJdFPLyo1+ub3eW54JB6rslwy/
f/U2tx/p2aZqc6lEqPE3aQJzBtiTU2OIYNXyhnDyVe0q7krk39O7emi/gZf0DyFA0Ii8HH2jSvII
ZjCFMl2wpaUxS2UC3gYXmsk5m3FEeaOVmMMHDHWTB2xk3rxdFm8UlJmcwLRjCxV7V1MIBFnaOQbw
CgmGvKXiSgXC8qh5AAtQpad9ipOC+vb7g0Q0DIWNtlVe2qW5vLPn6opeebbyoeY61hha4FVfJmWm
znGD6YlJ9TIHsi3ejMMC78WtUpiwXlqlpS/RT21JhsN0X6jvIM7f7qvMUvNgMGTBpnjb0Bzxt92v
0Gol/mRzi60ctzDPpgpE0pnjjHBM80RJ8D++l4d4YdkrS9CU69lASEBQc0NxJt1KuR5dErSBV34T
T7GCC+nsuLqWA4ppf4j1CFySweBGVOL6sQqU5uD3d7h+m+AO73hw6eKdjREJQjuIabKPiGtyaJtJ
qWuGDGPNQC2J9dRVoJ2BqbZmHvFGVVJHf1+jDzAt64qBs1PqceJ7WMFCdp1O8eFr2mwFIEm0tL9c
A2JS4PdfhfiGZ0sN9zbrpVpMbxoDO8RPKHuytP6ePWjcwGbYynt0FtPfnbcfgfEotm/DQnCqs3Lp
ZvaIiKSQhri0nuiWLmyQu7KfJYadP7oPeGwRt8ULo4N/7ClKpcT46pBHOn3mFNI1SO+nNs3EdYEh
3SyTDRntNebAHtGR8HFCoyPlTZGZKXwS8r7NDGNToHPhd/5j5HAS08YFPRNp8S4QoWUbqaM6/9pM
LUAOYhEc3H6PhFPKvcIKcWqpSOnUOr+lHBTFpzETwf2wZEWevMOL9fN9xo5WiCCgJuAxxs9NFHO9
EwY+vphvTL9yX8u2hk0zS0X+A/8Y1R57U7tVxYos8YxTZH/lCGscILSG00zVsiOuJjp1WHd556xc
yfqfXk970X/WMw1fuSUijvbf3D2ZDD6Gf452isw5fa9oAMc4Bdj+3yxW2yL2VZ62yKWbRma4Z19H
81TyfM4LYcbucgWWosNCA47qKrf4v3rIPCnO0XDxhVzShaqMkmnYD9eFM/Y+PitB83FTlkm1Sr8a
3PGuNPoUXxrSuyngWfn9vvoni2eRxT9TuUonJcqg2tOG7S3uL+MouBRVGAESCAVsm2bJCBoUsDpn
XpEIHXfo1E5pymNT7yI5GJMs7Fj+TkkCSqmpxSfvy0D++VFDZMwQAyUrLkioTbk7Alfqg1JCHe3G
hyDJD78G8KrR8PHker48b96S9OV0xji85xmH2zUWC/UhH75JBnxih24Wc1+Am+sJYkZ9MLSzdh83
+7YMhgNZAcqXDtIDHOCUmdblMpDZyQ1w+6P2lm60+gqFArw4+1CsXj48ZYFyjWOHtarUPS5w06pc
tYJZ+N3K7pTRAriTj6E5qg2xYJP6AB+ZWnWnvnU54wwJQhlJvL0SxdVNGuiI0Olmme9ETkJfarqd
jyWHgSJfdo/IXMy1jj+bO2qO+yYiQiRBsAnj6W0JOebKjlbXJS6wANAmQScaiWjRnTGxqdxz70H3
CGB0oXG58DW7MhY1yJO8T/oBAi4fWAc/68qLx2fDczpeWSdTr3qpsLupx9uLieDkafuTa2X1oiMg
GbX6reW1b6Uh0XJq5s6hM+0SzB82iIVAfL7RBuYzip5y7lFXSeLQB6x+MdVQ14LQWDbeihgIBUVO
HuVzDhTTF/KA8T+geH+/7xri6xXSaoqD3EHybEoWym4QQPHO/UqrogS17nwIeYgEIEi7n+YlvV1g
EJ64o+3NSK7RlIInWvhUV1rzXpPlGT9IHXETw7dDS8Js57LIDIhpumadDnDSf8VlrxlQ8nIAozal
5qguFA353XnhBTLaqM1h1V493jX+yT6KULOP+3syW655nlWXyrzbaHdbIoEVsEWRlWjdIhtY40AN
GjadKUw1TwAy8LUkvE6xeRR8wyYnctNw/LfT8VBjEzZKUxvgRDwAASTN/8e4cOLgu7lbDRAXdRfH
56N/BlibsIX+dX65NTwyvaNzrsUmChAc68wRAhcOdOS09fFETu6IJn51FaJ78TIaLe8HDslM8lrg
MWfE8WM6gvCyUxTy1dfuwPiuCvG+XtpD8MUDyzi36Wp7c6WPLadbXygGllGBAbwb51sn4yJBspfW
YQUwi9xR2F9r0Pev4drI5AnFl3t0VmbVVHuA2hvzmddFdZd6NDsWQO/KTdd5z1TE3PuRmNCdTy9p
08M+mNLNnD2VMRL1vP5dqT2ua2PINPWu+uXCE3FzumSPxNH54ES9A3m1AET2tE1E8U1rGslb/dNu
3978MiH0+7gMKlGY/Z8lDLBbZRQDGp5ohdvC3g3DDFle1rTQVkdDE1G77qZo2mOyg1P2lTx2NPRV
bTPlRPRHZOEy42Av9jdxdh2sc2yw1L5jb9ZUaz2lF2+vmVLo7K+tE3+ykU9F+5NUuJrRjDrAHPU2
aT2rQxd4zVo5DLFOpb74UDC5xu0CDXi1BPo14maujqZ9AqinRke+OXj0+osXtuyfxrSTbcfF66cr
fB5nqECRpeEzoUi3TpsI1k+TTLK0Fn86/A+cAmajUhJGuPzkR6bjI6PMMxahrtNOKy5OYbdgTjIU
ZEjzBQtZz/LI7My44SoorZtWAncFR7rnLMEoczKa09h211WgvL9j4bHUvfyjOTXOiQhx7PqvgHgx
RjdhjAeYUljdHcxNS/kMZ3d9coTt9dTE4Q7TuRHqKZtHbezuMEXts2kmsss1Nb0Z9hJ6Ud+PhvyO
NydVRqPZGAk68PYNQMt+NKg9AHDb7tX7xIiGw1hz1AyleMSK6O8/re5uc+g8rM7+3/Haihxs9LFX
JPTZjiaNqel3oKWYEx2Mj68Nq1atzs+v2Tpwoloyzf7DZ6nPp+pCGzQogK/0jnLJ2hCYc/PrH5fn
rJxyfKc+DwuSYz/4PKYNDTIP30ahaEypEc3CsnTHuMnB793hKhOn93wKUSxmZ7qYOPvTPZLN1Ffx
6AA8fiMP+nXdkg8X1haHaf5ltNRJHHeZf6YUBKmMy1He36vjVxQTvEAe7pv9jgXHSE+JvIuvKwcZ
7LMLLZRRN3iVIcsbjHwfJ1iqj3TfxRe+FqDwb1dn5XBU7ayS8t/zaMBbsZhFH2EUUe7y/G+jQSgn
lzINvK1/IFkokVdhjabntK7zfMZ+CpMVuivrMmzd2Wx0SMRz+T21RvKz7dgtcY5sFDGq58RWhX1X
gIkcWHOks2U0YvTuOqpiOKhtyxGU5z8B43ZdpCWzbe3neBln++3A+LkhB7CCQ/v5nklh5XCfkWAP
VBki3IAjS3QcWkQpuDh/CSWuFJ9CIN/JKfro130q5YZFpxhEaF7RNOgGy+P0Z/KwLFhKGqGRfRle
dbncl1BauP7PMRkKep8YwJL5m7gllCVlg42YxfU0Iulalz7FLMaZr3dwXhlEkrEo6wfy+XhQvRok
xJZIGUhrgeyZCo3Trry3B0wBL+3ELJLI2Ixk5SYAt0jZqXPA1KNL38t+D3/5ctqVTswn2Ph1dULj
qlYKx37J0Pea0lBerL4iSo9Df/3yVrUTmdnzlF28LhFJWqbnEBWGhGHs2wTRg9t9SacX9JPBnGUE
x47h9i+1BOQNfNyHaG33EEpAp+0F0QRK1adcVo8YL0kkyKpQ/9/llwJpEBbxPsSluFM8vsOomb5K
WX4uZ4cCCku/eXjnl1vhEthC/zLUi7iIOcCPkjgwKcq4nGasoMBlIAcugYvnQV7+gZyJZuLMXe+B
FEE/GuqTKgFfTo0bdW8Bn5nKcv7jIvLgazMISir4IL6LPswzdmWB3Fk33OQkg+DN5B340ZNyirkY
HzoZNw8woE46DHhGQEU0SCB23veK9nUPDSU9jCuotp4ttMkmcbSU/tTwBNeYyn35+ASi8aES8Q6Q
mv5bpEbj9jDWYYrS4behXeAfoVKCt+wY5XU+NDt6j+IgM+J7LA+NLi7PciJWOnyxB33crzBUGdMa
vglhR30o4aJ/QdoDmCIrEkdBIE1T1LNtg3f443Vrvsi3aS2KZk1wsjXPrYNBXvAc2s5wXwawP+Ym
CbM3bam4JI9KDc7fSlCfnlJvTCokzhgNryP9z2WEwZBFSijOwdxjxWX125LemgElOAD6hMKwefPR
x023H4N/lnRLU6LTOMfdNB04DaDWA9ulQ4kgzCQrWMwwqeqODOYqVPWu0XEuSVYXgIfAxUd968SS
fblrDTdFbBfJ/HCTiM5G5+r9yKOqG68ittbxNGmx8G/4G3GQNyGt3CMN+vLC6+Ugleyi17kguiuF
7Ye2J18Qm3dLjJopE4XHUqBPq3XT6Ia5TndUw+9RpebbIYZFGofKbFoQwQb4E2fHKbUIH/jmONoa
cEVR+d5J7Vy874skL15nZbj32iv6T06ZEFuQTSS8NPc+XiraA5GlsO8ybLMlTBZcXlFfRwH+tZqi
H5IlwMiYs848UW7vM67hir64xaY3ezZ30j/8dWZA7QmS+zCQU2fBywiarYTy1+1tsz6L4Vmbrc4X
hJAiWgQUzUOS4vp4gsGqX79LPB93N/9tqvgu5hwMpO90TOfYTi7/qUrbn2AwhqO82qHWZ6zvlqOU
PyFWnQXv7NgtFrL+DmhmzJ6EJNaAAqFubA9dcmdU261DiEEdfXggFtO/+PcrpOFVMj0EnTTLUcOA
lSqHkavaDx5uFLfDtiBFjH4it9Cm4Xm3dYZKRi83nrKLSea8+aoA4xXtYE4sYLODPrDk1eKTK8C9
pd+4PnjikpGi+qsSVAtlT4N4Db09yVRJbg3/b8fkboBUxgbQhlAjrB4yHw9Tn0rikqW/tKPQJnyP
G8x9ZH0QXU+5xl3dzC1eXWVkYdx4KlYvX328qNRgrNLHbvdiYkPmoWTMpRh/+ntdVHikIAm6ilVt
T512c5vt6vyNYKwPeKnGDAea5cCPoY1I91fHyWdho9g2Rf6hCyyTxC3wGn5t/XDcz85jlDzoqiHK
ua66ahPGmM0ZSWYscB9RxcNVv9/YKRLJ4lbY1dvuptAXoDFOgWv9NIgV8JScfxhXj2zukluA/dmv
jFnz2FtBHTWiso2oeF0en0f93OyaPurUjXXeIVUqfpDQObYP12ZEno9OMM0NJu66ciJdk+wxUwM8
cRwYmUBpdW8r+QZKntbodXH9zA2z4LCyQbAYcZET3lIZno+1G0JnK/shca6MPtb4BpCZ1ueCUqWZ
P+/7kFYNS49DsadyY4brMvtHo0tMJb5JMjhnwtY5rbiQmFEn4DmrWrvzQMuT/vfjGHkYhSGCZ26I
Hrkkwt/odcsiQb/IPDsv+nATzm4BEAEvgFQwyCqI1FG/7RBL5C9aGDI1TMr4g0MLv8hSMlgb1XD9
G4q4aIHqlRUJ7KywW6D4Jmqbi3sKP1Gg6kKMrou7c9JpVUNz/XGK1MEKRUwMjwvDJkBAuR6QGG/e
gutzOKlaEYMZiiUmIvdMb+VletwwsCU1ECgV549C97FkROLezcu0lgZexmYDSYrTaRNmWaf5AM2r
YVcmt+qI0R668WaUIQ2y60PIGhZZIc9QpPLjycNbHclmmwk15/7Uap7I2wsLp6qjT/faAx6jkbjG
hF8J+OhsjlD8nOGLVd+HaTgpk292oNwUYU33uq3/shyjM6832tZmWwRRA8AiOnSmZbMxFCahplpg
dictLwNOlJOrc7dpPTlidpa9zOjWdUhMYMY0ouRU6Nf4wP61PKz9JZr65i13gD2y5c92xgtD3afT
Y68GpfYnYTHDDdEYHmiXN3zHGTC7Wo+Ko7nF6Ec0FoSyIZDH9iCDrUT8NFb6rdQnzy01QTrRGjxI
U5hK0pr3x+zbjc+eociWqDADJOxDlLvv3uVUORB1IxsThPylec+2JKYyzM5KpAAQTF4pq2dbA9NY
RxypRkkp5KJSBTr+ubz0h1ywyuuX+dFcTH4tFAaSwip62s2+NDXZb9LVmPBQRoxT85OIY2BJVFaH
zKQt46ABwcOcEBWbyIB3GmM5edg8FYP9yU6VFAHBeQXASMIppU1NF6A1606P8BSv7FLxi15OTzIo
+cUmrOcf0/62lIxo6cUNosnFUttMESRbGXbGvFBySXhKpcBtYpeF/a64iaCpsf5mmRxqs2XADMO+
Wc3X58BEDBTVw/3UWzN4/fJqKDaSiHMK1qDY2JpkYdQGWM47fqFqU0FlT2gWfDhx6LuENIm+5MB5
OuAP6Lyb9IZk0wc5V497Yw1EKAm180FaYV2lDrr5gAmiWbRKX7IWvqtyPtzFBmbKrA2+f/lc4yel
n+oge4fllRN4C05kEaKxD1sKpqxxf4lMJNIfHuN/yqZKHRF03erQ+diCRIUtbecRp2G+AIWGKQhH
kWFQf5+asCu6z/7zyy2i8Pcmxj4aX3xDpytaUbQzjk+kY6gak83M7bPIdQCCf4ienhkydvH6C9U4
HsX7s6ewuQsD+ZNwMYF8Nnzc5v5/w63WQzz4x68ZCBf2QJp16QrwZpTlEQL/HUkNh68tKdoYLxOn
iBCC6YfS4VobQokCPrZANWcPcW1VZfnfR/6gtkRvgLves/MPhBNFm36q67g3Z6G8B4fs005ewxZh
2bQX9izxv/fMx/O/odqb/RIC8SpZ5IvFEsTE0EYvjaqa/Y54R9BBBK7vAemxzEh4pCGDVbqEucDk
x330TDaj4G/9e5vZR5kkW4m0bYpfrGKVdeU24bspeURL6LghKRlnOzFoTljt9rBdBuL/eY02lHqh
B+gvwyNGgDJvsNwsQrSvxHyR8MB8JSUP/Kv1hb3N9GCp8pcH69K3A1mflehO3SK+2Ot7kKj3mOLt
YZQynsUBJLdIhymtfE3Z9W2/vA/0Zx17s58EJsjJ5YuFFnv8PiYKBZK5xFNpF7il1gFzpwRxI8a1
y7ct8VrMCYIqSOf2VrnlrnyLpbmNzaowfsbd6qLWTNgsUWZz96tmcp05hrjCOGpmLV+XlgC4lip4
ggUFx19NVwMIIKxZ/71AtbhbvC6ApVOVobxTqNhcIDsj2Xno/b860FDf9Duh2jQM1IW/fNYT3wpR
AAyKmhqHeItxyph1VSLHGZx4omwfyVso9KURylT91M9lCCbOCFAk8/gc7yYWtT0O1n0HflxPO8Lp
bJ7XctLObWQakBr8iacWGbxf440eI2TgiVYg1Whm7CEMAX8p5nvRGKfDtiSQGbgZmz/1EeKztln8
oH9ZJbqUkbhjsjoDtFSQdc5NeD8zttb7X6h44+T7m39GCjq9rlqnVZuW7csIZff/kGV9JiF2bM3B
tfA2e7P+e5/FiwYZ/xfKZHjxn3KQvknOuiqMVTtgQHUqXy3wo8mDh/HfxXbXKDQih0V9xMMQw+Bl
gbgFcg5QFUEE4E9azu7cZndCrWGIQ/w2DbYVJ2/oMSbFjZYv3de/9brG7EOx1cXPD70R0ZiGRnH2
B5brQGImkNx34djRR2vr0NtS2RzfmKFiglQb1mQg1IojllNlNP8MBPtGllMNDiuf2veWW8/Ev1lC
5gl8WIYroHPUb2bZ8jq0SqLIo/ULpL4FAkyHvreUaF/SNZ0ulrAGEJNwhpO4bhXL6YB56NJ5U0G2
wHTDNPnUa4gfunBYmndq1A35c/cjNObEXMXJWpksoerWVVKPsZymhMlx0ovUtOtqOmX5LOfQIFDZ
6C50Lk+kwQaF8UAH8s/Ymi1Tv3WewntTy9QdZRHZNtODQOBhfJDpyAs/8nCQll50WMiz6DdFXtpO
OaNEC7oziLBQCkDqbrts5Bqu1f0cBNXAT78ckZwT5PIFa0EB/8DV6N3/RNjQqD3pDQauey5NNSGI
qD/SEfmoOZWKG1GNgwd8XrUPsyuD+2jop74JTkSsyhM/EeECEb1FXuBtXARrGA234VA5dPOTU60D
rJjVoIYUML3d0pKUWtFzhjBqvc4nM0fbXk7QTVqA+P0k2V0JVXjRrcGqjSdWzUkYZLe9BKppnzKy
UnrCaU7hQGdcey7BRAyPTjJz0N9Cxg5K2/etW9X+Ai6ZQt0xMc1DNqVIgqYYD0iZknZI84fnD+Ki
dFa/01AtWKK/ZtatPTGXjGvE+oaampCFLnXzKrL7hr7L1HVTE1eDap7B72VxFX/TBxMIFzFo7pEi
a/5HtOK0a6o1pi3CaQOD8IrgApA7C9kdqG/n99Kj3ohbKjLjBY4UxzqrtRwXtCTp/3jqRLJ0KxcA
8RlhPGPyhFP3AwFVDaupGdu+M4qm4yGLbm4rvjywsh2dzWjHP++i05ZHrTk4w4xDAP/tBpkJFwJ7
y0nQT3QApbOtr4KUuiFaJpIpawRLjft2Z3b2bfT50TGklXMESq7mwUsjpH/+GVMqcNo+F+pb6H7X
9awPqYDph9q5ONhd8mrBmsXb7hcHBvsasBilNndLs7hNMJkiC+IEmy3L2Bu+mhnwtfxqfKyiLzhF
hHfjxM+39KuZpNJuhjanoVMQ+oybSaGoLJmOtGVD/dDaN1PKEiT635L0G5ciniQhcu47Clq4yGj7
N+qK5SK8Z8J5U4OIZc4vt5Bzrgw/XwviY7haKgsOavS0MBvHQ5uIl5nMs8I7AT2vvnIWlt2N3HJo
EfLrwa1p+9n5x2OLfugb93rSaHE/rjwjJJxAFksgQVfP+mYUy+LuA+MW6NS9kUbHIiBWeYPu0/Ce
yuucsRNO9tPAg30NHtn1exLTMjFBPsmhYzNahw+nHX3sYs7uKDsTnQXWhZ9AzzPQnXVha2EEeNhO
fDVIjxalZNTDdaATvUROcwFQmVIxIMkh5U5b3whZIdu/216zZqwZ8goYUo+dc9kUHC6InK3l7xmt
nEyBfZSypzEzsfLR93Py0Qs5ArinN06rAjhUlihc7zGT6Zy4n1XIiNZnHKkbn/rCRCzhTPYW21V0
TSVJ5T7lBk4F2MuwbIj99aHdd57GQFubOc5FblF2mngyZrv2zFNo69zSFBcNnBP43RbF/T54fFsT
hWjvYYEIxBbnTXdf8anjRPJwskiGczDV3cTZsT3yCwrTw0T7Oqp9KHwYws367lxWeGhafaxh1B5y
K2KY2zORPZp2gHUtz15yXsUzcb3/rc1a1PJuQPXLiuKJ8HlRYqZe5bCwL+nrzSZljMDn0y9s4oFi
qkTABYfxMFY49d/AvTS84ZeO5rJSoH6CLYzK86PnwAehdzUE+av17hrymGRgFvVR5CxvEIfTUwql
+9g46SDilmzFsL6RR1WkRU4A3ff700xLABqUcaP/X3DPeaqmRLCgP5oDHsG9UiUgowBAUgy9Wpjj
S1B7tUXkVyyusjtNiemwSOSa74In+3rNcYeBevs9ZfXhXkXoZJU1NpcrSWDt/dGM7HL5oX7OXZTI
pOZv2htbuRDnhgiOgGarITHqe1h4evK+cw4O2zQD0XL73Mg+MVFogdz8ouUoX0ODJ+lZnOMn9S4+
bspz/4wTgXp0DPfMTGiHpQi2WWZ18WrPAe8n1q4Er4JE7Dbg0ThDlaKJ+rNNbke0tdo69N5PV0VC
4AR4/lqVB6utAXBMEnDOLysxBb9Iv9EjB0XOsWAcqh+bqPMJzPaB8XpoMeX0XH+cDduZmdOTPuVr
zdTF59WYP/2C09sQFiJ71+V30CvL1aT5hC2Uq0R2zn4DJ6rcP7AFpL23wAakfOOs0RcVFStaDm6B
weq3yt7HcJHSvPB3AZ/eelCm9l5eyuaEZoeqsHcaN/5AmoAxcAem4Vj2hMz3SpilhTUlZmGUdJVm
sWhpVWHNRalnIXKy2QoASYrGvZ92Gw0gz8H5I9rUBjR0djR+ticx9CGzwH7ooahVwi+6eulW6h6S
fVPow45AB+6xFKUlRNT8P6X95iKNCHgyaT9vhRh0oBjwfmGzlIdQilqnGiwUt88gM3G5xwJMTY5Z
/zBVtSjnr+XXmRMAwPJQ8eCDRQvd5CWTquw2irDedEURvqrDmXaF5AjRR/NB301Ie6KuGZwVkplj
gcz23QqGJz1YpqlembSVEmv/I0kgt9bSAdVEcXEeoUihsmCEpQoin7x/jn9UB7aBwlj++CSNj+Bm
rTmIjmcq7E5G6p7gVrOgaLJkU2ZmMjb6q1nPMSf9n4HLIBGWCMgTmcduib1VotHNfW0elFZYOsRZ
PilYJClXZDtlHssI1CYqE72l6cQqEp7tXRVPNVoqJd9dQqh5O+DCV2hdbIg6vu4CEKJ7hFtpjxzO
WYwVdab+CJTdIaiFPIr0pEQlfF4mVVL0O1Dm/MgHPHTNWDWAuHzfrNmIkkXX5z4j0qXXhTYkShh+
lPxAMCFX2akPpoqKTECYWjLHy+dqBCbVZ/t+qH6GIYkm1EJfQkNgbQETxPEcJs6x/8sViLWRjArI
vqi0T1cTssMZOWYLYfi2XNvMOUxcjluXS1a9VtNGdwj8e0W9ee8oe4bGyPg/yLNxBsFvzpJuqVcU
ecfAe0fWyQFkcOgSnxo5vmetTuXk/F5WeJk6lvqu+JbRR5ZX/yjgnf7IfzVIsLSFmZdGED0hzA1I
u4+YjJvgr8PJkG6SzddvbTpvCYozLjnnnpclkAVKohRW4J0p5pyXSNBx6T4+07H4Y5EfJ79XW1Aq
Nu/872FkoBor1Dun1+xT4BOEoscYTAxqTG4hB39KMpCOscijZ3l8KQbNLLZL1ffMKqOi6WxLSTaS
zH+opTsmHYUdHdpX7wm6O3084ZUExVCkPTW63UmTvR6Ql3gyzleD+izE78tkUrVuFQ5rduXGN0Ed
lMu3gdOrYcb/ts3gn070XpEiLzi3Camh76eEebtFjWpnBBg7hjI13KWlVYDsjxQtSjFrVVO0Y0qC
nZc2Ixsj2V/pU8BLClzkeuIDTF7fwZ+Vr/oYua/SMWXaqiwR/FQIdmY6qfaH/ytXBXlmrRrDMHzn
VuLaB3AiIxjbLdbVq38zpi+aRR05bOymS8LRvHNJo6F9l4ie1v0E70gpnpuOE44K8plutPtF9xnH
fnKVGeSDVWViXk8L9a4eUUx+DBrBlPdjuLC8SKHW/dPUh5XSuMk5L52UFS0wtXIDyideNRpEiqmW
e9myHHUKCFCUhcP3KKNRqt4TrfQesgpPRM3TDONkxC19h3nt3tS+68a3A2iN5GMJkJWe4zOuEkh+
sBJfEB4q4jt5RVFbAUsLTP1QmHstHYU5fuveg+G4PxEkMB7/2qqq01ahZ3EFcpIjBrP6etEKXiv8
nvlThnN2lT/y1elN/S2WWWhZJfzrd+mCjpMQBhN67pNT82aCI9XxHrfN6ewLSn1ODDhbS36kB9UB
uj6kyiBCP7fc0q1LQdRDaBF5VQJP0VPKrSaEh/brZrHurNWmeg8k+02AL8o7e9xLRh3RFUUGT/Pf
PBqQFU8Y0UzPZ1w36d9zag/atamxZR1iHmjO8vdnBVF/Meee514WD9pWql7Muz2WvQFtBOno7FKk
gf3FLsGaywv530NeKGFOH5ku+po+8T9MxGH73GGwl3ya3qSxdQoOh/3YJni+FpnzAIE9bocC/jSO
NIUKr3BpyGGIoNQD0pt4mqr+8dVUH5wIhJvOMiqCe2YLjfZ4mhiTZP/L4rfTNi9OleAk2eUUPVrQ
s084ZQWL6W23zOxNpLVeByRGh2nAxFGE77+OwT3BSk9GtdB3PwhEHziCaOorIpvQMf7MLTF54xYE
RsuHYWziH/o1/H+deV6nPFvkWMyggRBkEXc24EliBYXNUmAdCblLTU52mTHeqG/Hig/TrVQXezt/
rrJPTXpWuwXFWmWmV7+QbKA2ZwWZbl2ecP19tlMzqxdsJHfW+OxFYRUk9+Ivqjeh6GM+ZRqLfWGw
YB5CEofDRve+pIxkgT/xlAIv5xhscxzEn6GHC+3PtKE90zA8Jf1k3VeT6kLMshiydWZGrZ++rsDB
WtXixvutCLbg4qb376xDbA/pkCwZkIEGgkFGH72B3/xE0Iamve4ZkUeL7hV2p9qyE3qZVJ0GAxHo
8z7TQ+LCFK71o5DdTOiV6nXeJ2PqGk9bosFnjmOuoUCWHT3xR7Zub69DADdLgpAsy9/gxs4p+8sC
h6x11fuj6faJgkyeQJWmz6oGYvvn1nQVa0siJ22j2xB52jd+DrKXyV6GkroUghHB5bP9i6LeqNtm
n3YFF2F1BL7XQrJnghNN0M0dPzBMf9bGHE1S5NSUQzaraka6MlbmgnWPPiFlaUZxSseQHBnrcJ4v
MlkTQVubgo7kWJDNgTH0gZjUS8AVQxVOO0fFQpsD9zWDWiparDifoZqBrC3UT2vJ4cmAApCL4aBU
WOFH/U3t4DUS1NcgSG2zOS/NB7ZtCFl72QJdg0dU9JAeRCWR/AYjRLFSv9+sVHLYjPUdUUNgAGrq
zAQw+/Ky32Ca57Hsbhk1FjYwGyA4Mxc1TpBUMT2gP7lPjMM+R8rk9YkH9NJYur2QF/G/emMt9a6k
voY9W6hb6mFW5mLcItcbpfNE59m0zHJJQ0fnYENV4D8og5Iy9ZpTuWJWuIOVnbuQshlDhujpuyBl
hKsl+ItKM1mkOax5NTcy9KUqkR6rN2pqcFfOQtFk76wc8IX+ABahRj78y4XW/8PuCq83YCYJjk2c
bKtDsL4PNgPWRIpCF9rsGQFLIqkB7f2BaCR4mhMx48ovSpTgJERttsTKmpxdKwkOUO1/QvbuPpXl
22qRCtx3OCdxJ4yrK2GfSDhdlddB+nS42hPtJpK83HYcklSh112L+4UP5Tz225BIW8dSHiJBjD/j
sMj4U57dmJ4rnIMktLogT8TyU4XEOAob1YDP0hD8lfGFDLOnbxazFCSRdisfwVdwxbNraVNfeQio
zQ5QAaqBmHWhkKIQ2HybrX/J0iGggxJN4gzH4uo2pMSmkEGqFLCf8CY5nmZ/j8D9fVIIAPK7OqOZ
s/7ollrpsRx5Dc86wv+bg9oaTgy+H/XaCuhqeDvBcHxbRwqC+sZYzkVLqA/Z6Zn/fs0Yz++NowoZ
0J/6p3BVmGuUASFB87TD2zlSlhiomlpG4479CYD3eK6ZJj4tu9OV22DW7oai5g5Iz8VXbuupL8BV
se4lj8VKPAb9KhdflVrFY7Fe4jgF/3YndfCF6wSlFUM9InAPP3tmBLNHgernoHHuMPUg3RJS3wQn
WaD4onS+0rcS3GECfmUmaPuRwIUBeDHVbyZpQjeat8NDfPiLD+YLNDi7tnynRuJLlol/yIt/mUjO
UniN5T7UWIZ+QYN6oz+ozWElSawmandjWMBTSPTUsiz193YK/pmq3ku0DXkdlAZ3iP0uDFGm9ETO
vF04ex8R7p2FRJ8dGJrYwjQs0l+fEJC6CNcK2DJsZUuTmJzz6C3qRze0VE04prLH/GQnaZRXWein
v9STVzHqvhOca/BBdSC+qK0YZYiae1+q1vnDCVZryZu5zVjHZDN9gW27SNlQYopd1QFYDUxffX8Z
tvn1HBhRf5ga+OwTwF+OmQsRjTP7Ljw0b1AvZh8cJzfIyCWlc4WFgvni3Sn9cRNa1GzmOgFnagBb
WscUxyHysTNGHp7TR/P2vtv7QoIdNcOSfWhgqWAH1UV+CWzxHtGOPTwdib78TEu3D/yC2TIbj1Tw
YV9p0GEKWxYAnhBLEqmeye4VNCL4J5w8xJKg5pTe4yFYKMNgBYSjpUJ3tsdbelTSvtwtdYDReJva
vVQyMnnDq/HcEENLdrmv/mC1RE6VgItc/W0iXo4aIOoArrPT2G4qCwFzK6wQZVZZcSLnsv9LNFYR
2lFC3GWaXvGHXfz9fqpyNnngrapmigTl4nStUGD0el70vebotkGW3h1V5VbR84BU3Wf9aRsUUo9f
7eQQHDA8/eFB9YlzxFpEQYQD0roYlcTEmH6LB4cOnSr9B7Ju0DQVMqBBu41SQwzlVXRbqnGzCC4b
wP8JzCbZTo4+fCrK6ODVhHmXbc9bdQsSjOA/cMTkITL1/KW95/7iPinyzNTU291LqOgXa/WC2H+r
FfPvMJes9dslLHqtFZ6YH/BJHYO3LEOX+g5q+ZfRKYoW2+zn0ovNILhdw/6rKv++PcWPfXUjb8K5
5cKxZudMDjHVRrgi2haEW+2KVz3kqylx+0cjwvAknl8UjIfeokxyTOCtvYQEeS3pajCdHKDLaLls
xMLBhe8pdk6RsmYtB45Vo7SZFt7PeIFPravNHZ/XQhBxWSJ/JROtN0iiJvv34nPWX9JjpugoCW+6
rk23aREGVv9C+LhZKEbO4YoJUmITAlWECAMgD5DtUcTwFOkO7Uqhb9akbWHjY05moGUY00gCXZny
5w0mTJSpeptsIWhotlXo0v+hqVZq4MXlk6Y0vm8LJyKXOFXotf1vVECIPSSVVAeKx84FknQ8l9iW
diYONL5xSgxeIRv64xiIhQnHnBKYm8Tz9flCFSpy8MhFBMhBG6AItgW9Pe663Fn4mv2CK1wM81QR
2CDyJ4gccDewFjUVfsVI4kvrEyqNq6iYIq4o05ypmNBpnp7cgqUG0gDrWeXCLHt9VWtF3xl/l4fs
BLpscca7nuw5FrWIujmFdVlgxK7ux/I8QMqQ329Scx2Z/A0Mim+MR9pyktufK8LLibzrl0MRhhZ1
1uSijPtL/l6SIoC8kGtbnWHJ4cTFkEfM8CTsmZhrzcKUVi6tImxcrSSPReoWRvgz+LkOmxNecxnw
HSsShcsV2y06GNicBD6bV59psGKZZXPVrseUZIkmhnY/Oe6lk2luEiXOzY2YEiREDKRiXKsdl2Xo
PFPeEQDXwIS52vagcvRtettKU9FLZnjn0ywz48uyGKjBHnppkXLANrb7xnpRwGsyq5nTWnS2PX4v
YvXUlsQ2T34VzZ9KvNFO9ZlOF4UPJ81uygA2az/uhKmwCOqtPyNNXfhRcKKK2Wi7SXrlhaC/I6os
fgLqbKhlx0kwjprfRDxNgOvwcFM51E6EsdRkG7dTUFFz6o8PLanZbUvHii00GxRU7DmgRGviARHP
CVDQdE7NyJEB6Auj5zQIkWyDBbHDvBcIx9ygmSadLMizXxgci91Fticzx2BasbLOtDPArl5NQ8+T
bhZ6qjts1q+EIp8NonkewgeYCxGwyCFMiZFZ+i2rPdbY5+HWs3qK36f/BTYoDeAJr1ehfUK2+Xqr
KwuvzTaOtRdG29Kj82QPZ9sTpod0mjgSeZ7A/wqZL8KxLN8lXIj4R7kOJDOpzd7p2wpuGPAPYrg3
IUMGt8Qpbih4FusU9DyiDI1yFNuLzBKowxW2WQjmUxdjUYBfj3OKR3n99V9DPuwq5yicv4GMyiJz
Y/Per/FVALDwL81QItaoriYnqPxwCik4Rj3egHQ7jBOfuqMxqkF2+0cZAnTlPmGhTZsvj74vBGVD
BKy3njaOEQ5rjRWW1fzYTG0CH+2R1jw02PhDCBLYKIiKc7tIVwJ+Z3zPn9AvNPrLFffTl6YUZLFA
uyHs2iowBjO2712tdXMI991YMI+DMef0FRCKslX6U2a++bnv+n2BvWBYhckkBin0n+4KeNw2Fz1R
YXNbpfrPfH6rVxbnpuAkkudjZKg7gy9xdOGowCYVTjpA8kflP8++uL/VIAXchUSNnvdIjVJS0Xu5
xoO21Ti7Woesb1/eScNtbLUVchNnlBBsm7aLJKwMXpp+QQlP9Vy5ZLxcffjQhnPwwAAoPjQY/3Jo
dyRpSCZCi/xBkbv87y3Ozn1WmBpQNWxfVDNjD5bodzS/BbzRsYEkKyq77G8z2/Y1dob/gUCdswPm
YcGox7fykMebPEkZky0SwWNKiGWuf7WSH353kAr0eNqLMPCd2B4cjm86OSwGF99xk+WnyfkVVNYE
/VQ1KLo+P6Phj+wMdLfF27Xy/aPcyjtzVgBbUeJVDn0Wv2d6MVcC8+257TFfjaZtKRMeD8ezVo+y
oUopEbSKw59ebP/OOS/IAY5UDKp0nQeyEEFDEtdavMIqhNSsPZ8G9x6RdiuYTP6TLQj9D8k35o7h
FH12xOVN5qp1by+Zhze0kbvCP+6Qx2v9PMldIEBFno9rCbLIiW9QyDQ694fKw527MZFDEGx0ueMO
nlsfL2zFTAuoRtUu3v6FhOkbzJJnnaIlQHbxhc37Ch5Rv4YAZxhij2YElBX61f7iERcs7ddC38lw
aP1BfTzy4C4L3JDTN0UzjG3Z6uybxxQptoSWM3QtKpdZnB3lTSTJy7rif3n/mnPKQUreBwT5I5eq
Vm8QLPiIe2PUjw7Prd3+jYc+A6mxiZwRFXSD3qobKPsXdxcWWx+qHtZRXK6BddK1WOcLQ90swfE8
nDS8N2/noT1VWG8qapJYLQmRkZh3DEXcu6Sq7GZsdOwoOUuk+dFJvh03LX7fCknX9VvIOroSlm6h
mezzPL8VrANfy/sqYvSIWh4o/WGoAfXNAR3KZ3oJmRpKx9lhiMr49RDWXMejB0H5bvjQYEl/4G0H
Yf2u8oeQja1xvo06+Cp4B3fOsxS2xDIUhEQG9UcXfZ/TowAPPEFrK6NUrPGNDKo514Vzq9d+Tnna
zAvf4h58ltWYh4OFN7XyY69aGfG5odr4vTS9limsAMVyFKxw4E4hFt9sgKFFm5TCVd1PUWgC0S6Q
hCzlaMA4yil1DRlDzoZJtgpdov/zXBO1tyOyVL3VibLcJeY6BNtL1IyZ1BVgw/4KApNYSAiT3KGI
w5jRU+EwUET9czKZgkyTFG9C9ZJofAmm0Y1xael8QoPiF2J9ykOIvGREJVuWck7LJ3090TlSixqq
UYHZtJbulVsq3dW7kAT5H/7N9a+o1S3c2PkzuX7t8LTRirg6kk+gN3l2Epu0zVLFyjCHjvGnbf8K
AoyFEgdvNigs0QauPNSjOtn8xds9LFPjw7v/Y/IBnENGQP6ab1X+9YTsZoQWWyB+VhX3DEGCzqyK
mQjYt8VmWVh8gYjtBIUeWGKt8cfnGHD8huPCNtFyVkAIlO6Jx9Fq38vHP33jBtcmAAo06a5c5Cms
jBgtfLtVhR895NMXs8mXt4h/QN/KJ/ywvCkCuM7I4jLceXdD7JJrUAGQ2bii1FSNzlA+OIn94zPj
2iY43wMcrk89NWPuPHor7Z6rHqK+4vAgBwOFk93oFpz7AERXYHG99IrescQvrO21WAM4IIlhkdjw
IGQuuILWUkAKqq1dKk/Ow0ikm4oXQLtbCKILinOU/kHhZkB1ERr//H0X8Yik8+4LAEQv0N2v4r8k
KOebyZqYxsuX3VC6fkBbPlO+ynnoXdxLfs+jU+dMpiseCKVmi8Ni64ocPW0KATACHs0Q2TYi6z73
OS0DSxzu9OB2L7HyptLZ4sYxy4LKRG34F7Frt0o7icUPnNvmQehn1zHve6dT+m7vYDNj6xCMqyjl
w50LN0z1eEsFa0rlZv6uY8cwWyhd7NfFPOQyTM4RMNmPR4Y184/s2mxCWjuI5StiLaNTP8EucPcV
iiterOrP2NwnyrS1zZBF8jwGmi3dEQWAfyYg06AbcyWxgFKzImDCCHu5S0O4DZfKHWHStHn5BnNE
DaUiKo+dWRQrnP06mEVbAnjWzhMXloo6e51cptfFCD13YQjD4TgQa9YYwXSuEo8Eyff8G/gFulC7
rahCrrkIGEFCIUkTEmnEiOnN0f42mfVBlnvtdNpCxFcTJn0080rSJKtJwysxBILRXuiTpTV8ty5H
+7u0302DN2DttAlSRu6GdkOcfbFIMPUgZgn1J09h/XBrHjbMmuC5b3dM/XWlQjNkjWVrmhQV6zjv
lNFL/1hg+QpJAVdqJJiGiTzbZCOdugfq8hoiLjMe1o5V8jkghqeoxc+qcpVNPIooaOAiUHyoA46P
OyeuiQ/Jo+/I0EzIGnL7dmKUzT6EALTIpE5If7SfhrDRQzvxKf1t9CPRUzbvIXnHUaPJXrMTGY+p
vfGve8/oJAj4LJGDiwJc3CaLPaszuyKvqfJK/kW/Ui7D3CyxfX+zQUYVmo5+wA8UVDXSSCJaHeYL
XgQFnRqIjhfkf/05dATnNwgW8VdYgJcKhma0b7DI1J8J5dhbl3pdGfrA/5a0Gi0LVYDonnb5VoG7
JhG4nI7wpx2mot7rpMG/33BnRxzR8hnaZgzoWom/yDmbsXj/nNcCD0s5PDGi1Vd/git2WfG0Go38
v+kEgFrTIp0XWcTCko461kvsfV4W8dK0FPZGv1adC5DMFVyLrNe2tUXtNmY7nBTdnJChcyn7ndmC
TA46dU31E8Rm1E1b+ARFUdiXsjlkX9w+4Xa5bNf+LkHX2IJzKMu6ceD5FPJxq6fsAj2OGpZjmV5i
mOZTQ4E79SKx4G9AKYOTgF96ErMJi49/tJ95jV+V2Xcbjje/QjoEw6BN3g/OUKmDPHG0DflfEcVs
raMRyFW0/84jLBe1yR+iRxVasQ9CKburTOSgs4gNFw3t4iW06Tjb4oa7QwTs4DOUjltXiMgXSA78
PEWJRMot2pe5yWIsJK+yttG+IhjRRz2Emj6/yCTw15wxqKIQ0/BxeVKfTParCxOQUmu6jA4qfgOh
kp/+dsoVcWD85N9Vaz5I/Agdi1+xb8poiCmP5reo9vNdA6ybK0aQqU3fOXLPa2U7lXUtG/19UKbj
bVFbzmj5BUIP3OL0s+6nz85njwr5TfsCeMNMMsohBgqJ1gxGW7KESxRq0mBEi5FyjOvcGuCmq9zE
sGhc4YWEHe3vwdXcGTMImsaXBqrKY3d+OLkD3ahpKbRJJVSugHGzeMq7CwMyApI6QNUk5k7z8afw
wlMQ32ZK81/l3gsWR2HHS95xLflYxB/uw0vK5mFReJ8e03S0+WcL7nh97BSOHoocok4rIbrstfal
NuIMp+Dp+DX75/1HN6jB7Ta6h15wR3HrTUatxvzxeAjfdgJ9vONkOqzeuhkBLG13D8M/1wiG3I+t
i443QE7Ll3Xv0IjnMVX0C7eBWWC2Zo39rNM4zjhvaQFISSnE99aqljzDDycXnxqw9uXLe/Ixa2X+
loeES3QjIVs1aZN/ftp9SpTssL1C9DFHP1WnFo1mAMxYEzEV09zk5fCxduOCdBFTnCyQKP5gG5bZ
E4T39Dycew7VVvq87LC+uz5UqiJt5WhozUTS+GXvLZC5k+Jm651nrUH6zH7vxvLdprbb6OJ80uET
OnbuKILu2lRyCU4lfZdzW5NwGNhuOKULKgn2rHPq1vtVMk0ZmR84+vteVXiWfZeljc917pVgaGsA
xmD8rSi7cFM+cRpwk/EStz/oorYBlWNzMj2fElHQSNkkwSosGlxY+ZuFAFL9TDIgsKi0S5Rlz5gZ
MJ8pzWOmfquOnWFqH0kRydt/jFrQfxoGPZaBHJ7ib383E5xjrDMyPiAXpqjlb36EOV7jlpyIBUSo
L/WQ3lQS805FjHROyUwd8MAgnKpqUg5uzZNSFZekfcPh0QITU911hEsSYsbl0fq04W3eAofgNMM6
Bi/VOdU1xx0q7sC9ZNFUtrOPPreVbxxUty28onrhJu5bANNq1OcJreqKPzs0ttnIteKvQvqadir1
BJAypKJHE1bxtwMvchHSL7ki8botHCFV4e35L9NEJawIvQf5uc54o7kjiYPLM5S3I6LIVFQvfqea
hbsqupPr11vYwoQ69hyGRt+BE0QEHLbo7agIMPGCsk5g+cQgDDoKlEsVbRKfo9aWDB+ay6VaqFIb
mbsiG4UIB3G+alIiwfCyZQAyQEh1Knf+TkcCPdSKn3b9ugGTVnjkswTy6q5aJTOdCkctKl+0Gsrz
NaLNeSJOQCJXpKpaw+DsfECG9Jqxf7tHFl1I/UwRjYntM8uhCM4KaHkXDdgmvpd/Fnq8YyYY4Mjx
kRpTCPUxnA2zuLsDZZ0EqGlc1nhz4lkxWVBNi0rbSK50pkEM4MDDdruomV6K9xNyCROyQPINnZPN
dKgbbtP9BAppD1P6eUMKO7NgP7CvLU1y/gtribjUsQIx5H4DyvePQhHWn+PYxHlppV9JRRt05x04
nEMyXDtBrrRlenEIQBcC7KvwkBsbdK0bvz8GDNw7TbAX4h3Qv6Uh85Zdb2JZNztBjOIKd2bcVDWB
6zbMIBTsjPCRjltW0rdHyI1l+APx1sb+3jhe9MdgknqJPLVPQ3oGEVhdN8Qd9r31IxTWp7qUyqUY
xquxFEajV+V1uditTLDN10SPmyYCqy8ha/0kstPAOU4kfikMz4tOFRuiV1zP4xlZEHJ5w6O4ACE6
EZyX4KtHOCh6inakhAXfv9JxHFRnDGEMdVpiF0qswa6+Z2DJip8jrjHqxKOp6b/wQE6QKUQIFJOw
9o/Pox059j1PDvWIVqEHwoLeO5DNpkITyhyRGxcGvv12pZdreYPnLAJN5MYZveuVnVpl5rt7woEF
7QjOX/ARGywqE067do4e803P7Mv2RBqZtwk8oka19fImDijKXyGqoqbkS1nUc5Qk3t0xsrfc4n6F
cbbaJrV3BhGIQywAvkKHwC43B7LouueiMloNREaLgE9XuvYwqIyYWSMz18NBiQ+hTyu1QR6gWdrL
k6yW3V6mJ08Nu+YsmNob6awy3dkc5VBBFXazwj3xmgbDsVOVAbQEuwohtyEHKFdCIG+lYy7mmN1o
22UWzYvTv1dPEbjm2fvYxKF15d59AMB5z/k9CFiR0586/huqGkYiu8kgUKfBT4mJclxE1l0Pu559
979kmu4R97OfWqcTlBHOoOraS7IKzr0zMkhdYqhMINtY4dQBpLoA5C+qUj0TdG6fsJQ/npSUOBcy
v1CAUWcZA0dj9C15UENGR5+VwVq6U7nPHTNq2sHcrlxAuLHY9ZpurP+VTb5dgLjR4L4w65M0qpNV
PPaEyQybbhxYPMbB6xxbljUQrOKmKKebqC1DWo2NF1N+43gzGcGBAGms83WkJE5J84at6cnCqS6S
HoGq6k/ggRgd2Y1hJLBz90tegE7yb2g2EDw5/18mQtnxsl0fOCMO1DFLYHgq0CIoCIG6oVS0Naku
z5GuEToc0MswkP2O8D7VkFaKK44SDQoXe+ePqYmQJDOwssRU5Ku5bCxZgZN3oqx7ardaY0K7d+DC
bGwEpILhser2+mAXmztX4/Ky/O0XOhPKKrz5QJYO2G2X2mXV8mK97eMprITF/Zo4ewpOkfCXCiLf
nZ8loF4DZf2iayJgSnifoC3ICWcY84bBUaOjW72uE/QPrAqaLpqaFuUxZ+83/b4miEy0qr0CvmKE
eFqLmPxnEhEvMGw90DATv03ICjvxa8QnvvJ+1XWwfhNKo0wFaO/nFXuT6aR7hx040VPBHNITZlMU
YnlTD6nkDLVcfs8FDLWFDgavVC+wbJ1+NwAcNZ8PPbxPTjEGaDq/ZKmn/rkMcJIUPMHGJn8kc8Py
c58tpJr8P2MyvWuuIXqST6+FIBMoVpTdOvSKJirM0TTWCTjWg6rWkUs2c2u31SgxWUMfnFT96tqw
6veT8vAxobele98ztHc3OCY49TQRadAu9CnWU2tc/+cJkn936yA1Lu+ZFl4LFd2+QZZfnk8EmV/f
RHQqMDMYZ0LlB+uJOLNbkQNOa6FXdvjPSjbC/s3AZP0j0rM5+xiDhbrBdue9hj2axSQsjeqZw8wV
G7+SdoFLfCJr43O2kYvutSUAKWfs8d5GfRVyG8QOj5jWbW3jBgialwtr3cAolPvs20+nNCWdYDwT
eEkETemihCzq1hGRTXPfMGl9Mo4kq1tGOEuKwnK36a67GSUjryCE0YJtUuMD249ptvnILKzzMUmr
/5KSWL8OKXVtxJIHAZyfinQBmdzcxd7kOLVtVakZe+Ptn4dhISJjU1RO/LsfcL5bjFgHTrVunKEz
HxPzY/zgZiYwJBB2VVRWJa4vPTczTqVOJCEnHdffL8HbPnvDEy6btJziJaZmGONiEyrHE0D0s24+
hFd/2Y53fGJoIWBTth5p0Mc5t9wJX0oXFrQnj9MTxY4HfCPUgLBYFAsGqK1tXGdevh4/sFBDahhL
9NGXtl2gEH6bSHoYdgFxpJxDyyJcug7PB6boGsO4Osa1Vs1PsO/2DYYolQquuSX42WKNm61iRfcB
Akw9HhgtFRVkgkRuUO9WbvH/GCl5J+ip0iAr3nJctgfeJo4r9AdB1t+QG9POHiR8qeI62919n8+C
V4FpQH/TXZult6Uj+6LapNFbY21mm1Psbm92ZcU1YS41L69gpriTgFGHUrJlITGfVn/MMea9/6LH
T5wn80Loxzd0yzshHd00YGt062ZeA9PIyKuhZo+z31gnG4uWYLPk/xgjF8ABelfmlu6aEx53SYPe
Dcek27L8A+o4JJx7B+G+Sf27uxWFmK7ujA7gBDrXgHQIv4eRRj/4b1nfYJriyEOZCQ1iOMA4tipc
yQhyUtBuMG5U4SAWeIwk+el+N9Yfa00SRzPbG5Ev0WUTALq87rM5wLNLsLW/KtB5FiauWw4i2UPZ
+u1qrmcNCxvPRM01dM3EYoLA6RGosGmfsvplJocMQR12p3ZsKI6936qedoe+eUFkvhiHscOBmOx8
F8E6tJWqPYI4I+DP+58EdEYnV5o97qHebXZTRblwx3YIpaUF1+W73+HQ9VEvq6nWGiwvblxUBZHJ
80GiFfkr51VmUsrYyhowWqjUzvaF7Xm15zfPRF/gj49jbQdLuvu12B3Udma9cbkW95ZI+A/XUyGy
bX7Xj1AgGGoOWeqaMlgecB9SMnuU3zw0TrwYudtg6ZkveWMByOvNvdxjeYdO7Z87d2QOrrEDJ8tv
sC2QOyCi3v41J+MtwER3hLy1O66YqVX9/zpUytaBR+CLDA4yyORDQxNJJOoCc9t3iltxQjIClZbq
pRz1FlanhE0ZAkrdfMoiY2tUsP8rM6YhPdPOG73EnNP8JBriAR2RgXWGY1oVAgfHBpwRZ2wyhGlk
BX81QumZ8xu1qa+grUOKIXWRMSZ/6o5xb9oNVTEkEY7KR5dsAHCpoodlUgMsjZkKpUXTjdzoaamT
E/JI6/EVYuung6pJpC6Bpc+gziX1YPb5wSC8HIw4HiVSiXJpmcpl59ci8DPptVTsM9K7IkXAUjJR
rQsf40wYCAl+3mJ2k7LgSYqPUxcGpmz3gC0P2uYuYNT3bjbI2IziaNTy+vrwaNg3OZXqkbqS2DVy
CJaol+meTz3n2CvYffrfVk/b9U/m5PsvzF8GVE8gTzLa9p0I6oOoj4D5U16z5VTPK14XSlMM0jL6
8jdSmnDek8Avxha6PP9Bp0N530VvMif88WvAnmcl839ViUBRYiaLpwGZEPqf43WTMX99E4fonbCE
w70nF1LLGxHtLvr96EfEU7emRWM5tNtA3RPg/wQZVB9Uwwjm96eGoLh+nJCb5su5al3qC6fZtk/o
mI0+z+9TMT+h7gyoVYc5NBoje1ZrtnY/Yvg4P4uDMbK73nIfHf3QGGvL27vjaBIPRmOR7e/EIjVZ
9sFzVqyKxJYPx9iIhIVkfJwGuNhTlDe1bQTy5yQU4mblj77oIkF9GRgDwys7AD2WtCoyaLHB7AKC
BLXzwVDhyCt8G1h3NuwJQNvJ+fYKKfqYyJ1ijbEUwyvgNPOzlLd06Xb7E4gPlxBEuZlNb6DTD+Ad
sE8okGfIrVA0KsZQV8B1jVzq7FcVhEXjmXceo1nTTVq5TIZAF3NnRX+t7L+PXvEAgCXmr3k1sgKC
VjsGagfgpOiY4cgpLjE4T0oKQ1KBRSZRT2x7D3eJUGYA3RmP1vtBnZfxhclra2XW/zpCz7Sidx19
m5XH3wO4Y4DIoZfrAmCMiG5PdvzcDhhYjEg6Jnht3pPRVKorsBRDk5y3oah+ecwK2hGw+e0ZcGpq
oGotEqxsLFnuPnVulk3hbIcdDJlVpQ1aHu21MgFGkWxl+rtkhA/zK2o69ee+ewSnM0yk+bOcSY++
2wzun8J9l7xeUD6HyDRUOgSExc4A8AR2g2l9lz9a1QLzAV4WUu/Gy6VtJReYqcXE0tUjqMA/Nj0z
ZSt/6yBNz3ESFvEH4HxpSVp5WGM2+Iw1vyo2wZw3rYiTGLL2ApCgEOJCOf4hYabzt88zupwMiocb
PhUu6sRJS1DpMj6ZTiCAv/zSxOG8yDLfLv1dJ14+f3R7tYq4wfuuu9z80ekFR4pXOu49Jtj8gg8p
ZQ5i8f2GoGie8XG1+d6BDs7pfbLG42d0+Ef0qx5JTkNKQ8VqYRqy9MKPvVsXlmUoG4FpRWAVZP/o
dY+DBuap6uDKoVu5Ii4OMCqehGQrSAo98cMZs4vvzgUPPeiCmoezGVMm0TWNXN74EYh5RpxYvRkc
5KY/42ZtC4Fzkim/X+5MWBg8H4iHRmtXaD8NQp99oCwpYZAdDnFWX2xKjZEdGzKHi8Ca2M9o56k0
v/Ej0R8sM6J3tOWgejhIJFeCBi4WJVMFiZgmIFHggvqeMGOzX7MyPPFQgmUTFo98PkpCAdROnXBJ
kRhnMx60nVdZFrcaNNPEilXO/e8zi03imD46SwBx7SdfYHBn+1tkPMSZEkWC8pQ6W0/54SReYvc3
BrWMMJUxUO/PdrNO2oai5Unuq1pohgtxm7dHrMH3u6mycqX6RkoKxtgzUDOXHPvasTL9TfGMtMR4
q0P2rGKAYPvuHaLMW7GplCCJ/bGKhbcYhqkAx0e0yKRNtOR4V2JB8NnuDOOXHXV32k0/3DKPT/3m
JbPeFpLIk5bd0uugtwWeWsYDUJC28BsNSd4rkC7wRwrpQEhloS6l+feyxtyQqnSIKkKYiFo7pdp3
CdeMH2YJ+yyPy9CyaolGCaBPh88u1tNQQv0VrNvSx7u2WKL7sbVdM1YwQt2xngxhKpcrVj4iBHf5
ZY0yIqwvOi6AtPuiHXsFfvbkQPo8ls0u1JhTx6Mqp1vsnUtVCwqX8EJLAFChMwPBY20a6lXzMGS2
EN22kmcMGm1H/vFZkxu8V9ssJyRO4p7+zFZSC6N8z1VcWmasY/ih24B+21Zw7G/m06SZNsyncLaj
7qYD1gMHGHSdxxIwI+jPDcfcerJiA6unq0orycbiOKIxJKba/WcFwxd0Ubi+iHAWk57dj4t7Ghdn
6A8Lagl2F4EL1Wi7Y7uxWmsd7BfDvM5zCuAVN2amb9NAXP4CA8LRUWzkF9XDL0Wg/fV+8Ky0xw8H
tULxUMCtxGjsuFWDrTSFe1cNJGVvi0jUpLdtk6F8PblvpqNRXOnTRC3Gv2mztf/cp0xHlIHrCw9D
CxU3VaT2+ePjyyR1SeZpOoAwMkVnZ9/6HXCeU7Me65RqAnJacRQIh4w56wnKGjeEKJhZwLqhKZvp
FXAMgDsANngsAZDCAl6VaD1FtJlSfpy1Hh9eDolu23TcOsmNx/0j1k8h7nZE8j1cumai7G5O85RY
7C1lDW4xJhYg58iXhA+YTvRygTFDFxpWB2gTmQDT27vZTPqKwNsd2w2zrPIN7Dp0Bpp/lI9r8zeX
+PGL5pMBhC7pnl3/cE9oyv0Qu7BRLT7tiulFcnMHzWFEpCW03F4oauGgUNJzImA+Y+1hiBO4Q7It
bdzRbzy/0ZXXfOf1TXKmZssOApY+X+uUIKdAf/wp6qqrnnCs61SKKjrUqVePln6pQzYVeltpazNx
SYQg6q/oFVX3ZdfgyCmtVIkWrwRsVuuk4xNOMmBpGb94qGpkgzwkTrTLf47MYz1WqLKuHDfhq5Mr
+RggBA02W5v0OC4W1R5d0z7TztBRDaxq9lSBn5m3lLhUoMG3OSxAVTdI/dPEtddAQblo2F9gexPg
rSexotReL7uO3jQGRal3T0nzYNgNo6C7TxcDYtErKJBSCp3l4y3c+5DtLGBgHQe6OBak9jGT8N+f
Zs/paVlh2tKrJPsF4KkgUxrun/D8f+SEKzy2v44CziObz7VXXjTPH1ajIQbBX4YyEwrOz3oKNHPm
+83U3Bo6YnsqchEJedQ8ZjXcfJXsQkydnzmHkjWkP35V2dBkbS8FX55XB58NTNRq5ZcS/ZApq/lv
8+itI5jUonA/6sEsVtNHfiqioR6XijFAt9odbhfMR8MTDnToIWu7ciQCNBNgjzzAeNATLmDfI4Qd
vmuuQQ2bnB0ZqRh2y0U0hA3tzfGr3aAcVXOh0iNWq9Me5zC8cunIyEqrevdFswXqJRFwf25w+y/T
4w1NhT631j4tC5GqX9I0D4xCtLZl2ExcMMk7Gfq9i7ReBLLWH18m8tfAWLWen3g4hoQ4ZCQaha1t
AdB+EOTcIOjHxXLA2O4cWfSYuAfv8XSM08vuypXgQtwnwksTO5Akj/aedHwu8bhDymomK6ryc99Q
7k7cJ6OoURo2P1m04y/mtFKp4VccmBxminGn4zAl66IK2EGq0DSHL4HGQbfr8kArOvvzp3vFpubO
dJ2onnvJjbqpXlOK0auF+lj1tvt3Ws8mr4YvcRtNYADeQA41kpaxvNK/P4eUji7+SOVQODMe5AZD
cx1xPLa5nShPVPHm80Oz3GT6wfRlZsyGzQq3SufPwxmZE5WuQV/24cWdilt5C58MjL5I1uGO8AaB
m4r/pYEUNxGgKoe3qspl1VUyVYrPSlTSGH9E2V9Xnhw4lVv23UN0EEISljtGjZ7pbEr2xw+LWj15
wtnCKoTi7Ep0ittdvYmWxGwsiNZsTYwPqtM0KFSwBlL7zuUUh+4GU+mJJmx4N3gQhY36wMjRFDp1
PBNTY00/dlJei335RbqQkVbeZuCbSNi2XngfTCn2RKvDT3EM8SPVG+Y3j3DclgMIdNopZkojr2/2
5c9EE8yinyEydPMjBhTmikp0oOnglaECS9kgWOkHq8tgdBiEQVTGsTY5QpKJ0IzkaTF1XX8ZIVI+
D78V8fEk1j6PBWrvVLKv5NKIC3LFM2B/JtzUzkNl3xdnHt//wKTZ6x6iRhpTMHDP6sZ8gmueLxnv
q+Nys0PfVNEMTK1UJ4FUx2YwV6pel43O8XajuKZMmgdAWG1f29a/2oIjsyPrmlB3tVWMKXeCiVhT
bAX0QChj9Cs2gbKMOknVenuf0ZzKcsThvrZMMT2qUXOMjwsEqILCA6+Be7eMX8P423G00kaeMzBl
iUrAt199PlvH2b/5UF0IWWOZCK4Z4d7M60AIaPXs1JescibEgbnq5TRdKcBLy2ANv/qV+nPVhKJ7
HHwBZo79hrM2idJN1eGtDWL0C4EF5x1FbqG+CNQitrGwl+VYMw8EmVrcQwpz+dVd2QFBzOr9VdWM
5H0vzSFQe7ydSq8G4Nziwlh1KGgIIHzLf4x2np7cBKhfxXf5MMhfZJvqSWdF+jBTHlQjQ4UD+U+Y
Le34QVUX5bfMCqVDp4/NSY9MMVc2PPEIXbqt05Lb6TJlM4b6iZ73WUvj58TO/77rh3JofC8iTnX+
mk7c02OC7XAsfj0Mmnb1lVuekBp46MC5qN87zZDn9UPXyrDEtEEaOTxth0cE8V1UGVnf5QejmCFQ
zAOl07d6Y57kpf5EuNFIH6p6lR63vxz9jQhm4BVh6uxlMVRH6FD4LyiS4roda+KQPwB6iu6uHp1i
5yK6cVYKzDz8RnfhS8rrGHb+4ibo91XEryCs0inaGnQ8xaEhBoodnXbkKH1YffNaUS5X01szfzZq
daztrwGEu6kTnvE/NCVaFBrgbIwxXkGYkuzsFjTM+8D6nB5Fw977bj9f+NXomoNcCoutNaUkhfWU
bKy82SfwQzSVQZtrSFAq/6+cbbnwSzjQkAHBxYOb/LoIrVx8qOrQIF4gf4aLPMCOiiAUWatnUg1P
Cw+rRipQ/+qvCAPBit6xmcTcHFePwxo+GggCIRwTz2TPpebqYNEa2nC/zaLN/5LQjxfDetPMC6A1
9r+wGNmrzv21zsTgylnXB4FvQwYIWVSSVNkmjFCDzHNLEI2VobfHKB4zioccY0rN5GunYrknv2KY
0U7FyHV6PYek6dgDMU8xOGOG8qn75CGKJbsu4BEv/05hcYqWPkR7fjoy3yB8zGqvPoyCF7evzH9j
2MX5f2JHwsMUXu/MzPkyjL0rzP0oOQd3eoPo9fJBHPniOTvF7gCtjEQS0zyNmOVuu6AFBlS75wGW
2XAnCD+YtU0ydSzckSNmYe+PoCQ+Xv1tstnUq4APHYAyh16y7AZ4WujYh1p7SajpgldxIXrA9ojL
1v+q/ZsSnIuEy8q5HtY1xHEns9g2Inie5Ne2NqC5VYDF2sutc6CgNioeyMkk+fjW5ZIHFYQX1w+v
ntEalv3EI+oLGGSf9/RiyfLr7aeXzYf0iZ7RmvluG9pN1WqWvN8G42dnFVifUzOWJb64iEAhn6k8
4lTkfekW03lFYYRKVALgI0lOL55kFVX3tqEBJDnBAdREx0rv0AFvL8z/0LInh4ddscviM7/+q+wd
4LvM3en4BEbZdjXcAVsbtCGN5ZAN0Bu5tMrSBacczLgyGl6PsqFjf0sMN5ktjOj57nqecOSbBz4f
KzMMqSkLKx5Y43XUq7lskQw0gKdO1lUJXjx0OZ+FpyhuwTLtl1xm9WtspLA4HCV83TRkWjl0WAwL
MAz3JPzjneHRqhPyxNZ4TNA3bTX0mzvq7rI4Lcn9RbBl+MckYtOANeifJqnU5S5Q1MDsAt7kRQVj
Ic/JBbZRmrkwO6uVyETwHvDVtKaNs4asSvnFFJOcSePQwKQaHGk/j2R72jYW3D8n3DZyvTbCLUJd
0v+d0P5ZsIylPzm2mWTrLyY/2WqAdmVbr/PMCdtRmSoZr6xIT5cED6rBwlnweClDqHMEoyHiPo4L
e6n26RwZwGO92cGlGRMyr+D9YF6vom47mQWDb+LsXHLRW4dDADUjRZBeL7H6ihPrll37bJiZ8huh
hbTvJmZ3C8u8ZGRGGQQ/Qzyy3A9Ue/i8ktQVd7Q4VmsQZ4KuLGF0CqRf3Dm/GEU6dl5h6ADpjIkl
ThaLBUbPxJaqUSBHK1N2vKuwsCOeSe0jOAVnCNyxseGWmW7O7S13dLFZnFqGTOMpT4C5kt+h3Ufc
JvDNF+GsjTRkB8dWayc/xMzNDgx/SjokzYcNOx4DsPJOa68XrET/tMGUTRle/6aVMtqHqgLNlmbW
KnmtChYgzuoyQV+o9AmigB+xUGOgWjR36zJFVnLy0VOs1du+F25WBq6GiKr/y6JuyEt65jJy8T1d
n2Yih6d9+6Y9EUHFroZ5VXnupvxHmrsIPPCLxATM29IasO9S4CLFJOY2xwRFJUmPUdP2/Uffr2Jl
bl0UNtXhevmDaOI8hnJbYJkhWM233pxkyyPcCiukZkfRGz7NB3i5YwdW48svuq5W1g5anTCl4mt3
LStbwyZ1jAiGgHwAZT+l1y0sgHJfYz9wfiR1u4Y/lIuICBydI6erJF8IDi640BaYgZ0x7FHuL41g
L0IlS6gGbnL14N1ow6ygPFxA55Q6fiEce1oOV11Ytz5JD7tiJuBVVGBJs9bgKoGxoRklnyriFJUr
gm8AuWkekwbQoShJj3GA0GPCz/HBMtkRqc7Op1VE1zWJScjUQIqMgtRlW7k7Pn+iOTtzJTq7VDoI
t2Z1IVdTIXHRt+WsIrvS3KD1Czr/hqEUleM4aCFEXK5ni/nZ4I7YgMQUIQxvtxbsxcEhrV/gbGL6
ajky8yyVYvZFGgtGPMWTCKyD1SqaNqjVTLRdBL2Rte0VEd7ofzduKppOvILvd9IFq1yvVPaTACyE
buV06zecitDsxoaasizq5TWo7F5/hVp2lUps3DT38JpCWnAD0l6bcOGyrvIgVqiie8TjTm9lfWP0
6oTaR9clRfzUQNh7iDKJqf3spNjnK3xBrgPcYkpwj7YzCKdlbibbxUyEhTsJm1DBQBIRklVfZmzu
BPztXJIHCsdVdz++oPcrujhXE1ERBeK/NV54bX3sXjJoEEetSTnIc/+HqPhgFBbveRBsWmQUrRPm
P5TmaFlUfRnTmt3G4E1mojX1FPQSQnmVF0lvsyN+eSq+4X9s8xW6jBDcEXi9e5NYqfIgToVS3ns0
9diKaMsEO2w68np0ni/lp1f9fV75I3iX8hvoibXhyfNJ3/ycOwIr+sbPR/3c4oZS4fNChcmBL5u/
vF2GITBhvmL2UyOaXIn6FWMmphEvVlzZ0wbyhOBKWvlp3sk1Kp+x36HYoCrg5DlQc6oZ4iHfK7w1
B3vIzvzTv7psFUomZCmTZHgiQxW0/fPzfYEOFkiiSr1BwKOUQ7GfabK42IIWlKg2Wq27Wf46Y+28
BpWJutjLRb2RWPRHxVRy0ULOZUoV6pJXHJZLxyO2xM1G+2rtWJYGdicza6kr+RnNeLvw9Hfn/sLY
FtpyImUYIHBiI4s22sMLkaxdl+CY1tCKNzAzF2H+oxRtYERlV0CIypw2lktQSYEL5PcAfR6+cDfE
ExNsoGKdawx0ZfhsWsd0tZTVls7gq/CtnunULFFQn2hyrXY0Te/b65f+OH+ogmLvmERIyL7KsVy4
pTA3WG61O0m/2xmRwWWEU/19Tm6DDzp6yO9yghZpI9GSFVqlBHJ/drT3PO6cjL5UM0ZYpDJt/rv8
B936qwjQ8LyvICUJgPlw2eV89OeyWeggLEjvR/N9NAanTUDBkYfSHkToEbpcJxFoASS/cWGbquGj
u6eMhcaLkuowzrCTGmnuGp9qe6P3Uh2m1YNoEo5/QSElfLawvEwdDxnpnfhIymE/v+m2YPsV+m1Q
gyySgJU6wHFVadp67XMtEBs4TUPb7cBPpLcbMyNn34RzhwlrX8AxNAN/TQAguyDR9026U/rxDIXn
d5RBNqqkWH2ZtlUn+cOk/Iu4qw+VSa0P9cewMuwKwFQREX6fPJvvI80N74jMMRgU4nWaTkNvxNNQ
WK+Js0fVadmffNQBqx5QOA6hG5n2Y0jPrpHX1sZqPy9GebQSxmQSeZ4AWxfNTB+AKifYeZVWzz5q
Al5VvpJZrcxMdr5PZ55A/Mm/+9l85q0pV6ZQrKmakSjt8/cg8MW99ilzTh8rP85MDyJt3fN52O6+
1Lb2/plrFRpjPXgK1KVW9fKjgVoHdv9LEjd9L5xxe2J4hPrZ5VshSXTMy+WTDADvJlcPQP1x5Fzu
0IfGduQhNcJJ5IUaoHFOlwGUFBL33hoOmzgJwU6RXrejdkD97ukxvs5hjJxpOMqe69Hnbf1dsy1T
G+aZhuiv4NFmrhFn9Hi2qF40s2xVDDRpH/4g7gNTgTajj8m13v0PZD0e40lRnc49hSzso7XQRpxk
UKW6oiPhYu9Ed9P7ini/n8yvD+aQPsHDHlXTLHn/x6efMK+Qb9A7zChRbjCf9+tT2J+iSS1KDX5p
S+WtQhXnxvuVtWuKMWvZ1DId+2dh2dPLDyGje8o7VAhz4TZiGg82FnaV8Bf3inOJNYYHhaXQNrgu
casBibe9rrCKqDr4xrMQmiS1gpBYsvkM46iYxVUDnXcRFTr+BQJpAa7JMzMHAP59ZWvDHFTPn3uT
gwQtC6OwprjkQot+SeDU7B8wviqI1X+8nuh99XiKJSFqfMjBoNHPSV8MlnqY+dN3UG5cwLTQ2ars
Sb+TsXVq8oiNk6hqIl7qm82fxoPkkopvCTekl0+6q/9gxAUZhRpJYSdskToFrA1vJ8gebgZSVvTb
5ynrAnfmIOVkb/XWbtCdcZiYwEKNJwDxUPcSOuGAajegFKMDRT2HoLisK+pfxhvbL/3Yz0EGoksm
FfRjNGtB6IJRQ68KXAnzmMa/9wNITHoKCvZCm+Q2EsXsP2PUMz5TxmRyDJIHZvIego0E7mCbNnkM
0PKDvQ8PN2M5kv8BeFzNOQDv2+EmbZmxz/W470UPbiBsEU5l64CxYIKW9JHhGqKwpnZ0u+PWTB1m
03+HWyeUynaBdXEQDClJcIOqqM/EbvsjouDfiYBJiDWfQ7e12zhhixXogju64jPZ8mW49RJag5Xp
dADqEP1RUCznDV59QewsR3wm0h9nDT9t+5wM/QWfWkMA5IoIQLcAz01SjmQrYs/tUcZ0xbkOTpqm
14x2SjJYZhlPQU9cxja4s0edIJaGtEEMMftYMBCwBmM4NynbT0OoWMSO1YxM8LDER5e0Y6GDoesT
XCRzWCnBb8RDBAlOR2HXwJxwokF2VxeiYYTlizwvzRIZf0JHUiAnulBUzmtV/E72SHEPm7RTx9gi
4mfCMrK6Qoh5klOIG5cG7lugkXnm4VUabJ7Y4NesnJjM/zNoh6IzVUDDJMhdn8+/jxww07z+wT+b
kC9NoPSTsssn8lhORhrIwDlE0sfXt/o+cJ1I7Hjtax2Siq9B+5tKQD0jpboZle/Mm1TvBcWSeLAr
fL2jUB6awABONklXm04lKguffYYXOjEt+pDRZ3vmhqF/Vik6IZ4RsXvC1zNpbOo/M08kQbHcuEHj
t17wp71XZu6gKvf2sNeEYbNhMmeMva8wDRDvYVK/pC0UtKxONRl8MeAeS99jVEYx2ivaoHfjdnwH
f+jm8+8gvDbj3BIJpcsNSs8fAAmjV7AJzrxzDyxIksaQzIoF9/XVdy2CxSpB9JwS596xehHzwlYk
m+fTT3Wyubv8r6RSJsV/qYouLgOGl87YmU01av/QfecVaVM1NlP1dcm6HN+/teBAFjGZIdyw4BlV
ghBt4wDLfX9eTc5Q2frBV4amgPSXaTaOsKHrugpVZXZFWx7g2c3ZdqnIMHaxPaWJ6oMfe/T//Vlr
ncU9e5+hRj6C1dq+j/oix9yIZ5TcLAkU0kqmmQwEOCglVF+FnlsqH//WVp5LDBXbwWjlK4Pr5MaC
ev/7rq2QqyorT13ZLH6pP7AYO9drzDzvfDIq7FRBAm4Ye0TOOLpctlNWzfttJk4t3pGcxtidgrSJ
/9ACTk/kp79ZQM9l4u9ALLgJ5C4lk/YojfjwwXnrfjBvyb7mw8iZDr8Pkozn7AI/jMvMQx2Jyvj0
dsXCw9krAx+1TSIO1y/Y6BsVnTNJM8nx4pKGBQTIVdQL3JaEDj0fs3JFkKnl0/043D918EH6TuKA
R9B5iUxPqZTdmZBj8XYxIb6KAE59SrWU5fwhl9BUmGviDh9dpvdNRmgtiJjD5TFwDCZg4kWUaIpj
vv4l8TuSY6GJBiCU37j7J6JpHAa7bA9k3+aYnYrvaEMvcWLHNt8kZwUkdIB52Vm/f1SPGVz6wd81
snF4UR0UVpuxzsTjVYcOdiFRfMF0te+Qh10uW0eTvSQ4nHaUl7LlJORVPN+yRMQqUUroq8Iremnt
HlbWBu8PVrXZ38Jr3RYaIx4B4aI0xWpxaG+6Uj2c6UJmaRsZ0vZO7llO/jnyTTHdTVMP/ccK7vQ4
JPqHGYD7tjgjCoOjeMXIHqvJMlwcKjuWmv8xEjjgTZdVZbHq5SOWAfi9+S+sbhNvlv/edmB22S52
wmGOnHL+/i66CQXxrZYqUWvGbpIez0LdckrTjbbIQb0nBgo+8xC0dpsx/r0t6ZThkxj56JsamoCy
cszbrhlzGCv+kf34J+yCr2dv/A9h+0qWBPS5IuSliNpBRdor47zNlA83On+5rC4rNU1v2Rw14IZx
OVkvWXs1SVMX8mc0NgGhbjo+GXeuS4S1vDep6Cg8MYGGp0QgY6RWXKt/VMLMO6f1t+tC6BwW3p2s
QmGFUSdDTAqAefq7NyNivR+snNOC63mQl+U9bZkdcIa+CGNzpIgNdMdL+nz4RFBxdMi2L/MOBGFz
6lsXdnDMjECIOJ7eCsXAMPKbk+N25DxBLhU1i6zMp2egGj/aPXIWiadQH5pMHwZTg8oBKz+jVhXI
lV7VH4u/Fbut9p8ewocjPhlhbkPB3jZ5180fJZ88XEL1AOu+mEOUkqoVIUes5/PmkQpQYUoRustd
6hGpfHf7dTevzPKmfcK0eWaSvaZ+Fr8JklvJMR/8Rv/lqpjNbLAqPhSdOxsjRrKy7d4zKjK4F/Xu
IDsXGE0bHC0mx322UVTDIdgE+QcFr1mOX9jKVYC7MDLMQcZu+YUGb2ORnE8MuK/QAfKyXI2j+29g
6MAp1DCjQAI79gnng93uZ2/0O2fTWGRFtd49CZorOMK3tB8/OHfaozy/v8dG8WldcNDBVPBPSXgp
SWtvZonDuJAfOfElUQqB2ML9VymDy5EpPMOu/WPgLQKxmaEbOCcRcffRf8DCFuHXxDXbNZk+pjgr
pY0FTpocxN+hE7QWpJnvwGim0uAYBGv1MCa6fVZg+qJM1uU7kHnlw9KtRcVHBR4xUTgw3xImNT+i
9WFsjfmEsRgkJkJUdNnpSkuAdj3o4qTkx7yexPtQxilJkcGGAYsqbhr/szpuN9gp1bT+rTvw3FjJ
6OEmFxkw65/DxeEMxx4kdF1fyR78gztbskzft2h/G2ausS0gWWolWxz5CXgDvmGpjilxLT3uQ4m5
bO45ZwXDt7H7Cp7+SEM4NF7LTE1zXXfJkdQTa28gNj7kmqW6dLuHp5sVhmj4cCeOAktNaDwmGzmm
TP2PlbDAkzwZQwRSJx5KMn014+B18Y4I6kLvAKJcykv2Wd285ht4/I2086vP/oMurIzNVrqtddL8
hitvWdEQ4UjWI0bI0+RnohIwd5Dr0uOXFIB2HwszoFaeGuXJw0GGbPhQNFE28iguutRuifg8siBu
jeIR95ZzX2LUxucoIOh6C7wxpheEUFzeY0+HStnhuIUUuggqwI3P3Sq2l1Bghmb7ijbuJW6g2rHo
mC49pKIrTJy0m/zPLesoJlS1/Sg3Or3GAxAHb0OvoHl81ffe63Vlk/dUPafL0vtExOZ8qtm7di82
y00+FzxBVys+i+vgHIDZQzjYDc19M+FoDIp4E/cxhWv/35EvaotySafHjB88ucW25j/sBhv2EcjE
179gwA01WRmE0Hs3oKfMeNjPxsbwpQE3uO/birSzRJVmQT+Vig+uk3TjPomQYRI760OxKZU8kyL1
OGppx2+yOp+v0RTOi+XC2aMqksi/+4GWp/z2lrkIUlIyGddIZCHknYkfQdeC6sjTEqSsK5OXzOri
jVASmPwLmIYwlIkIIPkHx6k0wbXZBqMePlG0HXeyn/zaSYrs6YixFUHYa3mUPjXB12Zmv+SKQSPV
hgYcv5pWYgPvJJbx6G+z8QGC/FJzz88FM4jofkWje1sETpE/ktmcXFUCdRNWgg0oCJxHnqy10col
sustY/T7DCmlscMuj+ab1//AVJkKaaGk9MGvaukUQNFkx6pxuzUH0TB8jFhJkbE6/fumzqHNMWbH
vFFd63DDuTwgVnPqSEtPr1zVGjeomM0/7809hHo0KauykAjS8kHUC9BP8l7JkObDu7HX0b81joYf
hVau8AthvZugsYu1UiPneegYFt1Ajyywwd6FOBo3MGfcPFAzl77dDgWwiWBE0AwFeM0BQOJUGb+r
76MvntEYjFpyicPz1xKO0BMI9U+jW3aZVj4hOG5HOICtzb+ZwbH2V0RReEptss3WYveawg4j7zeu
n0BjLxK0/27uKtrQh1KX2c4hl+Cs7/AfuyEVuYqTleNHWYisY8kj04x09Sab7BkyL20w7bXS61zx
CUgDIFj5ekQ1WTcU5ZizGcre2qcEgy8fg1Ngy5zY0BaNCYOlMUU97lRVDvkzyonchgpB8vqD6UWL
8nqvO5dlbNSG8fU5wKNZ+/KpQEVKT93Xv581qEAV/x93eV3fYulJeQW9tLOJTw4hDBkV26QasV85
szkYNzcILA8N7bMuJnPVS3IkKoUkZJGGyb6d/+pxB+rySSG3PXeYIG/y785owpJEqfjrg8tP6pbb
qhg0TynzdiyW1AzodjayTSlAmUjUmnXu3OLvjDM8YeW+IUzp+RDcppNC//i9mj3NQiPHr3YHThJL
CHIZ8xn0pVE9dY1z/j26ABV4zHl5aaIJMki2iBw+Y7qu0QXaXWntzsI5KMgxAvA1tgHJjGUOiCNt
/10pGgtxWSqv6SLdk9OY5/WP/iGMY6z5SoBV30g3kSYTYUpFdhSS60xz4kCb4+yH5tZLwZZtplt3
rvADK/j2heg824hP83sJ/tj9gNrNpRxwOsg6Bs2OYdV2LnEokXhchu42FxzwmvPMcsW1l1+0ksQX
3RhYDKQnIwv4r+3qN5In539/jD/MfdYfQE6mzoZAzooo8hQYf88EnqHNVYDbT9fNkqAnfAlfwpF2
6WyFm/bUm3BCYg6dHfWTStXR2TTj+YjtJByQtRQ8O03cKigP4TfImzsCeXI31NUk024KXWeZWGpH
lH0vGN3sXJLrAhK1n/zgYwfebBCdVWzq2QW2mZiCd3lE0FqgUWmNOjxtU1J63IGr5yHxPPEWmxoB
nOsxLGF70zVQ36UEaVuXOXT18nFkzu+Z1N1Pmp7cDFuSYkKcwZX0HkrzgCJlA27zGDMWIjzfS3uQ
agwSSkZEMJ43uJy0dPM4DB2p4d1MO8+zmAlCozH3IrX4d0c9sbmH6Pa7ZbCxIN/JfxX1LbWE2WI8
WLPOY9PzmMi9DpIvGS+MpM918xXRr+WE+8Vr1VL2IzNZth1eUB1te0B+LDMsiNVznGSkkpisaMni
npIOlgDmdgVPX6awL/mEYrB184YwjcyuiH7yvb3cakHa3OAr/G4hKiV4aBFBFSKy5KQ702wsJnT3
b2aFobgsLiizsJeuBBDlTKlNdN1RNOe3zQ4xr+b9gxS5U0f7MlzxDREpNHt6rTdttHyQRJrtHCMM
u8wZnvppKvmWpEVCFsq67z6sCb6KPOYP2PMvdqeBFXM5ymksm2fHBLEWhp0qx+lS7147nz+HWAa0
7Hu6Py8y3wb4kYbxdyaTMxL7amezLqhdZm9PIoWM4kQKRwdPaGbbYRfOAHe9p4V73plXbBAT9T4Z
NOOvxvpSgr91BHxO8nVrwMak/scjKo7x96ybwQGjgKPsvjgOuIatyehtKLyvoBe+pEs34XCNYXGX
eGhTVM1IIxkuqMXaoTRyxPND/CY2A+/n164jpYmVg2SnsiH22uWu/yUaVaVIP2Pgc29qw3czbec9
wN8Yl19gMC/xMmdxrUro5DpP00TBshZJL2ErtLVHgI/AD9Zo6lmfP0JayZ4TVQJOeExehwEN9/Fd
Si0AOX1H7A3Q+EyLxD9HQw5gYgFmsmQAoRoPLF2gylrstaVx7nWsfGOCyZoqGwhDb5a1hwWT0VsP
IpFFkWEvz3cAg+n4hScOyP05xQqI96J1nzi9iWGgOdO2YedB+/F1nta9U+2WjHApajZTG9ICzhw6
7OyEFzULho2/Iw78UVOUGjrQr1MVfLkiWS9lRA9aHIddpuBfzDa/uZ6x7BrGphglkMKl5N3R7sjK
oEeBCXFOXnGbwYFLQmnYsnajTfg3qa4fXrmW+dNkDQRXYhSeACHzxSL8vBeFT3JGu0A3ujVFQUW7
maBbxZOzQs1xaRu5NDWYqkC+aroGl+IWnuaPpuribc55Az3yDvO+VrwlCIaFSmPNk9B7Fq9knLQi
EbXWlgw5MSSPAlnBbf3ir36eJdYiePYi0IO80ADhzexVhTJ5ZRgyyuZGRHltU8BcGQDIWM86stG/
fPkVAAIMSillwJG84FVeMWC89ApyWQko7snyWjBhhiaOBE46NwoiFpZxAJgxLJk0/oMu/fjDxl9z
Whht2Y1lU7vAcalbMCBe/CT4ZZU+vbbXwhfHw38XxZ47vLDvifq7fZ1rVh/gwtn0t5EXUoUZRVET
sKS8d96qIIcxZy/dHr9WllwXtelheW63UCty0f+G6WlqU204hNdSQkTQwWuYwpDA+mHS5mQZ1uKb
7qufHAhb4LrhKenhIlYDhaUlx9KN80U1trTbpK0MdIzw6RtH3IMDNz4aR5dhwSn5PyrQxOAW3J3f
5DqyyRSxWYuZuYsGKWoGCy31UQfL2GYboFsxeq0RiKwv5g6VU4SqhKaMms8xZnkAdRwqMNFwlHkL
tJdaHy8Qd7mt0Dr1Hhak+BZ9UkAqCimACeyag2zrRWJTQMUcCtedHFi151SoyXhSY+CG+YpaiQvx
5+I7iSRjBRbnR7ApeG/ce3+wv2qsmMK62Lt7cHZml1sVA92t0ZEzQG09kjw/19Vq8gzM/a1bEbo5
JiUKsc6FJ+K8dA0IEl1jKHkObx3LsLt6cRPfNMvOO2s/Zp92CDA3z9QNvvKemkClIUWftF4AEd58
UON7dlp9nwbZLNE/z68Qyloscbor4bJ8PuOmRIEwQSMIrsMRTSPYRtMZ/4O8hLy9EJDgUdf5eeTP
9bYAvxtWJgrYmPVlcMc7hzEA+Ej0/Yh2HEUaOdHVTsTP1HQphPLX99fFkzmiIUCqL1fIapuhqxM5
81tGNlF5NL1tJNnVWzSaSGsNlXtttsUeFLIhQlDm2OIm8jLR+dbVxQyN9GO/gGK9ourOICfdCPFD
C7KfgIB+22hVakjlpK+eO6WfvRDNHVRs2WrGHl+DMl6Ehi3umMbVP9GVEdjeX5KMMsN7xUiYO67Y
hvywWQrGn/Nz+stGiRrZ/fEvDa0T00rsTg5Ya2Uxp0/kZ3Dc5dapVor+bq8QQKR9uJxY39bW/ybU
JJZUhOJV6j7I2BBXwWKuXZp5zLZTc7dL78i0XlI0PDk6cxI1kH9y+hq9bZUN/PH1DZm/RUE46Y2V
rEqVUgcWhw1tRQqB7c1tvDRWWJJGcjkpSnP/eImFMoEHK+UhpNRifuok/30xOh8PvdAKfRJarEW2
JkVLSnxznebIBKBwjOZAlikQmV1JzuELNvku1gzPLqAt7tJCRWcCIg95MJo5tDat3SGFoutuSLDI
jrSIIuJnzG3biNWJV+af/zWv+Z4cUkgog3CMZWlh8L36akf3Ml7t1PzCeR5kichL24T2j4SrpO+i
STVtmMA3Fibp5pKoByxnaZky0eX68zWE3L9qC4jdUiVS/aICTWTGfQxqY9EId/5RaEZHZzDv+k0m
5gcT3mobqba3Ud/WJq632W6oeJdsimUVmDSR5IzW3mINgWiEBfRVQvomY/4uBrmQzBfSZW7C16QG
HCu9kASJ2yl60kkV/PHztwgghoYxx/qZzRapbHsJusAdvwgXa5SncFuBJ56F8gv0v9Hcd6n4Qwv3
3hO4c2yur6rw76EeJV2Lmadpbw6Mm1SUkzATl8jP+keoJW2sneih1QFa1Y36xTXboHTnEDsvu/y4
4kTBGEGRq4WlwjjR9tFXCihcsm0THjlew7W5Et869taA9+o4BpcwF0CLJa+iKgZis9wy1pqpGdOl
PAcVKrG7lwTQxrt0r2CvhV106CeMqIM6wHO+BarwOkNSETOI0tnKSkItS+lkwqFdC+9Di+jJfdhA
ZGsRq/n5X375+6pPcWpFLjtoIgnw3oR+NO9gOAn02QN1Rta+0Aq18T5e++P1oCAUVrZz/afDaQQh
06osBusZx6SSqxTv4EfMg21zNPnsv4ZdFVSxkvG6Y9IptdgxyrWQJ7Y6J7mD0YKc7WyivW5Lo2HB
V1/LolK6bYrSHXyBT1N7L2/S64syx8rlSs5F8Vs6WGBqVwMPGjYG6L88QdeEpzMbPyNpzfSfQKd2
e815bSP1d6un2gigUQeCm+IUeTxS+FxFtsDfY86wYw45cYRr+q+4NB8h8JumaKKNDoPvc5MaUkcC
NDcIfJSfXu2ed5va8getYWxlZgURSc7L2wxUriwYtUH8aWl5OE6jX7wehufzkUQztCzlSQI5UolR
MTcBg2DUp272bvYNyqv01Wdvl0MJ0zy3B4/Aoaeo5bdKFpYCYQAivYmqFh0R/eOqOwnu6XwJKXUi
oIUjaVoJ48tcbOzQfSgjvHp7Whv3doeQtbEWWeyOEdJ00LKbb8MV+CXgac7vvP/OqIm6IWE/73/R
UrJ2LruI3IL5LgPo+L2h4NgETbk2joTfjRmd8jRz1ave7TZBPLbYhsR9X0xcrzuFS0HSSkmiNxY1
JfTC0xPVFmDmC5nZtiZtLT1sOkb4QCks/+Se2TJihMs090ln26NwVmgNx8oSd4tsljdVfLpjgvUu
K7XRBYozxqDd/B4PLcjg3Mqe6gc8d1p+9gqVQ12/JQhtPO7BantZDUBt2NYjSa5erngGbdtreuA+
cDb2vRNT/RFOfP3skkN9wBXqwsbaAgnWBgSeuKSRVcEGKm8ES15Kcy4m57QPt32fduc2cbqJumyJ
dRQcCJtNUmdbVh5hYKD/uCKt9obze8xyOO5LXpqVGmxvjxBh/CEBFmGdtnd7gWC0q/eAibf1QpJ+
AacTzM87AEwqSkT60aKULND8XnWzKJbzKpZLZhG4oJeM1r/2xwj4oiYIHKlCJlYWskO/93FWdPYi
nM3fRLdm4rzWxD/EyK7rHgqi+/hw8QXX89zvh/6bnN5qeGmhUwPFRHQfjAAjui4HjIEF0uqPz6Jz
vCpz/o4KCteeHlMGqhGQwIHQya/iphEtCQhJqfjexfth7bRRa6j1Gv4D4R9uZwymKeufEaSZ/hCV
QnRRxmsvuu3Pll7LFZJeJlrOZvZNvBT2vbGbOreu94+PFIRSQqeI3j1nDO1PKKgGq5IvZC2mS28R
9PJzsT0fP7Chjobh8tDP5fXxvvzTGj4+5/5zEhxVZEnaDvK6r3QUD68z4EaPXxCjXVrQx1+Hz0o5
2X/IEYbD3tYUT/MRnFinjqt+8JeSqtwISx390p+JHOZzY4NTcUdZH9SRi4LtUcI8W2Gs51Iog+Lc
Vjag7qfVqVrEWwSJ4jWtBfTgD0LBaEdgVpXWu5AmBcqa1DeQbrLtdnvavAec1mNq1gurSMhdvSIG
Fygpcbpt7eoZFc9napBCcLdRvbndh7VQnja+HaJXYYobDnYBQ3pao1XFYLUXHVIJ7iZeGcZ4flOh
ePeKTAOacXAxx32LWPGVl/xMwetL3npK2bn6FQJAp/VmXxffE6H2Ys5DqbKpEEMWZs62TieHjr1O
QQ8tcHiCf3rM13OU2Y5gDwKpfDgAUIkKgxvCwkRqnLfyKMZFne7auA8mWOCQpxanWdX54xbu8JPu
jcvl4FffuYsbvkj4KX46DOQ41rpXIiTpAl70cCqPy6/jroHejDDyCRpt0lmZ03lWJ/NG/y2UI8Mq
zEfNvwM+WDpoRPFoxKim+hbXP9ALo+lgJVDHoVIOpeMY9tU6zVmen24o8JB3prTOqLf/8ILtAcGr
DO8B1+VMh5DeIH5MsT0XUNkFZ0rY6WuDrdSu3rLCePrjkAvmuJGy2+mLvRXkAVdd9uOwaXpk8Vf1
gDJU+O+cyzpl6g7z/s6V3LEDnmJX2Wm3Qmj9nk2szI236AMuyWqyGsjFw86f+rNjdds+tJAqo0LQ
R/OW3Qet/YdmdP0AftpgD6e/qJ6WkfLz47wuyVTTArbeZ0ofUcAwvrgH/1MTr5arHZQ7dZR4NqpB
41qo7aj7et6VzabcKZW6mSa69qfuXCCNmhTpAwWE6dZeV3IR1yQZVpYwtCcwVFO5vnLKR72XFnKR
rTfApD/N+LMd6qsPcqxpm7gtPSDMnBguKUSOONyrzkj4KZw5x9CUC/ODS6M92hSqW5Ip0RvpPMHZ
pB2tAuV9OzUzbTWrI5ZDCTTKxJZCzg/hymLEoGZZEiU1XNG7NJbPorRCtucGWKQZtNwDBxeIQl1h
B11qdcrk986bhX/tndhY7N5YziuMlTAli6bJwLGdL6gdvFZ8Ye+4ZmkoSpJ0Eqya/gKEoQaQeDLe
EFW6ygZLHW8x9Nf7Izi3eMLKJcTU0+TXfOHPr5T2eM7vdcM4NFoon9AVzpoL7qwaO358UthvDEk6
ZNsyGsuRvnr75zYxgeFm9tkCjW9L+1O0EGCdcy+cf0VZLLLjN1CyLDR/g65u2DLIj40Rh1uFLmz0
JxS46sadwAHRTrCMPxN2vu3wYcDU1dxeTAzF82irJrhS4G/Rh5qdfazaAcCAx0ATErgt5TyJRs8o
KoT42L6ZwmSgUr5bWIRAf9DBG9J43xf21eknQjSvV+VJP1/Qez/gLXcpHxJDJ2Fcpa8gSjnfRFFf
E+8JzeHZhnfOdk93ScReB8udC95E+Mdx0GiodjtPW+vbYuZfO/rJfMBraApBTj15epdA5LYwCse4
Tz5Xhq7puecy2u8SsnUsMwLZj20Po//Gdm1/1pZxZ0IqpdMRLCfsO8OLkBOYIJoVhsdrm6zUW3UL
dw4DRgOOyFejcIWHvZfqLg576tvSA3hatis7sWVPJlgYJvIMp52xuiwcFnJhy4/odQ3WUUVuN08R
86lmwCJApVlIUiLOy4qKLpQC0x5UdFhTptB4oUyqJJWNo3ZL0am0VDwKRDstGStwmKPIAlAoQyRl
+YPiDVu/ucNDv9r62d6LkZDV4cZRh0HtNBFI31FhfI7KzKYiueMDZLJKaDpccxFfkCOU/xU96wF4
aZkb9DgbYm+PatLqrLToXk/UzAR2pkABk+kVW6wlA5xwroh2zwaqUvuyOdVczn/ilzkuOX290u0A
LcliPiqBz2U+DGEpb0JBwHjZYKhreKWzptkC2rgim+/l7GrcHFRoC64wmXppm08Juysmcw39GT8K
4iioUvn87xmSJLSZhu5mQbBUwNzylu1AfKEgXzDnyjU/CPFLhEbeDbXjm8H3XFHX1mY9zGBl1hVC
K3Qbe66WRXu15btN7z5MGmnZvfrjuhvpebvCVFXG0Y3J+F27HPD3HbhGou2aO0W9gS8XkThO8jQK
eThpljuMLE2/iFymz4K5KxyUpELQWcCSO08K1bN3X0byy3GlqC6804gKWp5MTritVo77VUuzG5gU
BIV3d1KE93uEKjwuVKyzhdReLHXjL07Es556O9MHH+69imGpll7vYmDHp2CbRR2etN97J44GAQgr
88RCf4quTtX9NETBOLEIDQ73cCrvY00CRviy8gpHvZG2hRSiqNws5LeWZbLL1Yc87Be0haNyauaI
+9gVwaiChowku/N4u+pnKYMoiNYpviyPoIU8kN3ANHb50+m3hM/LQzoZEPpXOYEADHKCl9PLEPQm
uE9uVsQQQWEvzjb3aL+qjHTVV9evwEzvBJNdbZqT17CRQjxSa8lnM8DLghQ6DR4VhBuDdBpYFK/A
bJB9zrzb/kVC4+SzUEryok/xEKa/ykzdI2EXK/WOya8WGNmTdfx54Auu9ex6y5kdDTy2JyON/wiS
Bb2dBwwJd6BzvVUEXMSOcPyHJL1dJhF9aCu0/rTjT35hByw+PssmBgru7XMDiQEzPmvjMJNk1XcT
65UGybmZb70ysFquFNQszXKedJXwHnYhtKKFQoTn5z3G3416WTXok4tYk7pS3yNswM1LlMyGnUy+
NHg1f0Acbcbzx1nWcfmozcZhaBA8UpgBF/JY8styBvBmJIPokvzfltPlZWnjjG61Hf0DIgWEN+HE
T/WK50Tyee8B7eIyRKe30hVGIA1lTytHxNvmKPiNUMoipmf5UCq2geVbLeYb5OmKlQJnnZSS6YEv
vBgWlT+aREwFzc4HXFHlU4SY2SsqgS0nyvdE6ZQ+QzWAVu4Moyf3ouXvF5E+C196Vl754lXHYE7A
sRFBCqcPYqQUmfIJCNnuN78iASsbA5n1ghkx2iP2pbjzZjQVtn+BhVqa2Ks5QY1Zs4cibUlXE2PP
WD+irVR1rsxrdzRi/b9Pza6wNN8Qw0kQK/3p42GBPs4jymHt/yRQXyFvym4xBkgvmzhHXK1MukoL
DMZblqJ9Qz7v+D2QmVo0rFmRc3QA2mJxQb5SarFywAdl5aNFsCEMNFC9qfvxIeF8ZXp2G18u7ron
T/Dm8spBXTue/91uFdoXlelStkA/6N6P7Gmns+RLsB/mXRuTt7f9BuIGuiMehRkUhND4bBwT/txH
rw+/zlrSkXFB+Bweudi4F3WbSpRCN2UHQXoRujF3O3vS/HukQ87r8vTuOtjTPWz7Dq81o4uoHEei
e/0NaeZl6AeEk3gw4hASt+PenxdjpVDlNEATX3mwv0dirobPpieUGRp15NbNvBDElPnQGP1AUvaW
/zztK9wPnGnBZ199kIkyO8TTizKBz2Nkao/y7lyXADiqBnA1OcXFDvBMLW8YyQhqPk0EMmgOWHWG
qQ0HT3MNnRi8UBouQS0X42aRLcKmhSjZJ0EJUKuSvJjCOvdyvCrbufkSbRSj7KW+xXWVBBPFu5kr
4qAgoZsxrqcyQHwmzlsqOJsZw6o2nfHVU5oLLAcxiBqtZv63db+a5jrIWD1+MbCx7kv/zu58IIuk
8Lb6E4kThW0lWlVpDTt0tL4YCJe7aiY0FrfzNpMrEOiY5kBzdQ7RrmfSyHVgJpqMZtG0F/Ba+yQ4
xkDgTvCQ5Iu1ponaCsv9WAUsxh4V9a+3+kvkgkCckkn2ddw1uPhfILAZZBX+Wn/ojbbe/Nz3oW9U
VIR9g+bR7dzuzy/gB+lwChttJw5PTpgDFniy70a/RFg0I6fgkFzA+S9xVAPB6GGIF0By4B31gFuP
Kgj4gozd54WrHkHPMVxPvzc0PWZc7INs+kH//wBmznlJZABBOYYnvWhgMofYTXP3rsEhzGLYdb12
HD6KMWHa1QTm2yIW5SN8MoVnvCDzIgr89Po5BrQhVn1UN9GIXkgHYG5wQHfgvmCiv5xpOJwbbLMb
ALBbDIPGEf//mTveLmibW+YFmzTHriFkVueaABSfBSGJD+6qbKobzZw7meHFj05/vqdIjLd2u3eR
9YCRJHRqnuG4Z+AZi0+FiCqz8u/DqswMJvDXCCFlmJ+lhSW0lZwEGIhX8YPUz7Sczq6LJa3z+jAB
XjLIo2ChGd0x/hlKLn33lS/U+wQNzBt0EOxTyPjTuP1l0uV8LYqAbnfIlDESGTgFKVDos2P9pSeg
Sx5okqMAGTkzIyvfG53B9FwAp8Y68VApAgQDPEKVYM+PPC2yDUMbGcS1b17Bk1d9x9Ap6JE8tnj2
Xg5DFgL0GrpNfMbkx6sJxtZOQm8qU1Q1uoweUgsrTrqAIhcFYNqn8ajNupiW7pB3peLAWOlzK/oq
zSQ3AzY4X9KSWsxj1mOKS+NP50sd7UUB+A5llt8M8YrVc1TskCEvNf2Ge+XEfENhzy4e9hhYWepP
n/s1+6WNsxOzPfXfoHvqGQiPteT3UZekT++qd/0tcoalHLSza/xf0BLbsO6dMW1L3PDDGi9Z2efV
SjB7hOxwxVuFvWDbk4+0i95Q+anMvQWU5TkEI+1f4SXBm1F679/+pmzzbP7/DgfrqniSW6JiWerd
GcNRl53P4V7r8Mi98yUrIkbnOZN16BfsNRwcsB/e3y+ifn2jtmCnHvycs3ggRB8UoR7mLPwHZ/ml
dYOLqSvFLMHx/7ArtwbWxSir5gsiiZO7KhhTrD76mZ+6WZCg3LfZJr/VOHmhzWjSkyLuunu42kBx
RUjzrVgyQ3ncxb0kCLYJuVW7sfYk8ZO4SEptuQkJh9xO0Os4uWFmJFvx5eR4k2T3KeAqCbb+tAYl
rGCNxhawwj9gKk5J+0E90MjE+bfZ1u3VCYYU7C5foUWuY1nETZSK6/dNlymjKEwH0h3juHU8VDVH
4G4Bpl3aFGB8lU9FYe6+ApWtjk6udBUpOEZZrJrWs8CRLWToZzGN1Dr7RN5Q76BqlzpAj/WDyP1E
wrDdh3M4rsgsuuVkSm/QkR/b1RcWpi2Rqu4GmbQguLcTt0GA4rlQAvLRj3PvcplZsDvT2YkYZJS4
sVs0vBWVC7Ncmpc4X8eP/0xlKTyItSYDHySCO8nSIyQUgbSEggDN+eKsrDMGzf5yIHR3GgUaKrQY
7/H1z+7Kg79rT70cA/4jYx2cwIBUZ2CxIyntNT7Jayqk7ldOJfUqsZ5GY7+lr0TId6A1v+c6Hr5D
v2wceyQDeGFC+z/oLiNocUHanU/YOKLeCImK7uPZ3Bju+FP9AhFcoH1nxtsHk5H6iXneBI8Wh5qk
dHrQZnojM9esjWxzilnUoIfQLXnZdlJw1t7GTsOnOClU8QepzJ/Sp17WoFSG6hktQEEhqonxALnM
X4cb8LLBxu3P4BVE/qftoKH95Q2J/JIEqM9OkiDQ+ScbiDgj1LYS/6zCtlAJ/IQQJwEM3T0my5a3
SIcA1Hsc3CYsKImAZWYmcaP6ax3mvp0mpl6+fjT+c3hhRvfMEBzN1z6hGN6qJ6BWlUEviZ5QA0QG
sfdjgOWsVvPnFvduQ9+3OUDXsXIvbujrXssnnwANJ4Xef6x8Z8YXCKos9B3XzXK86A08EevWI/Fx
XDPhB5W+0p6c2JUSLe0Ot3sPX0d/id21MWO/ojiDMwKAaGqogiZ6Tl4CBeh8IkwSxDxOBDsi/vvq
Ejk3yAX3TQg1jOOiF6ViNkKvIoNUZR9ITz3sm1f7Z0ETYJxnmuAIJIv4au6ziSjml0RK+tAUnmbk
T1ZSl6aVbTJF9yC+yHBeUs3EedFOwSAAvbrrPa27zNwL0IKdPhXP8zR9KULG8bpmJF9pAOw5zgpC
bRTKXeU6yzcVW/0lv3eQRUJWtp+iwW6wmGak+4ZWmvOU8zCAhhGkMinirQ/aEoeBcyZFbeJb9bh5
OpsVRS2tPifZHXGs3K/7qxD5V3g13PNmaivU+NRZ4q/W1P3uLwsA5cMMWhEZM93Cf5vWAUL8eung
sl0qiHaYrFnJCdXyBIValI5VhKRe04RLsqclWADLzWhKET3E9Nl2unC/fd7oTWbkqGXGjy3+6KbW
r5mP2AumMd3HaMg4OkuAcDres76E023EgC4BiljHxaRCWyOMOU86g5HSCxrak8aFz7wTna45pXxD
qzc0owlwJKPrSNozuuEbyTqIHMDx0bx9+ikpHonPVQZy+qxQLPjvuy/Uc8h4H/ZF5m2t/Z6Uou3B
uriOb6MdPmHV6GMrMDIEAgo61I4/UKV7qTI3VHyHwmlx7a2MqHD44zB4nW3SGaaq5H+pjw/rdFHH
wKoRk8HBzuA+miy3wSXEkykqqUV/+dtj26N+RHmeKLrYU62asMDoqVzdrU+4u6dPMsI3H42xa2R9
fQshET7BwIVJ7YJmmUSI5NuN7cJDmNEIv0QRyNT0O2eSqh+pDZzzO4K5THIgCZKkiHglIErRp29Q
QQPxx9N9qyBbgrF4lw8hqubzteDWoCm599ce8Z82xGFiYKebRCf9IROlPIT0fr3qKkGqLrW5sswm
D4OUe0Z/BRAGJFhYcXgy36rWVLQ6N1wz5hLyLHBAkQ216GlQ2iG5m4N5gJ22iWgt5FCdnapQh72L
OABbfxaPYI0MaVZcTN3aHzdEjADa5qHez48/lgTvXd24hizblEXTq5u2nB67uHPLorrvyGBG54e7
d52WNDNi9y1VDqvNatYIXB+9JkiW2P/6wFUtgv0hLMbivAPfNE/Vum+ITunJGyx1CiUf2/c2+HEz
I8Bibi3Wb5smxwIqbdi0wASBppX9ZczormI3L3m0e061S8g80J0W38kjHmL6mOTaGWaUmZoQvsHl
W/UukSzTT6HSJpuc4RnQ6kEHMgddfvr9Bh2LQD0tI0o7KLRw4WjcYzgDHwETNoXwjqzLJBvMO6TS
Wrf9/JQe1MFVVdukYePMZA1tnxLBn308tWu+PCeXTn//889QvBt4KDLm61gFAnZOs3T9DLom+T8D
BsIbWTzwIYAvJIEEVcFrTPal03TtTuYt/cFhr6LldDQz8te6T5tmTEjjSVDREnFL3kdztTbOy1kw
ItARLx2PHWKy1eHI9MxvbuJzCI5z+z97AKJ3RCJItAavLGKlqcUcSSLhYTzhsYOJCqB17pjrzbOv
rMaDos1ePgMKeeadI2HOYBDwzkRyZXkdXgTnHNujurt/Dpz+bit5Viu7Zczp+YoTEGN21s4PUtCx
YQ5V+iBKu1uRTK4Z0leGgw3w7ijktj6BM+VcD7N/yXwt7drX1FdF376xvp5sWe1RObkqtqM1LHNa
c3QFzen1DYO3UvtR5FTw2DDVEKl+7koEQuKpN/5crJG2u4wZl6ovF+eqzdEAqxByA1ib0cwaRgFr
zVtj6h6t3LVDKSUId5xqRMas85LJbSWIWQcKg5goSFJbWuXcMxUbP9fHPwb+NXW1ANXergu/mZUH
z+J56ImJskdoFdR6juj0ARFH/4c+oyoNy34DvZkgkXp3oijTHTU/znVpex+f1Mtn6rSci9Nkkirq
lG2jpHiFWqvTGBSopcaqMescBRFcQUMUJLT1Onq5Fsyk73zYkIPP9VCqSuT1WKjlrqZn4i7I7/Bd
liv3+nr/a6j3GH/xC654B9Mj2+0B3DPJ+P+dX3eRZ/NZDDrg1crPeh+g7Gp4q5kVKw7hWgo3fGXx
VrYLfbExFIfBIB4vPGWL8Niui8XhjQvj8V+eWJM0TBT8uLHqvtqjx4GQ2b6pE7UmWYloOLST+yJP
fv+tEnIBch/flb1othNajcZLo8G/tVOkTNQVTc9jDy7rpQ5KeAjqQBJoOjD6VpMxwHvXnyYmFiC4
uQdmKQLluO45vxsf8BtJSOqKfjQzSeRsnE73Y68L+JM6ZhLLvMBU0siiIwkKi4OiuF6Cpc9Qn5Ex
rXGsdo3IfUah3foAD0Wdl/5rHmY2Iau0bi392qA780dzHBLKlgQMFi5vLhMO5Ml0DUebmxW/MBsO
n0Fjv+qW6dVkaPoqn1Izvsgwzmmu8ccenLEJ0b8tU3L8EPBZG+Lwr04BjjlhN8lDI4g9RQSNvWat
d6/tAHDHBubUPdoLtL9ezUiuCJWDvwE7awwTd25L1QJ+fY6ireFXkOJyfD+PaxqXP1nTegfiN6C/
VAXi5enc9qvDnKqA1VzbIBn7mBMugxTvmaYeDHdcd/svEEq0HyrJYQo8IjjazgSXxP4TdPs/05NA
jWQMN9m1pWBAWi+QljSmcSu1doXrFeHwLNaIwUYNU6hDtBqScyql4DIrWIXM0ihw9q/aGguqg5Ml
7CtP+NzZu4lxeC90ATVEYBOrYsf9MFFqZRCxfF+i+SESub6A66SHLizD1nOHjABNrbQaGkOmGMne
4UpSJJrhN7trZDmZznNUZ2XfG9jaWFaAvroZiPQeRqbyuyKtT56kUcOLnHPlhcBxpvCy8E2IEPk7
WnPp6ghIL3y1APXrzYSNhjz6ErJxiD0Fv3x2yxvVAGbTRALkx3pWObYj7uXKv3LG7ipplSMHyOPJ
fCMLbFLh4mCx1MExE205vP/FADBJU5t6sFSW9FuYtSyOZIlz0A+41BXG+axbt8jvIlYWKgsYeygc
ty30wKGsNRUc4es2+OcNP7qgaUQoW7pF1BnmTnwNmZryKTOW3O+F1Y1tUp+GhbQpCdx5z+dc4qkm
YzRCIBZT0l+Ig8VGMumuku1a0olpz0SKkrU6e81+fsE/ep7nx5h/50yZHu1eyzR2AVz2JK9XZMvp
6oMOzx+XvS5QTDOOVxQJZd6BS4N6aqhz/kFEliwDcv0ICcwrNKySOhJ6KtIYwgzhkRc3GVzCtfgW
wCUWAcou3stdhg/ClL6YzrMZFYg6yLDg+kdsO3FYbdRLm/bosmE7gnZcYW7lplM9YWsq23kQZ1ml
XcfpvM854QfQ/+E9mTiYXTDa0p6hvI9qKkx8mfMnQb7u1ZU7w4Q4zo75KDfzcB4coNghMhCoZP+/
jGbOelxe4oJbSHLLQOT1YpeQJS1GbGT6clLvLFNwaQWbQgUS272Mk64SUKpmFhpmOnb7UPa/Rb7E
qDaAqQUBa69qU+2z83Wu7U9CQfF8VOM4F+ThNNjsGK0rTiAi1hSEHtXlKCEHzP3JXJHY0GnlcfTj
8AHCxEvhsoDB+MGzyv24+J8+cuCvVUvqsilkaOtNZ7gUWcypr7tm4gcGDHGbLVxgjiSHZ8VgB892
fg4XBKJ4qVNpd6s/Gf29lXwYKm8dZ8fzAhHCNoAvAVkoZFbAaR8UM9U1zOizDxEBGYgNfmiDjThr
IIcQCSl68GNUQu4Uv45+CEvsxfA1e4eMhSAHNWYXBo9hRdbdV3U3DVe36/sRDZhHv/F1UwBUNtBz
p37Bgb1PjEoAFoBZ1NVA3KKH6dSQ7X2ti7Hs6ZmwLTL2bh3y0U0ex4Ro1ML7nvGbANnTA5N6X9hU
pMbyNjkXbFV0umCTQug+zWqic/NrnEPjTlwXz1+2OUPCDeQjUKLRmyHGdh4LLH96c4CHSAv13/HV
flim9kaRj+DybueBPe2KO8D/scnwpIAQXNV61TrYu1oJsyXpbqj6y/KpTP9FD6ozcgicXfMWB4SN
nK8YLignzlfG+vBl+DgivD79b+tKjh+dDXF/kVxSHmMo42az8+nz5WAVrmtp4ZKoFCfdFGLrG35d
XjIKTP4R9n9hIf7zbczmxzb2M9kwWNCUmjNFX9tFu2ezjUBmQoGeFDQsVDHiEeIoRT0d4/3Ns0g5
CqJ4Y1pq55VN3TZpZEHY8YwR1wHOTalC2L3nCJIWQrw6QCc7s7x+013GfWWCS5gqyAw3RM7C3mIz
EmOY8saJg4KJJRt5SXBw3m+qE9OA6y+4s8dA9hQBMgSXN3u0M5wOguMwbr4I1h27vhFsI0tQ6E9F
G44AwrChth5r9AI8X5k5spaJJNJSTAQIqXkSqvIRESJOPQ6A3C1hgvF+6waniXHos4qlrnVITgHz
BHQNJxFqvItIa/lqWAXOEvBUCl/9YQlFNT3XRaFxhnl/wIxo7lvTUnUlbHLhDyoxiNING/3zBMer
N3gFmRypbE9k3WhrTyo1KhQSxpWIu1omH7pGXm3zifFdO1DqGPEbUKw1BRPn8bpyXND4YrH2CavK
CLfHadL+zfvldKdF126i/XyCsfX8/VP4G9y9DBSpcrDYUYaWYeF2PFXPSL8fFFub94O430Z2Vj0X
TQgRRs2cKA9jsqOA2eCQqTQ7XCjmE3khsDq/5kF0IFrHY388E1z4Txv6s+hr/k3+69pYm/A5hR45
BQu6qnZEBw9O2Ykkz0/9uHNS/59IbFvfKu9OnJhASa2AKl3o6fuCG2ZuYWLfKUIUmz5gT/tIDbs6
e8jURurCi8wndy3tBvYT6kq02PVfaZxdRlQ9+Pb/Rc0/dpfg7pE0sMIvUrkyXKfUtDWsuk2b+mzD
kRCVnuC9Cm7mDcOKERrSA7oEZ6dlxvTn3ZQQS11/9tv70QAkT4IE2KjbW9USfZkm0jKTFX63dgNl
SxZ46S3h50wjuZvklXOYwdjV3R79SR7LQvOCyTQmtzgb37woHuikZSQ/Ed+4DYOoD7LaJzfrizbz
It5K21DlJOajG5YEOdE/mNJFSQddonzO3CAfVbjnJbmWRungZ+/0GRE35wumGvug9sWIfeifpdh/
d6/M0ow6XLWo6YoqcNARSIJk9AffIlN+tIQ7ElceW3p8DZwAWNMFzwT9tW3wiZT8q4QLRVe+DH6O
MJI8QyNxi3ahbH2fd4PZqbYSfGLmeqcpRlhnWQ8bWKWr8tfYytupjpexJEJ68EbZXT/iZWxukxZe
eUFKR3NIE8ZDjlwQLScOoYf9wyxQTAZiOmvPRHbRhTrDg+EvelFJQAb3s3LOyw2QrX3tZy7TGSZF
uy6u+Yzp+kpj/jtxB+J7MxZ7BrRlVsFG5hbf90RCabk9u/18y6fsh/FtZC4AACT+bwLbi+tWKQep
w9c+uBRL7tCJFiJMVK3VSAG01Se/7SJpJ+K8zVgZ4ot9bU8qw/2kADWOFpmusRDddjJvx8a/CxWh
0Qag0CiqGGtL1ByTnPeLIfMiXSln1tidc0/0B1whcgzZ6PZqApw8sUpccuOX6rT0axxnhCgx/Bj/
XzdJ4b5H22eO2Jy1gfjVarxc4lWG0oBvkx7WDiXesQh8+DuGat/DPWE4rAPfmmJTgfmMoZiIigF5
lGMo85UL3cVJqtq/M9lT4ca1VvjLvUg93yUqNjiQTW7vf/TCaXyWaM1c1K+n+m1+3MvIzkqR1ldO
3L4xIGbEeNEo2XVpVT17c6TGnVGkp+y2S2Iw69luE6IavKCa47oytLK3+Odid/RXcPdy2tvIIt7j
Q0xuqM5KmY5Yo20KA9VkZUvYqNCgEx6u5mtsJHnmAVtTSKnAmYV0zD9C6JQHhfeOWCYCaSv0+o+N
/cif32sbpRfkBQAJCSJEftO5a1lmzak16s2Cvx2hbAYRPa5RlkSFFeaWw3zpQDiIP/Z9giDVmKPw
hFBUNzyFPmFtdvK/hahHWAEsux5WbPUaXlGocSKAfxwwZHaGvZxFUrHo7M0Gf/nl3n+DBrQOVFKf
188ZEN4vo/WYGJhqLddLR1fuj9bC3qLaaOSrzpTb/wSO7PWQgj9GwFL4DiEYJJNL6s3wcbLNnda5
wRJ4P/wQLSPHKHXwGdiFL7eVvhw+v76sJiBDekhQRoKuIMJZS2kjbXFbSBrIclhXuiDwVL5PObsC
FqukTcVfE75y5vTovgCZPs3jz5IGNUTI+rkaj2TbH7gtJOvFHIgyuvjUJdbbgR8Zc6xJrNnYyAqy
vEB9yRo16r0fidiBlIFDWZFW5ftwvkXt4s2/VLtYo7JVpJg5xvAFcpEb4uf3kEJXDEtfpa4nVvDq
tg8CbZFBzJS7X3GX/5ihs+zME1/2ggWYUnLddu8NMM7DqzkGjXjXZlB5T7WECkoG48c6u34XNJqc
14i6cJ8Hc6vcIQX1mHyUp0zLAz/r0o0eIUBoOiAfqdZDkjqjN2G3XuvnnJFz/W4oQYCz7MM5uj+p
AZQcxvhGLBohoigSPwK1v7FDllOARBebuXvpjEMHgc3U58TQZj7xKpHC4UY3DGxvbUALjvilJexr
QgysZ6IWTAt4E1hLe391lAUeVGl3WBweVdGrZMGq46Xtk7UNzO4m1wKT3JGojzcC92JDgxh16a2a
mpCBJbrwWQJT1iLDKTYAjZl8zMCS1z0HiW/+uRYsiV+vawWcdY3jmE9odR2Hz4K9Ir8bte4sXMPC
wGOtET6tWNZvcTxWyU4utJE5WT0yttjk8A6VhWM3UEmZ1PlnjNfereTAtzlnOYAtsfdTzDiiPGih
JEQMWBnPz6IUZ5WA2M0UzGO19IzRHKSfR9WEbfNnhEVyg/gp68IGruo8yDPYMzhmqqnPF3wVNxgZ
tPnePsX6COJo60V4MWw8PRSyxROLlAlMi95f7tpqZi+Dr+nrfMpqGBzvGLDwCHn+xM6hkPl5s/XZ
QEWYknaaxmgKW5Ohxeiuw09klmetXwpUnqJs4Y8Qq/I9qok1hfhpXN2CeCGNQ5HG2X8E22lbC5ic
8prQKonUwq1XbzFZRKFgPZnumIKs5fdFuDB1xrZAlSP8TcEGd9IWO/ntuk0a13HuL45TKrUx0UMA
xQ96I2RzJVa+r8pdBsrhHab8CLPxHDlot9ae/CNYu2MprgkQ7exaqNCV98FeIhwx/qFVjB/9doWf
95DVdVtyWYlFWs+VHb/cWznnFA4Ivw9Er5fmAW2eaMXhs+AugNomao6MuNirtwgBHtigZxtyJQCh
VpcbjvUwgM8hzBNWmN+Ibq5Jtn6StPg49jSgNczcj4Ej4OM5CPIF+Ia1UdYsf1Tv6kl4UcW04qvd
wBygTMAkqWSUBN1AqtmJExGeSYHPSvUE9ET6weUZt79z5K7dI1o9dRFs/fqkXLDFGrRI74YsAYGK
YySH66v31KrrTyWiuesAG7gVZNC0LYuVZJc6x/VHz79ZLq+wB8yS7Ava8m4miwq1zWuOvmO2QNRb
uqFXUrJalB8VJjvdhQb2ZS+6r8eXI7sXZAF3Mh5VAlkPSxyZbd7cKeIZpkjY1F7OBiEQrA9UuIdh
y4/XpgZbQcPBFQ8ApdXUoZtqZmDA7MDJJFZRyWTMMa6lARGzowbtg5xks4aQCJ12jb/IYJS5KWNt
L0kbzr2Mt+wltOKhKVxg5Nujt3dtuZcLbiaMkPNVfns4563nw/1RIXJHpYT9Mce6yBcp6EIZMUOt
hhECYxj2LqJZNBiClrkBXTgtGkxH6jtMqKWAk5OjxVG0EfA7aNUqhHLIz2wgBRMlAgr+r0Z6safS
LqEYq8ZYgpt/SuJmki2N20gF7Y/zmUJ/ys/Z0xRIGqx84toTaH7stqy17Y+iYKVBS/f48YEQqSZJ
8TfqCSqKAktf0PLY1zcjCYqYaW0QfLLd+USaNRVoRDCOBor4IjP3DPGC0sjun/URmFJffmNMjsTY
wLBNTb3jU0mbsOd7mnHp41u8pPCU46b+j9B8dshEjUjNL1Zc6z0a6++6ja30wWB2F/410zbmzKcI
8qH7XAwz8zyKmcT3W5B1SRkNEmuS+xLx8Cm29DQH/azH9C/a629OS2gCT6EH+Lfa5DfRb4r1boJf
RUzYlmGcbnHXLkldpH+SUN+cVvqyunTXYXT7z76PY9Cq+y0dPFRAe6F8zwtIFQQmYDdR2ZgJVm8Z
GXmCPHVqN5OnBZ0mGByAR6R3mf+VHr6UCU0wMaYhgcZoNynwnF9U5dgucWN4ZPfcqE6qQGNahACu
PmMtnOSzT1mUbcwDvH9w+sHpBwQNRYoFgbT/rZwSzzJYfAjhrh8QsFcMkOk3eUV0w2Qo6F6gcFCF
WRNYlrlqqucka43NLUFiCnfihaROEgmKUUASrZgBT7v7Q8aziuWzGUlvLtppZt5oNYmlDNBXeUOz
8T3QWnzVikWP4suFTe60w/WBTP3vFKfSGXEtasej0wy8+q0o5rNhToaEHecRyohwbSl8LIcC6YYy
PWSfizSpcsnzClGSDRO1OrOJpokT+P+Tm3LHuiWC8aFfNpH2UtGTmwCTLUr+GbKcV0Y4dmGlu+UB
KUVXrs5Awb2p4ac3/+8d8c+pSl/5vwtHmCIzAPVItAgKFfPm2aRcySKJ3aVZHpAq3f0UcXTieD9v
SIwmCfF/oFldzBtb6wuPo1Y3y/8XU3Bzq8gpupWwnz6Wik6Yjup0+nK9fjUEKurXCE5NdghrmWRj
zWdfV86qJwoi6R2DZpSBaGdoKi6tJn8nM7J0mIkpF926eltUb2HN/IEbZpmbr6ImklOgUQIY470o
/zh6ucpxDDw8vMSapkBYz5OsNxM5nFkSptTCAS2EDZ8d7aOmsGI7Z5RSqqPZmwtCnq/xFsE+kBNB
RNkzLXCQ2mfjSenpLRx77NNAyCugWeVflxm0Q1RCEEIphPxtA0j+L4jQjP4PD22IetwY2YOnXGgr
fFcK4n04P1bvB5yBXYLWHnODNzfMnyXhute7gxwJeaKpVHdnh8x+UCF0VdNaGP7T+hH8U5urt78d
RBJxKKYGBVyVK9BXFvmPXPtD5eSN1wZ+ylYNeRwCj7iDwNGrAXTcNSZ2dXt8CAqbu9pLyv6Iljbp
K3Bue4K2CFWCJi560C+WS7jVp6ABJpShVCTVZ+xbSoCJOTdUrEiEek+ke1nNu0qIzJr8IMHukJsK
w/OJ4jt2wxbBa0f6sNYnax0+XIl+tcDGPWNHOvGRmrSArnOtDYcYRy9qAm0jykPBI+rtzYn0stVS
pvKeIdFxLWMPKmkz71x+4awSJvvIg3cD85o6O3BIQoV0cnxLISp31q9acsaFXwP8rHH8fbWnZglK
uV97BEAtuJzY7GbYOomPbG06qduu9CiRQkvaU2grsmAU77/QMiwDiZgzDXLevoCEV/PrSfRQ853R
tJrAP76NGp4k8slMC+Ev6xjlkyN0GSMk6w0FGgM2hGnfIwrIhHMSDUryV7ywQ/vmZAhKOcHE61vg
IdkSI4XaRoRwX9geoTi1jlZX0/kt3ql1sUKen6k/SzM7J8rO2uHegj0xG/jVIoKqa/3SLq2tl0nT
DxLiRKmu3Fe0xB2us8TFPQOTYseH4vEGvMgvwOmY3UmzsRA9cViF6Rr2k6ZlXfBEx8woFP02iXp2
LF5uv9mR9xDbNyOEMZJdnuEoi6WHPvFl9OgIA+UxX/vifE94zCB66q44P2u59bgktElWJJ26ZgKO
SxurjISFstXrVEadqsYN2uILLKmuM+d3+9vN+Y2batjB7H2bhdPavgM7AIRINZtf3KW/7Sn84IQp
9XkhxANU74q8USoOGP2HX5XgND1XS0rK/1ASARiALOMKCCfno8iNZF29ZwZlhxREwkSKCzHH2Y0e
Xj4DBk4keCCpeGbh/0+Q6Ia9ETE2wowqMAKpCRitSZ6tVY8ISCDQcQ/mOeH18vghifjdoHN7el5b
2CDo0QWPoZR3LXWpbmjvqdqax1AkW+DnumCMDKmWuqkAZTf65F/oE1pWgSq0ZGcq68Zg2OBc0TB/
cY9k0VR3f1e7u+dTiLslYsPYpEgQzQy5Yh6pUQsXWBju26h2BD8F4IbdFpnT546caLzQVhe5pSNe
XKx9MNXHM38tYjPIo5GyLQyd8x+eu/DkLmiBMUeDFso6muZrWN245aMA2Q+8SzM+miUPLiYXnM96
gSIjWBIFDzhlJi/Dm1NIplG7A3X0hnqDN3aIZSCeNrxZZbYvJcklIhirXHPwAKFtJrO1mrTVxeNq
7A7PHWSbEYsIgsgtoHHURW0wIVYgbzKiJDQVMN7T+nvsvq7gVD30MIpOLfe/gLBFmsesVzoX0TDu
4v3qZsh5EY/IPS/rb+HN7qLSOtqPxeDYgBbB/xH5EFE1sv20bYngmbtB8YAfk3joZdyUF9+bOsmP
eZZUEGTkks96eX+EC0BfmZPGMkKTF6zpBfed2nhk+4iJc2uqJhLse5tCRq9eoM5OycjQyw+4Tbpz
ZnmiK/cvpAhVVIF8fmoiF9mRLSv9nN7YVvrZmiIc8fdGS4vR4S+PIRW7YMqYmPdMZJd+zfBO+8GJ
/Gu7u/YpeNJEaNiD8SpY5zXG5es/AffeVQQUm3EYHn+d2v+mVNf7d8J0MHC6PBUdHTqnE55LG/Ob
4bRcAZx0lOmivn4sfvDy5Ly6UJq/uhclCC9e2XujaFejCVQ56nvtASmBY7zQd1EqZylByjYsbq+o
infD56qP74wN6Yl37oWTgeYzlRioa5C69vNGemiEAyBruf+fpCq1pLfR8qJgz88IbHPlckHis2mB
PbhaQ6+8FDFc9dvLUQ8Qjpm0v14z/5V3lV7bIrMz2Q2LTLtUEOAyD1ekn1duF5mjYmp1pZ9fOfJE
rZYYidndtIbX/mVkPEG9xIiBTlqpL0kfusdB/WK0sU5ZJzy5rVnu8wbO89ThIlfxR9sf9sdiS/nW
UtH9C3svhK+zWi49bX0Mn6xA2ymmG0iH70XTbzl1dWas+4C+fbSXBl04ju9kaXmFuRrrF3UCPRf0
/AWKJ8oE9+qHE95lQQEfvv7U4k5GYuS5y4T6nW6XKqLzDilZUme5zUbKJQ00H9Ye32kBaCMeQj+a
IRMqyfgrl35wgrKmZghvo+Hsv2MwP62DTLzwVJ/hEMj3hWXT5rXY75f0/55lnMSE4vvuyUu/lsHd
4QtEdDoOa8Wq86Ivkqdz++wWJ1Xg0Esd8hH0l0Vz+AL+QnwrYlr6sCMpEmmjvV2O7cBoZ+px/+FR
I91hM7H+0GQX4A2aqYcmdWubEgUxzoNOBAuRPMThzUiXjOF8dsH0kDP8Pls3k47vgZjoSUWReDf8
yApVe9fECyFWQ17lNVDKSItHpy/+dkwWAqX/kCnDOCYEiXs7NS5LYbwQ1KmRK7WzDsMuztE7H1xZ
hnaKN7HqAmX871VYnz8huEm641qMY3D1lBcHPblzEILSsr9U/NGLL3KOnPvVLNcfvkfRQSg3YeUC
fFCf+UiuVVCyPUORDMlHZkPSsxAFcU0V15eWOWRK6/KsfubSaaQbEpFSlwwgMPI/FM6PmIsILDNl
cAtB8cR4dtKoYFAzFuSqq1i+B+UTmpBKN33Wm9yu4x6fLBsRByCfp9a+xZE+hhYUsJOWSoDV6kAu
gfj5xvg+5bjHWy5qz/AforNCZPJSmyzqJJUbCtOPn0wDROxS6UgGfKv24Lc3aj1DYs5fzCf+O6qG
3vGe00WJMRyB7R54YQRkncBT2lfk52kCSZvmXBLkXqBz4mEmuqrsY3Lr9VPb9TY3Fkgmy4DuUh+S
RQAXWGx08gSaChOThzDKxXUDfHTc8Wg6vxcxHVVRWxV2jP9a0BPr+lxn6aKCMLP3mUGM5o/O+46T
esE2I4psewdUbjCuZKKVACuEtdhMX2gqd2cc3LUPDcvKN8U8TXMicBdITS6Wzdq5EYPUHGW86qxU
lqe9ceAMesp/UiFJGOES96VcrHrUE35E0K4dYUfRVXAk7RhpcL8auwhlgBmI0tHsQoGfyg/hXV6N
AQFUIF4hXAs/OSb2hyOwiw+tkrJ0bGl+4zGtN8h31SFCGhwnMvaRGl5VkIGZwa/2SwvTov/c49ee
wchOxsUII2KICK7V/a9wHrKfa7HR9oyHzhNgGGfFvwjf/g1Ma1IRYro+M3S6Tmd1FMHuZZ/eNfgd
0cvZRHZ6GqAWtdUrVBOKKmPX7QxxGbLBJewfBDaIzX74fefaSg6gxjpAJKAMGjsUFVzAXtrY/xFr
wVQWifv2SP8+TQqgjm5TCU0o9NWdqFyFEzhEIu56mPHWbzjHrQPuWr8v9bUMlFyTlGGB9yyj2tb9
9UGGPIym4boCseBi8+H83yuQJ20nLqhrL3/ntjlsKMBMjdZvuztV3D3sD6pa8xstGKtY3kPcFPsH
AFhxzm6pgUKANIEqA5u7fKpKcAAv9rEzWW7w3G4+Q+HS+hH3BQEhH3khbM3zjrpLKWFBzLFFI+yj
YR+vtxzq5Kiee4iPyDcUiOkaiI6uVN9s9ePCZy915RTq8BWtPHnFxrPaBIHur7FkXZM+DPlQjbZ5
UHKwYecEHmbq1dkoUDDNW9O5JVunGA2Fp5bbLTZFKxUWahj0bQke4DH+1UcCIz+cE4eFBEeQLEyn
WGf6S2ANXl+A3+vQJtCEFRpuda0H3ut5WPJffx/xoqohlrqgolL0kcobV2IZpZ0ZvbMVRPmmw871
VA303UPNpQWmylaTDybT5aYZtAqOrdZubZcd3pfA76jrTbKdw63n2h/+3yQJxpwO4e7qIzOffyLv
QYbqkZq3olsA0RrCG/oVtobYSbkotNikYsmTk64tZeHSfw/wvTM6YF++C7q64SjaAuGlsG+C2j47
uCXHezFYahWjKlfjlaPKvEKXFYFQGccSGr6Mm3ZXmQngU/PE6g57g5ZbQk1W4IoiyT0Dury+ADPQ
EmwYbKWBO2GEQYdzDt41JHnJtohSTVuYCEZO25YpmuT1k3iBB8XrMSYQ8U8INelzW6yLcP+54Koa
6PKkt8HdhzOP8M1/q5McdN7JepVGoEC9wMdmKJcvrksi/YQHnXGmWi7fX0fCnDThgndfkHdYZuNF
QlOs80D4kMT/+ArI67e3Dm9tcBAb2lWWYb/CneiJ4OFMeh+jKztkP3DIrWrp8g49aGvdWVQNkabS
Ui43u34hNhz1V6k37FRIPxma/VLbvqmBE7fU0IskTYJ6MUgkpF9R4cm7blRGvvXcihNWe+Czf3PN
0m0w8f5JMP4ii/qXFcBrhoN87f+NjvqlBJye0kLz5QPncAVIrfeig+oAFPayMj/DP9PFSgxiVXwE
QepGG5HiQq3cLGb1BZwZO1mUy18HIB2EsMiBye+fQkHLg4G32iPSdYuA+xzSef0+SkpkkHNPMfET
4S1Ypj2wy0utXw92Xq60ygo9prg5Z8fAUMUVT2DqdfMWcZ3+45Kx3Wp+V1rTUr/dOZQGLWRGUVaT
g3fngOJbdpnaAA1zEx7V24PNvGBvGPiDq2d/UAUen5bPHU1sm3l0/ICfa6gpkpytF39EJJ0KchU0
UG6mkiJTxnG6vDE+QTWwHeuNCF1WsLG+41wqxQ4OgfpD2zKC23d8Ot/UvSb2IEyYj+1h0yamyqaM
RV+r6usa25Y3ye3qJbyLMWbLwQ41zjzvwDRw97ye31TocgArv2YY0M2pNXgFM8DcXfL1Jv7teqe8
zoW7cf+agyanNGBlG0mMeiQQ2GjEWzN3/q6JlCSpldTT/MU/OYEYjC9KxP8LRmKf6i6/HM8xUNbb
Je9QA7mlTHPIFpk/y+JcuYO+/vDAlipxJKL9xsUdTda/yUzBDKIhCaAwKWaoDNGqsG18L/fF8Bc0
oAJhT4JgLgph+H3uZ364kosHYYf86+Ot5EaoxYH/rJpPloDShDuJSTUEojxS1BmLk1X96kc3IXoM
48ezuKntBwnmYyX6YgbLRZGnVAaLtCysJjCLPan59q5M3aPz+d77OXb4rKEoYOLk7QONp968RqEK
EZylwFkSbuXr8e8oLNq5ZzcfkpZ/oupFLBuAYi8XYDZNm2VSizxMhNDWOul8wqWwvYnoEtU23gEZ
Z/wMFH7L9kXHAAc4PvUUNqDHg+S1GLRMZvaTqG4WZ+YGKLB1EYiPwYpX8D2VEB0K2z2drd4vkqAf
flj/uoer0Dei3q7/Gq6Q210iDtF6PxaoFNlXlITerb/IXguQ0Yd567OXb7W+QkTnbQl0YEf4TyoX
i/eoIyVuwRoiydYSrC4O14LL4k4eb6NkXtz5FkDcHowEwzc3u1YWIYVhIeRTg0LKJjE5ZPc9z7D4
2wmgn0v6oXS0P5a0VUMhvEV9OEuYHh1T81A9a8xlzZISHW45x1KbdeU0XI4riZpDwiM3/ad53App
c40oykpvMcuG+vJBOp2BF8MRkHz35bgsNjZ2j4R7S5CcH2DkMkNBLKF/5KPvAHcdHQ+UX76v+RJc
0ukwbxSWdASaBHHn6B3j25UFzf6Tq67PCtRFQ+37jEUcMOAry1xCVn6opGftA85KV/lrFs5YnDC7
8oc4SyfMBXmhtLdSYqciBtWIiUX7PCxqoXOe9zQCEv24zh6EllEzGWh71KkWCYIfzrmTuGW/6OPH
U0vOXp4jA/bF3rYm37HDh+j6/8kEEjKm2foB3ugp+pYLMFk4u8SyIBWgge1sxGfHaWo7Zylcv2Tp
eRRzD6eBJIOmYPKPHSs1v9m9nXocg8gQ/QabKgoy93lh/xKIufyHV4khJHw8N4AuMzuAWmkhqeAJ
xP/fQoatbfmvA3iZC9XCDXYN9gskwmSDY3PF0UWhPl6E25UmKW0pA+wn6XY3u/ffcuQ3unyQ+JGd
yKWHLhUQ9HdAp8ra2xaA2MhbWUDNAQNygRd0aX0SQQtyPjVuOt/KTUQRs/wokNlm9OPVEN3Jqn2E
/oQHNreRvx7rm7Zj77//GlHYn7DDF43DM8+JYQo8cH/iLBLPTQj4W7410MELg8KExHTvzYsmmN52
lbVFsisNmHtaeNfaS3V91kAHpJ2Sx24pGzcRgRhZ5BMYjs11dH4+BtnUERrzSsVl/hqkNJMMKGCW
cjXxIl4sPMwhWBWJKiv19KpG/K14bXjqF3IY0nn4KW1oDGrM3tpHF411JNYr9Cbq3nqGAPxC6lPx
AGYMm9CCH+cKZLlwi8HeyX6dRx2tbKJ9RfJrCaRst6sFp+aaHpY+FuArgkfDk1CPiipuz4yUZExu
eK1WE0Us9YqhsUEWzZ/q7x6Sc+NNCkSJTo/IAtTfDUN1BkSI/3hCE41ByJkjBLT0A+uJGoNaTGWK
L8Y0m8QA/bQd8qyRQeo5JBrvLx/6zWQdKEGEVLP4KhbxVykpHCr6D04qLgURjlSwpbih6wedS8UP
x0cUrM1BzZUWspyDyqYtlCq12gyq2y5NjxtCpxaTk+W0LlgHPf/299n1aMDkH+81OBpxmo+xuh3M
BQwgUjKnK7S1y06taL1rR0b6P2buHTCeddpXv7j59dmpF3m3Do8st0b3aeOvv1PFJ8v0fte2/Jq2
Ox3bpNJskdfie+HFKihOTnNOTmP3IlzpnT5pLWJ7j6ClcvDPYJVtX33cSIdjoOf/4uqBpV3qLvx8
J+SsjXXO9hi6rm9U+XZtBC4kQgyqYVstRChfDYm3/SJ//Bt45fH6iKq2n8+QwCoy8ZAJbNkGFa6h
NPvIzf3xaqSqHYPa7JPIOcET4WGkQ++97GGAjv5Haj/kpx3jC9Ef89S3oQ7WYCoacUGj6O5eJJXC
myImmdAELuaGylsu+GIuxukTLkBiGN/ELQmRajfi6Fjl0CMyr2jGdNQXMJlQS0eBBDDIWqX9UJRT
nZr6Sqw0SE9CcSXLacjSdFJ/mJv76HHo5gon74yZ6vpkWJZei9mdPbdrtWdVWC7tt9RGrRo/Y6Yd
DH/5a0vl22Q0q/dk7Df72Jq3+rfvIg2xqO8y7clPf9b3CDzIE+/p/bLW/apAqd+04LKgIpKXBfWW
ASk8QaLOj1XUc+IGgHl3ylbgbgGdEg44SjNhkxj2DCoIDxrtpyWRPEg9NYMDbZ5xpWceIvu4Od73
0vbvKzPcWsqnVpyxhLrSczTl55Y9j8yBM14BW9fF05+6pjl1HljIOwrd7Km1StmA8rOzxF7/z1Bj
c0A98ck5ErL3t1VQELJ+4nMXk6F1r7/4oJ5bvGoX5Q/yCUB0K4/0I3T1L5j+2VrC5up1wT6v0QL/
CVZsrJBAZ0MWk2F0jzUVs7oUv3GKvtzgLzdVIg7W4un8VCQcZx+iwKZgpbMZpyQT3kPMBQwTwr0a
hgk7lbWJdWeVczQk7YcPriGscDnin6gZF3TdGJ25XJ1Erdstx8DQ+kbD7h8mz8D7whHU+Hxu9seW
/qjd4YHG3dOVLIMcDeQ1ydkAGgDRYwmGjd1SqRIOIVXkhMEW0qUYIRxfq4TWVoOTamvgxJf0bHNY
r+zqmNEncOPwPdgiAHvFLBXjDw+OvSLCt5DopZkcquzTVkijDXz5VI64K2jUaXNJaPLoGhSybKL3
Lpy+xQqWK3GypH/fdyvf0i55evIGTIgwc56XWmgVaTCqC2cqWeJwj5KtxkgwPGmCZA4gA+EkNngh
JvmvHNLcdDr2AnX4++UqMaLpAmW7upKypTEjjshiYdkuQQTKtXUHYnPrtLcDZ+A37DKOBunJVhKk
SfsHLhUe0Kzx9UyrpjNdNe7ASoyhn2LF9QAEFBjjo537+w9Rej8lR2KP+v3PG80o2rA3m8tsbVGo
5zVithINBDDeEBPhb+AXXegkGK6o5UPBLOOfD86JcLyZ0lNHwLCGeb3snyabgRXTH7yo4M3yWRa0
phQ8clFmT7VaLExj36Drno+43hdRK/O1B+LXN1WWl917VdMON8eTywEaejCTXPa8z4GAg/rto7xA
rhTt3qUN451K5v4p7mH3lLKiWTD4mJI+QvgwMPEZU48h++IW9cQY+XtZV7BWNxVJEtyg/UIJo98y
r9sRlproXnKWKcxYJ/jWGCBoNo5OCHVWK6Y/UJ+wnDU47UUIouPYVhNthQmj+mS5NDMcu5/NSH3p
hRHURZ0IPJp3FE5UMh0Al+maBQHocJuIDEelm76WJtMIka3w5k4Z0PR7VV7znf6tzGhxQmrv+TJj
eGhdyhEx6V4yyHY6Wowkr+MyMdQ0ilIdpszOvcJYhRgzt9Q6ZAdVAiD4rOInf2kC2siDO3ZWU0/f
FOI+4+TQ8F9HMj+OPmmORiwczvuTuQ5I5nJBnfK2vTd3X/QVUYxvlZ4n7BH7lw2mrTNfyxMpdvFK
90V8Wgz28ipFCnoG4Q6gn3uusOaAj6R21GB48u486n55f/YRDyda5wN53PY+WFrD7NShWZSNGDkH
cbjI/KGqvKQcat4Obcf7lmxV3DHcM3+h9TTCSuGSyglAftulgWaIOkhkkdwxQNx5KqcQPIvK6n9x
W3RV56HmZywumTtGzrgNPSzNOgB3xwBcn33tYlVpZGYfBJNEHX9zJY/lq2/uIWbz/OMBrBeKC04O
umm0Deia6F8UXtXpOyyThR/6xiTqetmi1zmgvSRjXdqHjeM/4xAXXkGa7b2NiFlY/y69+L8NcDjh
hREQDFFVb4OS2CpALoeopUdJqVbSvmZRFj6JQ4Erfle/G7m947WKgWszBjCFay+YHPrL54c4Kx8p
//Bk5muCYcfuURQOegm9TJPEMeWyVm1hlZ9JEydaRnVc+GIQ/tUDQj3LI3CGAZThg9S2vvfq8X7a
ESwHaWuOALMFXnF49vw8TG8Uxjnahs9Hd/QVTo0BfB6zcgfPjT+rJHtIAUPHhK/TIkzMBZzVBlL+
HABfVhQWqrMbio662jZ75z8L3oRjaKWjbNVbRoWt1V/uUqteiNgp0kKe5IQ/Kd/uN8O3/W1CPMfu
vmrlP3M0MWhnvjoUyMoOkuFkSC210WulJVNcHZDwDoo/wH/dW66y69YGIFB0LIt/ib8KRiuIJrtZ
sH+jg8qWIxJ6LhYRkYs9qjq/IasoZylgzFs/02RMUIqzfFXS8azfwqLgndOA3AGDTbedIRvBlrF9
Pb4itEXbeI+jgOZqQxjl5jblHkQrvTfCE5/f6iy+OCQ1CsIT9MoiJjiRubHH297f2JSCg8eBb3BS
wlk9UtB5mNCnBpUcWm4Ef+PARZZ6JnfsBBM2AoK1Im9hMLPZum+QG7Ukcnwqeq8QhRmr1Bl37wjs
XpQX/LS9eTH37aOrq9mm7Nx3Lsj+fv7orcoP7PtC+XEnV0LBievvM3k6eJ2aDz6dZWgQ19RI1uvr
R6mskRKIEzEAs10Qk+g66jB2wOGE2lW1I/81QUfcvkcdznHdltv6l+CXi4imejOIm/8YrnXIsxyV
KYBNoVgUQZ76GRYtfFcHR7WVQfuV+bEkuuYlJByx0rXrM3YCUop/bVlcsafk4KW8PpFclMAqVQ1a
V/QzWvRgplVYhXun2rgDTrc/GsxG3Q7CNYaopOEKOqlF5HD3kaLvfXToZ8KwlMRExGQtuqHMPI4a
skXwuNnQtog5MSh60lmdR45ZxXOWP1EC0mdQ8oYVpwL/RTeKo/TXIJOWEGEggEvuAV313qaRu59O
vpdpG96WU/DUADA20nLWQxT/eZC5zu7BYxxl6rvtio046QYl9Bw04gCvF5ImW3HMouVngsl24zz4
bmJKG9jPJlk9i8uLAbaevFSnFgP8XVSDW8SWtwGbD4gb3dCo2hBgzpmjskjDhG74Uev7r+juLnvV
YppXquiMp6khJErMn6a3/ZAATYxnRf71TTZ0L2yMWSnnz6IbEPTB+C8richzsLsPO6fzXT/y7QIf
oycCVRl2AIgDS6YGX5bWkHN+TvBDTtiK1N6h7DDdW+dyk6NkNrb80u36MP65rg47sUrnudLbx7tI
thhP1Ty9o063NzLznmyunXuY0hkBFSYt2cVpIXroNmVuiwqOMbWXupkv7H3nDsIovKcxAneZDmIr
a2O2YZR1jwHm/PuhGmDfhNh+RbAObDV9hGJy61F3ihRh+0F2HZe9K7/NwseUDvoJXLhloo6S2weY
fYiPRKNhK99doqdFZIrX0HKQsBH4SXWaQB/DlJhdhHSrgPbTQMz2q5fQ3AqWeOrrAkhnrOwqe7cG
r8OiIEwIY6FhmDI6Ye9R1ITgGrMtcKY6J7PyuTBGrOWACtBUsXmrQQcjCn7xJiwOn8PfkvZ40g+3
vzvGhgNbmWf6rrFg8NtA+kwzDkujSOcIrUgA4SMJoFQhNi8kXLgiMIsIjG0+oMPXYxMf/aWpdgeD
fhpR2XdCSOK6iLFnrbI7tWrRIRWpIPp/dzPErw+M8WKWZ1LaEVYDyFWPRa43iKm79B53eE0R1QLU
M/iCFG+AJ2jEFz30CdLMLKo+xFaxdyHTRz3FDRQsV6Xky5VO8daIRIlOlI3x7jFUfXjqBeoRZKOB
O0VAZ7iyJRLdviQc4CUSC32pR7+i6grEIrGinyesWsoj6ukSGuFDaLsryNuRLLgx9Vkzt6tpVTJN
d/2VmuEsYFv2j2zY34Yh0B2cdtnVWFWrQwM6CTJcrLm6XIkPO4Q3+a3taVSvhbWJ6hkkuZ4bgQsO
1IOImhMT82ngRG+VbUSQSt1EQPrxkHABZ2tuaM+khRddOMk4c84aAiGTM7HJwzrFV4Kd4IvdYA4f
dnolcI4jCfB+WMi3lRq+nWxTb71W6FGQYp+1HAmY414KaxebRvvWph2EiFMP9VG38k7nhQZIf+lF
Nb0dhSDaDmr1xJ22Q0PqFW/sY1Pu5Rgn/+yQdW35IMlwv4gJMtNaSIac14Uiu33WaQYGGbTryCtD
RFy1/UUD6dGiWTe6BstFKotGtY5xnNsFGqffhZmY+tTgUkm+Bhdee/bIUZ3aKirX4eqaAoK4/wZO
VqeUam8mcbNcRFbgyNrbTMz6CTfgNJ+9z2m/VFa5JID1KFWsmjc8j4WzH+QsmKmGZjA7K4m0+fYq
hhvBMR64ay/PX82g5JTJg7hujBi5rVdMNUuFNFvm67hQcJv1vyWppq+hlK/+8J2vs7F/a6Wr+vTb
Ww+nTCD94Ty5MddpANPSMdnZlwruVpRWqShMdpfJW35oLj524DV+iIVd+i2VdPl7IksEMQAOiZkV
h5nJEK43eK5YXbBQQ9AaGSy2M0zEHrb5iDXz9NFichlccaXNdOCp7wxGcevXdvWlXbzTC+fXocZl
t5TKD6t7H5rxupIS9t78Cz8wplNbN0thmASwvxYBj9NO0f73XD8O3Jm7utXVsXjuTLkDqrc6E8Lc
qIDHa/RbJsGChKDrcRq7jEXVMOG4GbGaunTcizdwHywJ/vVGQSsuLoWKqy3PEHBkKPvemeHIV1Rq
Y75X/aXoNBITcGELMosHc2iz5nIEMvcnnZ0/wZMnXGTK2oJ5MGvM39Rr/eXwlALXDtxhxQRKUcR7
fkplF0fVjZWQYOFq0X+R5cmguwoCV2yLfIANfav1qnEC2foL4gh2oq0y+pB9/VxoTdL26n5EEfse
8xnFRwAwK2vHyIsR78s7oj7dzx5zy61uv2bN7Fk0S3VueZPzmQ1/hEjKUbcTgSSgTopftacXnC+B
peIFlzn5Bn0mGidYVC/du2RrpVDNRtPs8HOpZGG9KEPZaRaLqT+DvJzPZ3qqc0OUb8F/ewCe59II
c4RfZfXnv/DmOMajbsJtMplmATpvVR7eh5RqFFdT74fl1FHHgXVV+KVJjDIjOnFCyJR0K6tcpWwZ
rHaoYInEnSaxIVxI/qdP9BJDsIAvkJHnL0nvAOyzJhBDh+R7gFQI68d2tnETyqiYoG96AHTrRVya
AknReyXIcZh1PqnEUrmGgnakmfTZJxdfQHAMdo5fnWObuf8gn0VcAepprOksxvE4kDqD0La9E8LP
PTZPIBq1kelYqH5rFBQ/P83WdyZ5v2HA1mjRottpbYRSP9hI9j1Of5xA3DDwV0DYFHLl8ZNDnGmy
QtE7M6MqQUYBNiRJkkjZMMas7+7fDLf4V6nN4VmM63TrBTb7xuhpLCeagQal1PsskmK5azGT740t
fNhMpQuM5eCepZTTBQAy/ePBk3DJK4Y3WwRKNl17eoCzh9x4hUG1v6L/miZqZ5JGiuQl5k5pYW+j
m0BT6pHByNIgac2VyE0siRvYMYAnt/9ZBFlsLqNkKeKtzDVo6N/wBGhIjZQhEFXBsB9Nj8EpF9rA
VFOlnXyso6e+ghw9NnyebEzKjTVb2EaivKDc/HJN8H6JqGGzWRomZC/bbuDQqkGhHzHkhagFj6MQ
bsd8Ba7Y4QodkYWJhIHwHrmOSv4OQyV/0jlfpYZrdFJMdcQVuRHMC4tV9M9z+E7Z8zC+v5LCWswX
75t9f4w0tHxKuQv4CJrxXw9/Of4Vasmik0iHsyZendTrwekWhQzH7YSPGfUUCBz9P72sScGsZV02
YBTagszbMkmjwmiizvmlFdsFvjukrKiHDhPi51uxfeVgs49t/KVrVdr3TaZTSQN6vFx6ob8HHivJ
eRslJt4rqDHk+GR20JssLh+tQiKJLtIecKrKmAVNoRviD9oHEaYuiFLUCpeBcUSwj6xXMjAQbywj
PcbGDEOdJaWu/T1PwxcvAwNSMuRJ4orbCMTHPoD20oiHMxrjNTci2FmVBo/Di+TNHzmCeqJKhnrg
3aJaoFvYduF53pS1XuWa9lY/+1Y42HI+/uWIVo7++epz4EjlpomSKLoudTMA+4cybcT+XUsMWa1k
UW/J3TvGDjyGdjak0aKGmlVFaT9ObFY9I9z4U20HCmgtZh5PixBWP9u68Znjuji9Gu8U4fTm1yK1
P69b0OvcI8D4Af50GNTWiu9QA/GzaHWm5+eglgoevLpTHolDouC/xP4IFUqz+W0ywN9/4aj2oDPO
HanNaPEMIANJOgDcdHsnZKr0LETWXNv4vz1hcFShbtlYPEV2PYqN60H5gdTkjlo7fpsb3B0xRbNF
WeFVF6FXogsK4xzf4DN7cosD2BejsBOiOtcmmLTmTHbp/UWa1UIzugDfCbFjv8T2ZwOhigel3kJc
DcrN3zfx/RyGcEjv1Spa19cBgcCzASNfUueSqAI2NsLHCIO/rwf0ufDJO0dW1GH71Q5clvXw34C0
osJ9traqrsLPxui6PwEW4FXvcTgU/helEc8TKK3BODe4c5dUvJQf4/ix8HiIK+uoYnqVTchomiw6
A1GDjM7ziT7f8bo0HTdhwZZDWfDfNxb0ZooXwWtGzkpSgF05PTOmqDfEWA3TeMCfyZkR+2Bv9yk/
LW/d/XxuqcizAgwdfSb9c7PndzraRm/vAVaVA4Op4LNGXpLJ5ZQ8D/HfRH6xhSIMJRuw7D/Oiruu
30ekyIdnN275Bc7RqzdqyULYOh6zYGVhtBXKjTt/AJRSs32wVUdjN/BbS3VqCpMOyviemWYKW4EI
h0MPMGOkyroLiY3yBZfM7HUk7gfI6T2AauOS4Wgro/FvMWAqQWw68oW451KTbGKTSMQu5DENY4Gn
G5ujXmOOEODvyeP0T4PhmC3+cbXwH2mC9K3KFv15Be+1WBYSnU2NfUJKOKsp7EeekSN1tjnXcZHy
kg+OtIriARPxezgOEw8vXiXh/w/1Go19oTcAV2vUKWCi04EfNGoPgQwuYCKxjA8lLUpN8Y1habQB
MVO+pSRUbOBLSJttPsiW9HhCI5UmifEsnEJLh5y7teZj0aOMkx+k9sU3W+yQgj1ivra20UQyCEJg
1GHT5LYKQr7Z63WnRKUMsKglQdby8Ba/Tlez1YIzoKX5ViNTd84PXAnPCcNLvZ1m8py6iuxnqlh6
ORRdobsNiFT45i36BTy+j0fXkHDgEPh9S71U8pPFFNX4qDQL5vtQgDLEaloRyO1PLdnsemHv0+kC
BWfHhGiOQkfzDH8nEjMWbri+s5X+ar08MOuIz405h5mIcSEzJoRXz/MzxCOBfxPQTdo2oHZdHmUs
DEB3+4PnjB86VIJNFiP/loT0qMAfMp6OQg4UVqodX0pUEEk5tz6OV9iBFgkIkNVODGZkjHjKcQ7J
LA2SSKxprP5/mAePGnBxkLdRHpO8rF2Vy746EHyfqeejdsQeFJ2anFaZ9Gw4VOcKfwrxj9y8QK3y
gFsj9S935ssr4Ykxpixsqt3WwaeuRHFCIw8BHy2NZDlajh+AxnTGq4mso7m2vymigXtGQ1jjzGZI
nDxXNY/51kEMOdjocRMEgvshDE/dcW+o4tsmOv6UZ3G4Y7a0qbb+JfDw+1qKz2KHGL+98z5TFNyf
cfXRPBnRm3rQX8he2d4/rIBS3shdorGsX99WqFE/9lPkkwUAcct0pH4+Y0TjbYO7ogO3aIMie1yy
KGVWYvkhTgk10M7QdOZ4J9C+Qn+k7WCqeshq6RrB+jZLWQj8HCqmP28ntnY2qc8BlK2UPmxDNXwC
rSf5oe3keoQHJzwiNLvsNAFvsTQuoC4w9ukvs4fa7v4RrV6nnQpw8PvO/oh88XpOz235qnzWc8vv
eZphEtpgvT7HMqX1T7HeCLChTIlnkP/1VCBIViGI+rzvh71z+taoEzjvheAo4seis+aFdLgjYxYH
ZdunSJa8BdXq+urV2ePAB0yeL2XSsz6LlTiaHrBnTMbTgSVss7joCoCQUW7Iq04E62R+hkEIj/lC
Wv/iGiCelX/zdjtm/KfqgVQaI40+7DBNMVbK1HpdJChG/hPf80Wur+MAfKBQ67+WOfrJHfFkS149
fZBlX1qoUCZsrAOPNGOxqhP/mPixVvHucOrphCq/ruZAb1VrofnQO+eMELrTdRXJGmghv0BSyDST
Epr2fZ1cS4ch80qUUBK/miQ/7I83y1UMtGQosMIYbfcwPaR8ssNWYSi38crbzANXFSNbc7jT889b
Uu/tWBfGznT5OdCZ+A+B9DlncFnp/l5blSdFjBqVOjFcJHMkMP/V1Pmt2XDunKuCN190Pel7kXa1
A6VDfZK8ZkYAm/hXqdGUoD4Pk+VDoHAPxukoJG2eTfxvSgMTa02pVNn1zxKUNlBgMZdJjpoH8riS
H7BU8Xi8ZTnUfRy6GpbJ515nC7eu9cEfoeDCgn6AVADacD/2vUeguH+ElN/VFGwzTFUNbZr5MewR
yuQhPvSGy+VfC37Tfpyv5JkJQK7/cMHDe8LBgkBdej5A+8bfYxuMGkLyrAlcLiLK6jF7aq1gaO+/
wged/DxaHqaojTQMjmV1wDuioQwB2PEOSabyVkCoEvUQm7bi4zayoJyBaDsIaP1rh2hbzfjLDZPn
jFMSCdNpoVhKxzsEnX7h4aPPkDD/ng1r9BQpaX+vo7nMRbadOSJw+o7hI9RP6fu6+D7HWRdRHmG2
jDfO0qnCL3Zwpmg4/43H0tWOyuls+aItPY5mGyRQkJ5UE1QUvpliQJBG0zM4ElmPpt+hxDVP2J41
udgR8YDOe61uUApz+HNWaWXHnwb0oIr9OcXJ8N8dcPHmwXIHl3qRbQOvE/zZgQljsofhjeBRUjJo
JT3avhx4BgN/tJ3cBspvM0EEASPLxAPXIUc5BskhKQoW3d6g8rkzJBXwd9fRShGsqhToItKV3da/
iXA7H8Jp0o+WXqYZ88s+OhgKR2Jqlz6IZW8poaXwn0xmofJ5lvvT00xnt2gaUMa1EH9lSa98SEoL
F4Dga7xY9XzojypezuzOxtiPJQ7ne6hsFiwb8mcZWi5vn6eAXcreZfQRz+iArzp1oO3yFSUZ3afI
TnKFARxZ9XfVUHms3JOU8guN3R/rlKKKCPiaK5Lpcb5RZAnmm6E6FhuXXxfAauolJoRFql+NSpup
UwlP7eV447BLU4DlxhWWS9rahUKJZoQ5KPLy5osOgZ0frmw4E6gysU2z4mNsK17+eta6D8t/paDB
yBWgZieU1FeG8ZuYDyuliS+GUcPN4qDJdLeMNIfMi1qYAQSuReUCNV7ud4kVcCLAoZ1+65SHYsI4
tOvHCebWu0Op2AMd74vO1d8pNOlfL07ADv2uUqBU/XtZrlv/IUtx7/r65jIfEHZVbV9HypRG+6yE
H10jsoD5iAYWhwLl5yXleZGJGxpqYes7u2gEgbqy7fEdjpyHAAYThu/sQIWd7VENHGJnb6bLf/5D
9e/h2MxIqapOzPK3UNIUD69WssCDqgen3nA94+ynr0n03NCwl+V05fRRwG0n//wySf/Lm2Ueqngi
K+5lr7VkaqMSCrkrcUwa56Bjm3DArNlK3HO9msvDyRo75xykIC+7v3itIC74qPEqTP5q4dBcG0Pu
Zp0VrqaIyS+wZYJlHr8fNy/fjB05rKTVwhMJKPS4h62OztKS3a2C1KhTmXQomznZe8jWOMthiIrz
w9MPgrFB4YOWKIFieq7QmwO8ogksX/5FCFcEpqtV0ORPq9PU8jGvWk5qHzYd6f8MB1aq8rQ/xkuv
1uILvb3nqpmw6Awtrcgqv7JR1o3L9PX1okbScdbCyBvJVkom9jt6N/FH4bVf3j0V7umxz+Gnc6zU
T6nII+uJCpZIEJVF29Fb6IVFBaMPlAsE5+Ca68u91NJ2iBJshs3uoRoisAs0gK/BJMR0kblOwUmy
3oCXAmoFENS5z7XhGNoAyI2xqSG7Ki1zHJom7mqTV/xhh9qOQtw1BKVlAD50CbCrhHJkHntPIWpL
UbpeFOB2FjhwYHKq9tvDQWTzXN6kAIPo6UdN2TOkqwCTiJ27eRFG+440qNJMwT5vUGmpPvPhNG5V
k5aTm7fNl1DIxrjzrP6Y1E21tA2CL6oV2ubD3LCbFncEYaXdsV2ulONzM+B8Q6B/LOPj5+hA/HGu
qInWszVXkKWmM6uDBxqk3DV5c6FgY1mkb6i8687JuDocx6uNDqfGwDLEsJ4MNe6unnogxElkeRoa
2UdNNLl1xDjIFGWdpLNFFOCOmLU8QfNWhqlaX6+GraHm2SAJ+pNla3UcWwIF5hHmIrEJXk2E4r31
Nlctm5mYzIoK22QgY6RLgx5TNdzpUOz/dItmCII6lwAg+kHnd8MbQcRdV0pa629Resy7cDlMtNZ/
7wPVmtJ6yGSL+eosmzzpkTk9R07hHujpza0NBpMmmJjaom/SJCGLs/Np/PM8Hh84FJFL6fwRVmOm
yv5IV9Op9DyJvqUBGYiCCFGq3qsd2JYL4Wzmdf+NpbnS0DLokLfUKwTlNYEZwDwnrPsxGUoYnqnM
rfzfQVNTF6IoOxcAGvhaZ1Sv82OcTrD8+jImUah473w39gZCOCdXv3U0qKrpZvofxrOPhi1e+hyf
Y2736eKEUMBeQ8MWMDTFXpX+P9cp5h5mBA1v55SqVc5zaGXuaPOjjB/fDm0HqC9Qi8hbSbZjNLdc
MPt7ICLaz5+t5mAzIPph/mFG5FobXn3h7mMiXsWPEYQEx4DURP2GvKPU0oWLQ7HHSTRhOg2EWOSi
6FSAyPujZzHAGCU6/ojcxOdsqcUgYgO1dvvzzZd2ZHnAzm/8byp6pBa4bKN06xeZ9MB6YuQRwqU7
QUIknUo9BFnrHeGZ/wNBlvZJHz6wAFxhN1bz8ZUNvQPZGhjz24f+3as9i/apiQit6smnOzw4aOpj
8MVrBGzi+toiUy1VLmSnggDTN4AAFUYwshJo/Ng0cqDvzJmqLGn8d2O/htrryiCKm2sdbohrdTRo
UmNypeI5ueDSL+2HT2CN29hLnBwaI0Hhq2aI2FxMqhff77qmguhqSupjqaNz/e5gLHLfcar6MC6i
mJL1UXjH9kF9L3JXQm849fRCVaq77gXXyHzy/i5kqhqYo8C2ghdspIT74E4eiU4LiXOCd6peYSo9
2rmgBipVqcXT28ArQaQHi6cUzmjEtQchHLiZwr/VYdWpwCih0s3UmPehbclcrbRUOEe8I9Qu6nUM
vp/rqyffly5KQ8p5NpaFoSlkiBfmXioEAtaE9+4Z1qgjK4sKQoXdpRG7F3oNLToBO7QtAoQpruif
h3wmo49570PomgNxOkIty5bKAjdsWKTdQVTbzHHEBaTLftJ5Fy5O3qPeKSXpFJdx6vMG/wRiw2s+
nWtTgM9qpVHiirxa4J8IeDtX5QVgvXPAYNpuMQyMEvWVi8OwruflWJZYLqpllbjrdQWu+GAYEqbi
5b+31Tk5B3tTRe/uhsk0NvaAPZcTGxPZoS6noPWvC9nWG/5fxoDJCL4OpdRQftNQgrzBWzt+IfOa
gSjJrKRk1gWu8FhfZQ3zR9A0Kz+6cBqk6tHqi2tAmq9Wz4AMYb6j3ZsOhcsOAC46xao/Rs93p6SP
NWeVUsetLfRtiSApSfjIwcsL7xDn9oClEOK0mgHhAjirk8AIIlnv2Ss0JXOs8TnHZ8W678w8moou
LXIhfjK3hgkad8AVbp+8mVFZxpPzY1gypZ97XJzFYH7MdxbRiP/1l9QRJRMRKPczdIyC2X4hhH1Y
yaomgDPr4SQYGtsUqVDLkJPkbQGETpvytzeuqEVt6xinmwZYFXRIjaWGs2ERVx3nKQKJImUNci+w
Zm3QkFIWTTM8OaGgOxGcjLQr1tVI/ru8/BSrRDB1HQICkyWFmXC3LoQl4AcanHngQVg9z+/WB2vu
2kUEzTYMjmAQ3fFCTQyMijxMlIKCAK0SUP3skLkHY9KbBl1QX36OnqShLNKLitaN8SwnTDqWDJ+C
+PeRVEl6j1PbcPPFWOeXRDp315csQE2yohgarvn011skbLpoeVfGExz11LP6Sw4A2pXDQZkKFAyl
0gAkQiA/quGC7Gb/sxfhm8mfGnj8ZaNKX4YvqGQXTj3G9gNkdk8ZGd/VTgmxOCVKvq9r7QEpigFc
ww8w9ENNn1+KWya+XwaF9oBJ2KMhOLTrabi1XC3jJgywYzir6d6jFS3SNSlHBV7j/bj3axEaQXXK
8sVROgdfYaMAit7YJsaujqiKynAU1Qvk8qEAjgF9sb67n2bhFi8TcpIcAldwhj7x//oZAr3CcvQD
uQsTrqGakXuk7QijdyA9OWsybUZmqt+FjW/s5npW3IoxdgBSWoOibVdZ8/sgSCHFzlChIKfjvvqj
yIsZw31ee6VNiJeY87I3nQbcpzHPON3qc6+UhIpwVD8YUIQ079ovyHkXQTrWapPtIXkMZyYo0NFc
bcub3p62hKajv2daJUkMI+6/mB1uLaNynjalOndKNG8vq2xg1A09eplSNx/gyrutKcJ6Ny8PNMQR
G7OXdZFvSWS9Ba6hiz0oddN/LeRh2erHZ4FKfQvLQvl0uhiF908gx+ib5mJ5+IB4axcD8EOB0IZk
bbZTUIEqJDONWybgzx3HMVp7mcko4GybzDnD1DrWYocU4gYNlAy2QlI7jXggBeoT1geQVeOkAYOd
zicRyBhb6BwDs4ozNAnAvjNrtm64FEyEudCD1bDrGk8XUg7bxQPcgNdi3ia0+76O5yUIiua2mhaY
3l/UkOw+GrPvfgWfp1NZrIIhBAIv4f4eJfVzjWQ0VRLZHRj+rloOUCZz2jijYcnzAXXAMQXSw8Ig
wECzTUU+sGQtzArfBKYyichy/QHO2/AvV19uFyAs4CDkW9LVxivLsfximl9QIIKy5rCV583mXIx7
567qDdAMvcZaNZkGXyRIVCba6aaSp5wBn9d1l7Ohd2/cbDtKowegxPN5ekP/UeYvn8rFhNox3Bvx
pVpsPbukwhMjDRSxHgsXB4uGoQzg+XQdpYXeosk+aQLigAdQzL2Oj/Wd/upiep1LwGbHDfOGc7gs
jnSRniDiO8/f0/t9SHZtfhnp0vl4HVWBJKA121pu0pGk4nh8dxaH9tiqGBUnI377zpFY345kHpwI
SWgqlD0f3T069TD1XpFzDt0GoQLH3xsQnH6TBbEsom2XXjZvs3+2+JdqR3zE+IiiJjOG3gUTDQi7
7S4N5x8oJhpP4cAQsVQomM81Lw3OI9cZm5nNx7MHUMncqOp8vf6DjxFBMEjXG9ausGjYBFYm3EqG
SEqSU0totN5+ChPba1UQYWZZHv1dQVHaKzFsQwdl35NJL2H0m7cj0vyVOQWI1Q0YCW+SKGbwslay
yJlm3GQvOXS7cdjnG5Zjy2ExTWqkzjpudjrnOGl75qZJuMPL0H3nAB6+uXLT3yDMZhg6QVWP4m0a
B4kZfi9uU3aHO2LUKI0dEPqr6YEMmxt22m2MP92mSnCcNk4Z24yv5tDyQfrTNr0WyS4AE+K0ZiBm
+mmWxqF5CztJsagRIsITnvVc7azcA59kXVClTHy7OCLduG9j3iLXuarWZIquohELv3LKtcdeSzc6
Za7mT1ap4KcRNJw2GW4d8daJ3aWgFmiipvm+xddhdOpuh2HZ7vgSxNFZS1JQqslLaitH6mPBQUVd
Wd45ljdtSuzJR8Kkrsi0hFfxyzFRfJlMe8ajyRpv/o5UB1P9/95WnRpR7XaoK2rXmJ4zoxSTMPN0
bGvILxXugUA//4are5A7Wvn5tt4nK/S2mKSnYiMgB2u+0j26mjlHEfOYLqexzfvmlSfT5+UHonPH
DhP1InrO2fYoNd6XTpfxHcUJegf29IRKLyre1FkxxKtzRMc+ztVtS+jlmXjIjErNsOD9Iw5Mlttu
KCn0foky913BlQLM+GohZycroArTkLowI9XllCvM36WRz6KayntMsxkdCjNDoyqwmSI9kxD5HhoF
1e3DbsA6htzoe4fFbGO6W0ImASsJPqobfPC81F6UG7mBM1A3Z8bRT3FlDlwwfcmgHyqe19OzO7EG
a7qscp693TzeXnu1jukL4cnYp8iYhLM7en7YAe4B6VR8BVYyCK/bP18Z1vk0y1z8T/TakkGBebkl
irFvl8r4x+8oNFhAbx/chu1pm0F3hT63u0W/BgxG/bRB4jhcj0YZWKkhke65LBpaa8sBMf5vtRrQ
fmjz+MogcAaunKl/sE2vBqTSBRJ9vMvyqovXCZDn0CGS8r+eQSXX4YpoTlqTrsC3+gC9RZnXXlYi
i3GGslf5rH8oHrrIYS6es7rrKUtMwH/Fpyiu+AgLxPzM8AIzA5tDOvtwmlt7AO4+hX204JvhjZf3
tiLmO1it5yeD26VXhw+HuTJWnwcTUPGuaLVZPrtx7Yix8SZypTFeZD+L34ysfrEmz68f5HDeJ4ae
NNfK0q3siCn2FT5PRV1OFEVRzbY1u9GyuX91CRqb1uJUXIOdWD5Na5PHtaj+BY73cihdk2uKMfJ5
6A6WpUlTegu60Izrae+7DcQ4tZ9DtK/2Rx09gvts3SEvfz0YNvzXo/ir4ZgCKPhYSKlPDtEo68qm
9uwWDooHn8HTPQCVLmgIidt/PxIwAy3SQPMdhfCUyQVEwoUoaq0nDqXjFC47F85++ekgiHz0gWJv
P+HAd0HHkB9Kzm7yYPb8hWNVz4N+m5cU8BjCarZ0qpEbXuKokFXMikCROO27VJNgVk6u6FG2z1S0
GQyYEJnpRAuWKo44UUuTQs2eOxk1fmLla0lGBNm0pdvAn8EFetiuyFm6/+u+OM6ToFkUsZ2DaYO+
oz8Vskfbhfle36JHo3i1nJwtTJxwOC9jY/7uex9m8c5iGrlhwNUZXGUaEy9H6M7pGgbrZhg39BxO
ntLFaEhBQ0KCYJBcqo5Q2ohIteusURSheHVYKBy4fhBjLWqufHHDd4cwJ0/RmnX8HD64P8HmzhKm
7XBLxtztI6OokDPTrBN0XGlEuAT+zcKJ8+y4QLsxvVfokhtHxgFjOWPzZMoi5phvuKjY1yb9fSBk
qXM48VgyEcALRT8nRhBxJlH++rn5HeUraG6RjaCPAl73Uo4jZ69PhjceIf+q8bj3FwWR5Fr6Sz9F
Tu+v1foL9poByrWTUSmyo9m/59klczdxNK3Kzgkkblk0KlvxJX0YzLnTZ7YC6Ra9WyNdIHXBtH58
pDHxbXt9MQfQmls30Qnf0psgtZI4JwR4tCDyjvqJiEQunq3r6kXM8XlMtuxLGZtOqxqP6FHdUKz3
OUpQhTY/yB6TdNri0ekU2lf3YH19xX+Jn/JQfzGPRUw3co+SCsB4xRu9TutfrPhp25dqkcUfnetO
m7djptpW95+FzHdA1fHeRl6TVwH0E2rJks8zZ1Ay7P6b+Doqyzj80KNrQA8pJKEronlEkSHaEdDA
Jbq4GASQSTk8TACMzGlWZSXcfMaal7gTe3/ulu/yvXott78LTRZLLvTylxNBMm5+TkQngjiWJkZD
4Todo43zee/ZHPeaEXFe8YNct7M3ECO5XkJ5/0iVkO+dx5xA5k7gdvnCycW3rcZs02KBeyW8+JxP
1yKNDNPQCqt3Bn2gxzuNVEr3n07cTTfbx29lJt9utnUXdE02z5BLdJ047i04l3OLXWMCzlc/ko3j
0uxuPxHBgiKgfAm5H8TCgZ4h1+euPJf3AN7o88RuT2XzUZmmv7tXggg/R/JAWDlgA4TvgTuaVbXC
t552dyjK1GBaTJaTZQ4/CETxVblKK3YQSAemvnnLv6Yq9ucKaaETHxDbhkpqmrgPzWPMoqjpfU7L
gSSNoCvyaOetHilMVOJqaqoYixb1kXifFxuT8gkoO3HBI8BjhqU7XfLBtfAd1PdMKrGZDVkvNoTn
Z7xcfLF4fMhMO7weWm3cxy5XbeKKd0fqpKehkm0+pH3/ABWDB4eoFD8bCvtryMz6cfpofbOChRHM
kBPec3ewUrbmMUBvFyPlNMikZLxCJzTPdHEnis7EsQ3huWvRgbeLYblWPSIB6JE5EZhGCqJIe72Q
Mj4rg+iTpHUIoHBZvWLMRRVrQ7FSCLRY728M+iISZPfHz66+rC9cNeI4FHRQcL+mu05FcaQ/MHFo
MDL0UwCK/JPTmv3amCHkeCVhkViK0giey7JNS1DS2yfQAc81+B6X9/qNA3t2w+sbSuGooKZZCNIy
K1oh/jiRmmYibOQpW6MRvxkMax6bWXOIyDm3HGl1pj+S4b1abvA9BBWy7dGA3AKr7PAaaOoHmdzp
btGM1ULqhopGW+Gruz6Tk5QVmkaS3FpARcHPlgqER99gSW1o33BWYQvTj1or9QKQkTxMRK93TMr2
w5U/xAQAi2DpzFfCwuXWX5YkRI0n/ENnq/TWZZOVOcVuvDAs4+qAHg37/0ib+UoUQgNazjWVJ4Su
rFNZvXuDMDlLrynCYBl68JFG/voKJpZz2DqoU40uTVVoP6xP4un0ZVYemWJjqMtR++bAmiY//Cpf
QNMMDAQsUIPLwue5i/PM/EqwPNBbiELgQLdO+BcexC4VWBXtY63K3zE1gR1MjIS34eTSQm7qnNIN
JaEJU6hd9Py0V5ESfH9jm72txzvEKzRVbMBb8UWE32G9/6bQQYy/5sOHDKGqdzCVpoAWvfK/c5qd
pjen5bUrio0noWaWTMqAnRzp5b6ooYzWKta3UYV8oL2IeOAXLLTvXcW3ikOhfYm4YEOqGLm56gq+
NyoOf2yXa4MI5VTzWq8td6dYfCIYIbN5OkZAY2woboQhmXsXWvNn7ChwVXKv3/T9+GbWmnvaKdqV
K9mnYbWJgo8WH+DkVlM6LHq5lpfmXKxC8cr9iLNYBaaOEJVGtCXA2yztlfILd7SxOaKCZGifkDkJ
GPNk1iaT5n0lRjv1Ey+KeD7UDYrbfDhyHOk9QRRq+sEDObqrei1v22DH1sdnsE+CdtMtbc9PEjvH
POO6nyNpDVvyffTO5tRZCaZ5MCzcy13S92U4exaTmRLxbSFO+CbxdNPCyZbE+8sGD2cP0MTzJt1u
FARU5d9N8Qx4NBuFv4TZqadZ9HU4vcTzwloLhvU1vvLTBZM892JgGAmbb7LHfB9d6uFVmcJ8yqmm
eZkqKmPQcPHdh/kxj382t5e/AbkG4GzWKitmeKCmj1jFgRHJzdAwN2COduLPjkRWstd++XYtm77G
M6+BQg8mKNLpPFuy8JZGvmpMuBTggMylLxmPCMuLS+VdQkxn6IxhcRUvZjB/Cu7+l4Qm4ShJTtuV
NN690vB/zxUPH0NMEBfp0z/gV8ibTtcC/BzsQtG03wFPggNQgZeuSYVrmozbGTGJ8BM4nrfeZG/Z
pBnAn53XuCVodHcY673lTFuwJ8OVy5FLchuvF/WY0qsPcwFC2/CYp/HApdK4mxmVYODpl1Oao7Ja
W+4Mumld4yOXDvAci9g+Zyy1uQssHQWduH7Knt2lALNgnuX7i4GvcJQ5YDiu//H1ONclWaA2q6iw
WZzIBaZdpvI88kBDusLhxjleZQ5l2aejNWdaCOWwTmj9aoM6QNHVhoH9AWt/E/8UIueOyje6LQzQ
A3ECCn7lxNffD3g/sWI3H8Yp8PsFyOz4HoL8c19TAYyE07T42oV3ceotKqLBVUE6tksanNovTAcR
DPox4DUPt+S/MaSfzN31D1xaFYehAxr6NjFemprqHYEMBxAO7DcHn4XgThaovT2HoCINlxwofQe/
KNoUkThdcYFcz6l5oSadv3wH8sJxsUN9Ni5cyXYPW2vCHvjKKYpgiMmdWigzD966F3aSI40CHatH
u27lLPSyRIZ1wBXNQAIiQyhtDyUW+CSK7y3hzqVNzVpOhtp3CtBjAMGD9KsEox/oWqW3qN32Kvx+
c1O3lQafcXeObJe8oNIHIRwgN8o3Pg4BqRqCga/IOufcdib/ndPRA/H/DSDcjlCnCcjKrK2jux5I
fBIYUxbn+khlOBHcYEjUkIVDo3h7h9cj2rk/FeYf2NPpptJ9Y29ocuk3ZCjCEWYLVUrsqFwAAZ1R
5cOAU1T2VFHaUnnYgK44VyYCwscb+R88Vsz+/v6oLrFLiqQVeOpySBf70Rq+baXgk8kb653xmnlk
BGDHprKK7mFj2RcdD6shsqmwIEVXC8WC+d66unenFljVBY1GR7pm/igigQjQalU02GM64gkASKv4
r2l4GkK/OAvh+OlL9KlMDoH2clQqbtZaNrzpOWZmEX6IEfp2sIt9ttCKN2ONdx3SH6N7gEVtHeEC
RGuwXFL7HI2zopomohWxmafMIMH9T2tVBEbl21bTSsMjIgLpuF22n+abVuu1Z3tUOqAD66FZZXwW
ooc5mofXylDzGiWufDWwlcGaM5UVd+C4PF36r5z/gWpcHzeC5rwZ0aG5V2k2d17MuW0RPHOMyB7J
EMfzfPPF+JDM6qa9gSw3KWpQjQWjvBAYCrywjtJYlvWPQZeFcOJaavbwIBySJBfng64HHiJ+Xe6U
c+48pJ+Kn4SUCGC7e031XPf0pJjXjahs1U4quEr/NQR8v6sVzIm+HJBpY4sS4Qkh9qzXJIPpARQb
zugn3fU0+HUWGg1DuMOjit8krxdPkjKsKwv/XZvwv6Hw8MBb7+FJz6FH07PE02nE3gK8Vz5WMIrn
LvZQx1pqwqDcfIRdmW7lXYjOTvGdI5kBkphTvJXg8GWE8lNpuud7DmHWzGN4EgXgMcm64rT6hOyv
sGVzzBYCbzWi78W6u4p9FESRQk6bqOesoc3p/kpeECgVK3U3qThUkzeDzGWs2R8yNX68ZnHwZO6z
9+ABipKPvT1uxGVRBFiW2G7qYufhTwx6uA2yBwAizFxLdCa4dY+uQoEO4aV1TSsdhvU01Cx6gj4B
TI+y4MjvV0ARheAO/W0pLkwuU7QSQyzqButU21U1TzVrz5ntZf2CfV41Yve/NnGGPH3/P6AG0+f2
9HY4LCIwd51SP0x79sZmi20o/k6chU0IPm98NlKJzzpM7IMdWMFSANkLYkMS5Qj0q8dKCWA9JlUm
aYfYCzdwvVvLRS3XkQnd2zdpcGdMb8QP+C4I0XBswT2DWEk1bf0h/4jAodfedUqf8vERMJhxk2FY
sC1sMKgZj47IYMAsu8rMOsb2oTil4U1jDQ/Vrpi5wHQGoHxnjp1P/GKQZG/IZqiJ2o0mrLNeHr4T
8MgrhjSoy4jg8Tfqef9rPl0tgNeo1w/dkHP56DWsbG5F5h18bVB4AbnJRz2FtQcFrg7Uk/ZyKtGh
HQvCazy9VGgrikrY7Gjm/lODu+bEcZpz20ef3IZZhb8Q69RvHPGdkzC5o9nnnh8ucztE2pPnbqC3
chpJlGHTWp0r+LS/t+Z0x65PQkcDuPenC7BCGE2g18pq8mE7mYthrr+04+fDEZFK9Ur5jFyDhwqM
hduQxTDrm0O3hHp0i68RQGnhFSrkzXTnzcGqvWvUI3+fU/eLuIIqExVuG8bKaAaJEvteNDCQOgJj
7Q/ABiMc0pUIb7mv+asnSmJA7+AfoCZj16kcm77cLJsfwxy+Bp24brG+kA0HnwW+J1oJhxvwTgwT
c9EuD1RFXjf1BaixahZREzmFaXQ7XY4GyNFDowZ/tPkK2mF//H5mmZG7q4LCrE+homKpCe11TayI
gEC73i9+wBQQZiw9Xis4aTmSvYN7qGFlqp8WChiOBLo04/LtcnrWJegSjJlGiBxwVdKQ1WHZNs59
G8gsbIYjjpECIBdsyZb5UUg9y5ScK5jSgK+dKlSOGFw13wHc99E9naMzRnODxE8u3Z6e8ByWIPf6
c91Cp2ukNkazIl+Qy9Bgan6PwYTtkIG7c24Q5SW7p87mN79ng/BPlgHGTR2ko1nhLEgJJyCwFHIt
cvwciwB8UIunTEqAdT+H0x+7WHEG19UiKr1lovNySFy9Tp6oYMF7hgVeAh+AqWQTVtxx7pzljUYc
7o7lnjT5dx4rRIu5Hk4rGw9/lH7xDqv4QAPD7S3DmOHOHopxaFxY+qXOYr+7iKNumj8z282LT0fb
07wO/i0yZbIN8B8JNmvxK31pXjsaIddsLcTrsUZav4rHyJYJtqHaYwquMYBgiPzH+6hAfIdAWCNe
KFbVjky7hQpzb+UyGzJYxfYqglqKSJifjZVf4/1e0O9qOlmZ+3r+ZbA1pN3aysH+P8F8Pi78QjHy
8xI/6ttHiHohZfV2L8+1blT7UiyrpNiq6WLuKL+oyDR3JhPJ9QyxH7CbHL+Vsq1ex8FllR78VGIH
ODYOppMBg6ItIl+6oozViV2IIeaLgDB6LpY9z8k2feORqk2QrcSaGmCK9M6mFNRbcGLcwQXaB2bG
9NnPDZXWWDBF3VvdTG2yeAL62bouCklhiD0Yz22b/uyd6NYq6a2dzhO6fynCWz0Zt+SVBgEpbkbD
alEZfh9FMLXON28hUPkoEMqUPTvd6P5Cxm0r5LZPKTVs8BSjDcNKL309X9qpDAaeAPVGvdCAFwgb
AOvZLsziCyRRzHpG3u5Lpm7jnqrD5wfUkldCyS6d1JJXbwCkDWDU6+++UGjWW2xBahMua+bFoCZj
E0zym7k4MMcE29JiapQ7G49NJcTMZ6sAdeE7eY+FG7ffhIW8qJEYRdWRWcbAftubkcQMA2pQs4k/
c2PhhMHo4yuxodmwSTj55mRPVDsSqq0MrLASFn5kJtVhLtnUV37rIlf+rsKc65jTzw7ohKa8QKcj
5cSyvdWGFlB5M8OJncGO7pAD0+VGnEzJEAiF+KBObswr6wueEhlYKe4vsk3V/s2G1U8OX47dRxSN
QEngTR2GPQWJdF7V3NPVMw6YN1648sAS/AKz+ytc14TsGBPNsMUXAPwSpJ3cbWLkLBsgxbbQyfiR
4x+BmFxhYxzxJnxJ6Ce/KTa5demJwICR/mfvFMTLcIqdxmrrqU6NINwN4AkzZJS3c6R64qgQSitp
CCjwbzjYZ8KDbiC/LPjQLV+cYp8jZr/+4CCQxJzMd5u0ZF2IU+FpeTOporOjOXU9ZXF1AR37YCvZ
YWqj63r8pimly+u3c8eLeuJo9aqCDxqyic86XheVMjCCrdw5iM4z7M5hw55FoB2jfE2QwZS0aKot
blREX3CRIeq0Lthx9QzGWfpgyOfmageWON8aSybm45BUv95JoTu2+/32uGV7uenPz2kcysHi/h8T
m3731JQnE2q4QbK1O1VKr0BSMVRdGNKUlpX2Sa6aSxcQx0pOYIBpjBEX2457d/gFsAu+kUsWmRkV
YUgxg93qY7W6Mcn0mNV2CL80dbnjR6X70HfLSOtUQ+NVhS7cZPtOOxPoU2rNhBdfjQVB+B8TONxP
JhPW/O/FQb6xb9MKfSTqCbvyoyrg1Aym4LFGEJ2IoiqkexQjYbOfoG6Awx/gTQk0mHQNXX3qixKI
67pYV5oOd9/sPhOoFJ2CcvOHpu/FVkfGhkfKG6XpxhvVaG+WmUbK0yYxqdp0OtWAEtFlO7aWIYgK
Gwt/fRs1rkOPFkRYVs0daA5d50znQLmLzMN6bzEBukDoe3hopWTJIUqWF9qIx7MMSRJ4bYF91G6s
yM03SWx/XfT2soS+e2Vwl1C2R5R1DT6OxjbFseDOsEIu14gH2lYgA72AnhQ18E4yMOa8B5eI6KJh
gSOJkpSG+bIttqARUccc5cA6jcpRaeYMFR61IoUcUYGTD9hO7QTLTjgAG9JjstwI+grG3dkfUmpH
XN4RBi6++T/dyaW4NvynZv3/76YQn+hpQnoFmfpUn/inqomQQQWkkxnpXqTwUmc8HjHWcZcLmgsp
XKOkYNW8/iFoXYWjKQw2cqBnKC9NhgrFbzZUBU+mpKk6i/arjXuCItsR0glSwkFG3rEIY4KGZOoH
6y/ZyZKbuy/PyoBkH6xodxHC0EmAyjrVqDwaleRE2WzPGgxWonsJttzz1Ghq+SWwOcPJGFYXKn4E
ZdNfoeDpQxq4NgFwxd95LFpm8d4+x8CLZrJNL3AJuuJt/RduniwBE1Hk4rng7fVzVLr9HinT2hDF
PSdM+fQ3YNgi5SkEGtK3smNsll3BsEZOvOgWe14W5By4Vweplb3woztmIyf78y9ZzPB08cD6qdPO
h2i0vRAAkfn2V6qYRwMfMJ2CgqHlHwV3eWwea0jNAg3skilBj2nZdKMWArXSJ0EJkPqrIFylcxxF
H7odf2EN00nz4sjckWLy6QTlH9wBp9xj7QxhIwzTSno4gLHBfs80iH6onOqyI2inzk/npbomPJyd
o+RE+U4JE5h/Bw12kEidQrVlU7pDePjVxnRDKpBeb9CM4EA3U+W6zUo1d8rsinPqwEAUGuY1b/u2
joEanoP/y/lAelCfLOpPGkYrjYIqpFpDwPFQ3FQQtKxaYdEY0C6Dg9/BguS+48wYBkFAg4BywlZ0
sRP/BM5L1xTCoc9ayNE8kEc+9RUx9BwUiSnQZnmnzU9otpK4Fievb7vXztcEqPsbynUCreswr5m3
zo++YzGXGyXscnRKFvPn7KpcBir0YieptOFLyw4bEUqoVZo1HmRixsMJYfMxXS3Tg2jIww0NELSf
s35K/XrJxOaFHFP0uboyBsmwgNA8Px5tVylv8X/VCCfDaGFZX8YEDhcsF4Xk4VtQGAQpy2ANEWnz
pvGkVWZdSNwLb51d0VCqVAxXUJGz563hV49PB4j1K3Ud0g0N0sBusEJZamd/ghYEHZnT+mi7HT8e
Yqn8cSrottHlgC5J8f6LHTlzmBhJeO6rNj+YuFn/yeWVXyY/R1DMYtMIvjcCuUiX592Dg6IHYhXa
TPn3efgRtFYkrL57TkEZSIzpF3ZMxX9dKTOSkH0yQ8+sQnbDtuY04f3Z/0YD/vN6VHuvILPSXaUB
6kLn4sP9ofEfa/p9h0UTo+cRCwnZLeSbIdifqAf67oEQclKjIax+UJxuho4+mo6jBhchwhhnBFIK
/pzMzxARIUX7Qc8mnwbZTEHz1iShT4Ns4rn7rxz34W6+D87VdQa/raPhyUiTCVueQPooVqRjKthZ
KCoa+pfubtaAHJVItd+kqa4i/9VGAKoL7UqkeHlkX4PUhoNdb+nZBBRsMwUjwbtsJS2GV2BbSokb
SwtBOqNrOOI1T1GdK5mdARjIhM/Y9oS9fN/Vm2PZcpnQwkeposBi4kIUphOZItfA1UghPwKrcWUT
UMhReypQlrErxrKy9Y+F9gi13JXywiwvWFJuP38wrpRErZGeJFpBXIxLKHFSqsoBsQX2aYmlItwz
/SqC2D850Sd7u215LgG9tbeWQkLUVyNA9DesjtNUXCu4WkyUNCGE06A3oT8QRkAyfziSImOTGQmY
nCIaI2sgiwlBXcoXP6kMfUiHE48qFxjjSfut9jn2zIexBQrdqB36GgTVAXFxn1RPIU7zfMmCNxde
g/6RGG+o77pVgJD0xApLOW2bIsdNTl9zO0sYW5NaX9arOSlccs1CY4O1Bw1ENz1oXhAvsSecnwmB
J+dbApWNVwc+3801zD9iceP5sPyqOGWjo8yjCl/kJ1ZypHtuxk/tI5hw9XnTp2ztxLBcMZdCkUet
2w5Y0r6FXPZ3FHWIOOaLqDLsnyFkd1NuHgvaHIzczi+BcWofze6gbxs8Ron6V5Yc0JVYwwEc8ECj
l4VOIvNJASUVmgRJQLR89QGKWjiWzJn5EJDAC0i0TrrBvkl8VoxV8qz7yB8Agmhmmhc/Vs+FpAj1
D0ox43yZgjsDLlORTrxjrtFWgdyVLjznZpi+tndmhp+MAAsBkDEJV/FeJF5JziYI0fYpRJkKLQfD
6AMOQ1+GdIJlJP0lO1jww2KkuI32frIu5adR38Gi2kqV9tD9zrb6Ca/qd9CboMFtAhI60ZWd0Jvl
z216cmt7EhaLDPrd6lsV83bCCeP3y0w7gyz9h/Ey2rsOZanU44Jv90H6lJeBlxAFarLdpRIP8nCi
U9nrpsYaUr22Ca0gqrEgxMfKpWZT6TNacbGICqGfCFe9nP6/C8ZPb6B9mQJ1V+pkoEx9oOQeWNJ4
/FI3wccTvN5SOHBCJLvw7dK7yg1vdQuFzvgxcO8i4IuIYZUO4M96BGw5850UGTNS0nU4d1ZEWtjL
Jv7PoXLsdGsA07KCUp3TXM+Kx1tD3vaSC6K1MQcJYzeVoKtxIlFjWcM09EQ0aHgdiIErMXRXkeaf
0vugf4Yp0GhBdmIluUzjQctN3sgGGprHtbWqfy8qQxfptjZtUeNF4+kmtSchx3ADzQgoRRr4Zhbe
Hn7gP6xi4JlGd3Qt6KtdDS6HpNE5m0h33Hlp/avQTk/OtAdkWB2wPmY22vBd0YQjPKO0x6+9Ywb0
E9iWC/UX17haKJI1PQXR5ReWDT7yw3rZDS/yU1569V7olZu0BfBki13zG5JJA/NiAI2uZOLWd5Bw
eWYFjA/q3Ka7AfKTCGEjADpjTqOmmtjZIbF0CJqEC6B7CKg1a+Ou3Dw57LqUdeiM381v7lfNOfFF
+FzAsvH7kV+Ef4sTtP17YEhDrfDnAuEok73hDEYbIRZvV5TJXNWaVmFv2kpYa+nD/tC2m9sOxmeP
sDzADrH83NA/M3z4/mX0VTOIJNWKa2NspUPkOIjKE/qSW6I0aP+oN+1+O8CuzzG9s7zpob6ewFEM
kxOjKpHnFjgW5YJ+klGQKgBE+cFX0w11AR1dNcRuRgHF6qN3WkqqHz/58rvbipuisjQ2OoUoyz2V
K3/wVJ5hHDKeM8uBhxUfQH6PQ67CgaDlyUtMIumMJ5ScWiydrllgO7PPMQChpuVItX4HzFeJQf56
zoCGi87WhoLapB38ZFfIxGvYSxqNcii/WiGO2d0SSvZn18CM+p29wg708AnUaotrDYd/7Rcank9u
13b6CKgy3MwJrbNV12ubscIxMD/Cj730fW6RA5+mqJeHl26B1DkyMPuY7sez7QNuhChiz5YqKch7
kzvuesE81JtQg7dkuA0V1L+bPF9sO2KiOPy+MHnGUxRyPpSrP86oxTm0xdAUnllEB8ixIM32jKbY
vTuDyqh6MSDbHQdaetuGwD1iQ1VxYlwy9t6m1l4jduI8LyRAvFDm2z+OQmSq7m0rg+GfPeYZGjyE
lrmuse5ac0gkyOHUvV/uAdrVIv+53j881O4iYPQZPW4xG4G4vwmtPu+9BDGQ4/Vpt6Q9x9Rn+dPj
VVscBEU4w4V6jehbGf8D3pML0ZDsyz9ggJ0fobXcWLu/XyArLG4RtFSoAMW5EvbnURqZZX8vliip
fdQA3ClIs7RV1InBM8VKvN2zc9YKHW9a9c+yIsMGgejg3LhougjhCABVqB7y3sZg6ThRsaleP9P1
bSrrKstki3uwFjSgcUcUKTGGKI993tKscBuhN2rUlZOsoWiB9kEs7RIxkmubIpPRpANuobbjrKMQ
QySyTSyr5ypulH0aQNRFDz714jLuBON8DNXi71WNjxiVS3lfgrf/XIZq3k8guFZywSy5C4Mp7aDa
weHTM4ht75piFhjylrxN8KN3dflbbXU62PTAP4VioOfsSaoKo8Z5Zta4DsjC9U8QTooPzC/ATc8t
/D7IK25pG72VB5I5SsDUqc8snptp44NuBaVpDuqJlPsJIBFQ/YdJL+AyHEkTF1BO3221Lg3IwYfz
urnJm9Mw1xMHDx76sGDhafaohLw6FyU/m6YpuvMrJFnx5ezEI1eZtaZnprzkrSFwQdWDUjohTm4k
Sldrvey09EeDDKlydySElE/Rb63tGUC4Za+CbMcdNSqGh5kDyM4u3GKCGT+E4snjJh/7ShGkLiNN
B+tWYuwhaNAqymaO6RADGfpQzBK84Me+KI9qfgAqPfHBYN5E2NNvvUEHrsoKip9/TvjffP9mXXbd
IRurIavEY56u1scqtRc3h9ywHthzMEJMUSdK0nbFcLheVzctMTMmoxnIdJD0dGsWOgGDDK1Auz6U
2vCSgtUM+Q/mHEkEj4Ewr0vqO4P4Sm2uHHoy5QNPv6GEa7raHmuyhMuI6OaFupD930pvQJ68d/ah
y0fzJ52cEYqCJmF2oFZ+picdAlD0JTzhEJbyPXvfv8O0XA2eyqPhaPm4j5Jy6+iTt+1Brxnxk7gu
g0SMnuQZ9p2p7t8Kp7GTMq6o2+MIi69CEV2wNAOk0TMw5HoA6i8FO1R42XijyCMQcOHRhaLwkkPV
mgqU8VfCCgXm+LGjQ8MZRvgkYE5We7Fb2/1KqcuBu/wERB8EWhMMY0GNm6CEfxFv3T5KlOAn0COw
UpqifMSKGHRtwVQhdsUUc2fOK/ts1Q1/HppuHVpMQEqUw6t+gZ247ZYPqQRJz2dw99kfoszYDmsk
HWSOUluDqrfhA+Pp4e7x6AA5erAP/t7PlSjFIIj9IPD5Us97Q1EpowbaFUTFWqwqRT2c286ETbWK
/I7FJY1FrHk2x8kGV9xUHpMj7g8/ipU+wdKo6m/Vjjb+LuXMU7ybC6aH0vhojMeLrbrADzmPzp2b
r4I8eF6jmr5AuLwxwCJijMVgft7mQMPNSjoIGQ1DQKmVD4pfXcvsGB6b+Do3tqw1YUMmBUW8vYTz
ohNpAzXkxulrd++0s8QRK/L3Uy57vD+ArNrplOrRYOdLkjX3L2bkA5G2fVzC//43DIeqpNsJCDQk
cg6alAGglHKcmlHWUv0ZVMQ7YdajRKCUOsoRqQaA4W8MNT62GF64MXbgcosj2yFH84vk5scVGy+F
+78y0bFcDd1MP+/5pF8NnGOL0f6TMZurmz+82SeznkR3vFige23s1mI33C9gNAQa7R2uYR/+FZH2
eq4zpP0mpkQ6pgY70ubv88WoSpS9+wfJ8SokO9kD2iPk+VB1PuREqislpuYz57XouCegy/ZfHQ97
QzWs+CHLEJuDfgwoEgXeg4ApiS1/x9uNuxWmu0HCHSmt7YtPNfBC73JmM+vj1PawMF0oblCeFnuA
+pspzpUxBnvIt7OK/yPWTcO4GPglEMwyrnazSIo/LRx9LwmxTGYhuxT/hHoJJJ2SjnaYMdt4OYxA
IxwWFk7MysS1Yv697yrqQBGIQ4izKoaO2g3lQ4/TnM7qdlkQ4P0M5rd95GuHyF6Ses3RF4uR5WBH
FruUXW6UEoIVU4Z2qzlrIZ541mBbfk3tm0iYmAV7rdPcIKaDZgGokyL/YaAMURTvlRGRRL0Axx0L
ZpZG5gUNUpr9xc3U+hgER6K12QKII/TA6az5k5lcSgs8eMsCzeZixOeMOh1l/bFUC6QbJa8joUb7
+5ExmFl0FkZweHne/2Fx6gU3P18pJo78ZLvtuRgAykwHMsG3Co1ymSEKWrkKm3/r+ZavQGEqTCFI
kR5zzJZKMS6c0vGgPsvdA8bP+ZgB8ZxuSH4QcRFaE0ijoBCVCJTaEzTGAtwBbVepTQJni8oeL+6W
Dz7pc60o/fkcs/9V6Z0cUSiFgGz4v89xPsCMBN/hgbX9jHs7J80dhOIIOOA3AXW0kDB5LIDQa4fY
zjhh6JgWIsvYOf0PntuBIsyqoTgrCcFFDpoPJ/KgZB4M8P2wI08wm2g2+GKMcpWwBh7g5nZ/ZNCI
mc8c5/mrK9384XhviUY2bf4/yA+Qgr+gfv7DaXtPsvoO1wgKC3F2h8jO/35n35tOmIfTmwYn6ezr
N9QZLIxl6ditJYj3wtg0ODracinV/XjJPsRL/8oMuHevs8yVHc5V67BA5hIvNEUQav/6ydD/0b4I
9+3BQSyRrWp18rpjNAT6QbiaThAgihO2QvUNHxs4NgsOrv2j+50g/sLp9yy8IuvQCG2M4ipOoHXx
hdpjtDu/U9JyTIZ+IoCkZsfzHI1U6CuJ0s6fyhcxFlyaRNnLXxoVWn77q6Xk52HlCMBT1ntN+BZM
mv4C8F5JWQYmiTSZT5lR9oxPuMY1Zb+3hD4QzVFypOOfjar6dLWTPBhnp80RdE97P8gujDdk5tSH
0UXM0GYOZgmJdX9svDwnsdrxyaVz0XNwYPn0vqXtDfIEp4UKp1CAvkILQk7FSdVO++0wiWzt2Abo
lk/Tiev5EsAmdX2cdk6P4W7I9TG5jsb4ACMrPe2MTxOa1Prd0mIegiDrWBdANklna8nTZGtfO2gA
MWtvW0WR7wx9KC6qLWw7pDv8VDn9aBYBaz+7HuvCFXLGECa7djP3Gk8aAId9YqZhUcfzUPi8RDKv
dwOOYfteamnfdQJsQPntEpLsrQqj/duaNN9aLGJuJGRk812Mh0wnVarD0oOAVUusXOwVob5elEr0
aCS3QcyJ4WKXZDWRC6u5BDWHkmWlyPXf+cBgZWLffOa5mjLVlUnbqkysTs7VuSQ5ThbJ2vIYcwK+
3xoy9yLGNmqUyX6cc0lq7v5hIXxg9gYPedQIiaVkrc4zKhmurAAxdGG/5zF5eQHnaZyVvkQks4wK
fLt0ebIq3xhMpm1EUNJJ0/tKZWlwPsE572UwDUmdMjWqDqGqfvZGnVNPmahSE9JBF+6k40yAY/7e
AN1gvL/I0a9KfEI1/ofM8cWRBKj0jtegHM5b8VcieA7PaU6PXvAyUjKcqfkls5SNEZWyj8Kdt/cg
lNXgUiCpTGD7Kw/PN9YCMTZICcQooMW0MAMu+ndSgbZay8q4BLndFFYV7qUEWtjLhaeAIKg50zKo
mZ74HcAzWvrPuGTjfNfiQR6Yffg2L99iFWfWmhmnArJJZXhcBrVIRIam8hPmSdd4Y14bIB+YwNKO
Z19UWJpw43SdE96inMGnHvb9CBywPhF6hN5dqZHOgvxOHnjqnR6Mo5fy2NHa6LxgRlAC/U01VLmX
Pl9BwOu2wFr7qzxnmFF+ml/KRDYbylHTEwAbpiBwGNh30pYLQCDVtFcKCUB06H0pm/egkQmbMk/H
s1iazl5nuwuV8lRUmZO2JR1pOK95SIbLoypvos8BF7J8HbQCRel3pt6Zr3P7aPVjnQsTAk5HM/Co
rDqqPCtM5grm0s70xejPG+bt3yPgsAqQLIMAlTL01irtFO8I3tXOyGMM9esA8kJQ/lCAJl9eq4Gm
rxNfwjnGwe7YMYS0CeRHUNotBMNcSess9nh1XXUQMVq/Vx5Jnc4mbHsxwcY1A+FFv0zktJ9DeJd8
fhzM+ue/31ER3SepySEekhy+JrwooZBCQYkV9YPtfvzVKOS0KIHdB1mSysNarV0C/m4P4NAa4ZwS
HtS4yPaWlEHCasF6UOv99B+XE9kZww5yrvxEIToHpXMDBwz6mP7kyEkl0zusZwnibIo6EHJ8BkJ8
21H/LgHwu1pL8jgX+byUuMQ9B58JIQ93oIDy+IbDFB63M7c5xjes4kqFuynuP0Psumwn0LtzmgiY
km8ZLDTniUPD39OWcVhDy1oWg36aeO4ftcrvqIePG6VtDggkn/zExBRMycwvHpnk7BHROSdg3AyR
zYPhD18vLCTzB98MYSrOZht8e0n4xXtDBxS2C3waM4A5aFgQXRjo3ZgfXoSnwV0thIhMwRd8ncLP
NAU8GHwwxBqxZImsQfbJqaTvzWmteup/54VfcToqLfS8GIGcRdUBFI0PK/fg0lhnN6LJtc6Dt88R
PlxKNwHOaq3FhWUlO7E2bsaEn/S4Ge/CTzE47OCP3rNNeIQL6LKjaiu8Z7cI5i9NR3e19OC5LfTa
lTYWiq3FUsbpcQPsTpH2wsWxk4vra7Nm9KPdcGZSkTY4JPE1bE9r/DOWS0aO9xtvUUoHQYdODzj8
E8eec39UP0Xy8okgvldlDl5luOAaCIAje1j1B6DSifJA1rlxtTOXgjkIrJL71YZYgmKAVedKCSFe
tK7xHLmG6elEnfcm80YxNjrE/Yu/IT2uI6+9eQCYfXzF6QL4aCRC3y5/9TqsKfpyoSovzjlCg70E
hfkRmxYSWHBM6DuFGS9NjhN4FLGjLA1kWdXcMKPILiZquFE4rvrtqLhYcm89tI5Pv4kBjm75pqyX
qB8bplPriNcAznAanzoOHkctuBqr6jCDKLUoU6TqedQMD4zPKA5E+TJHzuGrdKp0AuiD1Zfl63SJ
AM8h66tAuxr5H7IdeYYfDXQD/yA7JEKCWRrdiNUTtbx1UE3JEE1/SoPpwaIz6xy1iY8DWTLEF0FK
VSjeQARNGCms3YiRKiidvfwF5gWyExFn5jCqcUF0SE3XMrFi6yVoJXb/mQF8HVOS8Fs9endQLMsK
WIHsJNfg1CFD0fLa9z4KVXP40R+eg95RBOtFqvydQ5ACBLJE27tMw41sU3OIgg01l7+4LlE4k/NJ
pQUEksuPDrN9g2Ftt2e7I4oEat917D/A8WZlRqzpIZ5DFn63jwzM8ZbjQr/RQRLAMKqP73NpXi2/
6DpbsoLlCEpWfOz3wg0UELwmEeYr84CMVN6k0u4ZMUF9cU/9ZhzP90XrJ4Q8VZqHWw2sBcjRrzem
5nYxOUqv4uE3yvmnvDebiZ7hcE8SYGFRtRLxtqA5Kc8XOJGe1Ds2xcIQ3YZgseP5qhPanrJ/SUxN
3GARGpwCgHf4MavFQirs/aiFGvZJJK4SIb8GUE+wi0jDgjjdT8rxhwHdRIBJaDg2TcfCjxXOGeJO
SdsraPYDR0X6P6u2ztnNXZx6B7xUKJtA+biYTSga4uYlpmnCZlZK+0+XtjBQWDWFA8CQwYhGtMaF
4zpOSM4OwM5DeigUoQrE50wYneDGUTMPxwAG4bcBi3tSaksMTrKy5qSJXqwqPYG4dTJSGwmYTi1m
u7+9U5fC+wpMe5imVz8AMOpc4IdtNWoKs86PpD86MSVclRhG/xeXze/3JIo4OvWuk5xoB4Ltt5bW
U+ggDWkH3nEQomFjJUWTg7zE3F4ylaFgS9FhczIS+QWDM9fB+7htt4wBSOsdCeDdTV4wTOQqELHc
322QlIeQPhASrNyJW8UtKWzhju5KvSXHANFp7AjxmwDN+PBnDS3/TzEn+/TjsR3oS4bcWunTlGY0
DMJ+/3DlZ+PLw+GUmCgsDgXzmuvfQabUoh7Sx2yEIici3ySCPrM+O0+r8mblGanwzLw3sQGqM5Jd
c/GemrXyOXoYEZqeUr8fEtdq3BxzHvj6PriPsPYNH6IOtHgC+I0MbcwyITeAQ8SXgZaRmOLPjs5n
GLf0Z4Xi57EEHqjhQ3GXLUT8R5lYohZSutUjgbesLrI91CR2yMtUaP67q6MrEzcLDpQD25GYOLE6
FGoC3fZg3CzKI5N5tMV2NFJMU+sWIsqrxULqG0TGS26IDjx7+hfl9IqYrPnF9dGxLc0QQmFztWeA
IlY+ttf8fT6nKQtinczdgIs+kKcrzy2H1X29dcOseBsYN/Xv7GTrkWjMuDYcTEGYHx6YSG7YPSrM
sXBpIKDvp94OrajJtSxvPB0YvxQYdUyGkNB+pX/yKx/+ObTiYrac21N/XSXKn3PGjdOlOi3AARd5
43i8kN1FloRecdIHLAOk4pI/Tegbcwa+s+Zydcfyt39JjDKK7EqbRBfqNpp3BRGywVQVDXUvMrQj
TWg9lQlA6Fif/YmyquI+PreAZBYC7Wly6WqN26v8+ByVOiTlKMhUdhQqygRrf8M1aaezullTzQpQ
o9MQdCfjOsvUfUOp3bFQpzMSRmH5fKdExNgRw2S2HPLzLkH8kpPAv+8nXk84XylVpDZePjVjJrpV
OurHYY9ghsP6jHuVE0hVQO7RfvRgVtWVZvKfdpSJ6vJAqulo32VksH9sMuTd0pKb/Q2bb3Oq9e9b
+oSaWTqPW9ovavNG35O8Kah44l0VPMyw47f3NAqvH5kj/rr2DeoKbI419qBRF5HnUmMabPlyikIt
Z0xNxSHdmhdEQ7scJBjz7QukUGwtHC7jK2ka6QIot6zyd/JA/XCXqxIAW9qW7vBDb9LNtZ4GuHhE
aJe3++YQ8jR2PACkONgk0IkopBTm0i0m4MsoRX59m2AQq3edNJWna8zT1YDJaJlbGOkHsSZahhUU
RkfbKdAyUM2uAKNWKYY6vsPXI5/qGTE/Jeve4JI8mm2FE3aok6bSVG3yaDKWlVzGEYvI8WjRrYql
6nVyARRPAxHuGGJQ6JpPJbJqZrlBUEkg2GsiAzaxwEHl4DvfYIVBKIIP6v6Qp1+n7Ye+XbRyrfEM
O3LYdYUcY9rkerN1y5Wp/6guR0DoEhPL8DgpkparqWNhCnzDFY1IejzemUIMTb/AwIqnsvBm3z0R
1vgTacBW2zvBuFSiDTXnvhCVYhXkpQRGTRN7EOfJBO+1Djnsa+DXJlE6hD4l8P8PoGVHCO27LpnW
/iOU5gOArO8OckP5IQP2C+HMfxPkrBRUFPTaRQ4ESu14AG6veYm4V+KddvLb0i5v+uP1H747bOkH
8g65eirYNMVswhWH/gJVhNl7Px7XEwsjy510DW2mIqA/4O4F6eHkwp4Wvmh5WuqkErIaHZ3+TfKg
lOQHHLKpiQKa2n2AqlEpqGP07UvyZIAGtZy6+tGyDUF/mfrNnj+eMqnzp5EBZoMaG6L5YhtVIYl7
u+GZh0nhyxkdVHcZ/Oz5/8WtX+vfSKWQgn5Zx3MwvNlrE7l9ZyT8BuBMf96f0205n35u+sxDPIsl
ZKAjr0PLZjkVcDhqgjcT/6KeutYpA6kEAGCgi09FOyjylHemQ/WWIP/sgrHQHYtz4owejHkpCXXh
1tQhHy2WQ3nSD3m700nhw2gmKLEWOdxsBFVoAB1H/4R+chsBPuCVDEEjKWPAVmRBNrXnN0zrxj2O
HZO3n0+07jfOp5dq3WBRQVBOOohEYgyVzP3XatyzsHvJhQiTS3WOHELboae4VPVj3z3XBxCQ6dRI
c3juyZkzEP4MFWN+1oTq03wK8OEnh11DGRu7F9fqGB0uL9BxWRc/QV2YDlyGHHPUpmrTxflHwe0+
+sOsuxgdgeUa85UChm1k5w3yIADmClvoQ57tvPYe5UkxNv+ruU70YLc1GcIZ8eo9aMgIB7aZvN6i
/wab+QmsRHM5rHB/uaygH/7cVHId2YuKKEonw68Y9FjAOCd+Cj8NTMZ3sFP9mXORH/r/P3NFw1Rv
cX/90M4SAA+JY0xip21KHm2aLuPil1c3wDU95WkE3sJY2HABUpPZG7F3E+vhpsEMNIcNR3WwT2ae
jHUTXTmcuJxxkyCJlaTY9yJ1CHdb374SkxVX61QHp48sawdn4fGnF5jB39st6s2b6G/JGE2TvQFJ
MMsdGM7O17MHpDnsTT3+25OcJCQHzuCFxXm8zldYULbsorg2n0zrf6ad+l5OOMFjjKD75Qy6qAhg
xwypBMOLZT6wpqEtncDH5PyDrJp8xBXQbf8igpvk9ummsv2HEZrXcu5o+qpI0WTQSqQxSltfJ44r
Mcptr2JC72N8A/T7J0SRqGh8mgj/tZjRAJwlMWFhkVluR3eK/4wzymI3BKMUw20IyYpzU9oNCqZA
iB0gzkUYs3NiH5As9qxIW4+sfaAjjgNaoqxakJL0G/YTVr4WVOd0WbmzXifI5DoZgNh+clEkhEFd
mfZG9yKQiz+p/BSjhwNt039fzfJBZejGPQE01NTfubC6uddWMWFLOXiPHXi68bPt3esXWB6DcyBb
dQ6al26VEvKnhZhzD/jFjLK+y39z8+qXeH9ms2EvBxo7PpMFtCRVy+IhNKIjYVJv1j1PWCZekBPk
iKz7EQfENriqFlwzDvOcaNaX5tZOA0ccArx8qRn8ZyJLqqXUxtUKDLzK4voabBlC57kaZJaAf3Gc
SwpfLBgATCnOpSpefmMNwLsG85ix9w8TaQmKLoO30lT4JOdKa5esJO3MyjtKD+3p9z5T9GUhImkD
/5+0BdU7NlIbEeyRhA26xt3rPqAOemA0lgInTQrcxoqrvKGnfig9T9qmad55jMo4/3sa2wqkqn0B
Hrp0JZBPc9N6LChIY9C3hjF+m1wPKkU7OaV0qW/ZyExhYHvf5+BBMY/qFoF4B7114nRJ6rLVsvbV
IDdleOi21IrXIsoLKxmj13/zJd6zPGtnYNtrIJ7BvT7uqj5HykXR2MdC8CEmqJp0Eti1VXL/JwIl
nanchbJWiNiJVL1RVlQf/1L31hENBxkiPU2z8DeO9j24kbCz6zmqMZR4mxQey9PBHtrH/2ZaC3EE
hPLYQP2rcv2nJ3H/O8VdchGPqRPHGDUt1taiXdCafuY5wzrKUt6FAc5gqgeRcFuuhg81UV4ch8US
LU/nDS/ci++OhDm+PJVXtvEL2nUJjB0Efc8XFLLwvFyQV9l9opIxyRTuy05q+6GFVoj/TgpuYNIl
Wq7bfFyF+MOUJ5OsGsIflnQzS1A+2gDQA+GLpk4hAl/vSLHuKwfMu+L7Ce3JAeASzxMBVjhxvrJE
tpft5oj1jyI+BMi7WuY0g4zMJvW8Tnpvexw8uinKeWYndyvPNKrA5ArxUz++N0TYi9AjBsMoMan0
xLQsKasYIgUE0anTLTruGoboSUQ77igAymkhjA4kuXkcH4xEmF79kISDnUn/3UqZ1trBjB0ohND+
T8ZMQ7Kivk/k/3pfRcMRox+ZJvIkm1AfjY8fs/07hiBdEsf56hL2iZRNgDnnz9nPdjeCfeCFHavh
mE37LqyNRcMbDwvXt7Fn/xJTX+IgUIplkKLeXLk4RW6UIsrTq9RONmmxi+ZBTVr0Ho+KbE0M9Bh2
QkQLTci9MHwC1EKz4ETSB/aulAa7bmxlCkMBvnyByCPmcf0L9V1xLf2zcK/Lwj3zvhwYKR/U+uB3
EThAsjEEe9jZHTVr8LFquJUTn4SWEsqbdv5ODvpU14VKX7BX/ODO+C8dfNT7lMLH8jFFL7/7Ggk0
z62JVNSveSPQSd9Nn/i4nGn3d8DhqnBW4DC1vlL6lzUqy2Ax/kqPui/765hv/akRhgef0oj4QUmR
v+d/7grx3HlymMrxPNQDrEGW0BrWwj3Q13DqVbt9duw1W+yjRvOXHmT07K5Fhg7FfLPQUkU6rt2Y
CEk3H7j7P9EnJ5P9cQVdKZzd1VxkzmEIlB0+s0XIBjPrVDJymau+SJnTB9BzaWoXmaFWM/YIVZJI
u9i/NtFdndySSScekhkizxJlyuDqd8D34C0ZJSYoev4q4nfT58FyQKO7/br5zDu/fA+yjzKirbL7
IPD8Ad2Fw6bBRe5k0wJNFo+wYyOv2eaR1XS3SjtdTBCbHypBNb1NZSO6b7YhLAV5TzzmvUkLn2Zi
TwkgNH/nW7UdF5Czzm0gSFVywaIPYKn2e8EcIfqofPcp6cUWVmxyFrBw47McKb8TT2x5R5DzX54b
aPuLG9LkoZZhc/KmXy7RJoCjOOJMJgGW/GQ3ZdQ6blW3+wrX3Rtd0+x1n3jWm070FRARxyWJG6DB
0jbimf4z3NBLpOd0HNPWEfQuxYOay916DR+nZ4hX1zI0AOEu2nT3MsaffLiKIDe48Obxqn5qWkLj
bqWgRnJ7llojFNO5qekB5ROlZypyho5GWlmfRVhSS29tPima/xbDHz4oJuTGKPmthBnpJxcYN9+P
w3KKlivP/ms7SMLKj+fE7cFzwahRbAlfsBmwNCBmCD2+EE/e4TYHG/7CL6GpYx2ACM5K9cMImzxQ
gF2Fao+tTN+/I6kP6kkqUJW3fav2gTJSYXQTod3Z692LCAqdNaK1F40ozTp0qtjnbI/T6dpssprq
cBYDQgf8asdXKhqRTs4eWuaY6m5ZnWpJuVSuRDuC1gD0JQJRx5EYF+WQUsyy/VrzF46ZycgiWp/i
I3RAVrVpLjPQ46eow752kpFbQBqjrBWT89mrw0AfQugwm7epaCiAduxppUydbP+j3zITBV25+oVu
8Ps0MGpKd8/q5XIR1l8XaInTWGDXivSXktSZKwkXR6txv9yyE9T1eGARI/douGUYBfysNbqQgnei
9ZST9X9K07dqmNukLlw01UEPZ55omR1kxyO2jaOinqcqt0A+WIHzGLlTG1R9RTtjTIkewTAd4OZg
iH1XFDVSMPqN18vMCJhLMyPVUi9mvJOawvilyNLRAJl6ojb3qR2Dv0JWox5ST3rMN4xT42PtrMQL
SNetY1juYDaunYzogYrXTHsTjbnEcfg6FjLFq45Gd6kNxrXwXUqa2n/cSQ82HBVXNA5MTKwjbYBX
FqSjqcILXGjqXplrmI8X1tsf8UaUwpLZcSmWdTBC3QeqtEYRQslnVvNUl3IwGH4eA108Ux0wiwDi
rV623DuQU1W49ABLOYYUF0Q6EN4/MNcd0Ph6c2GnY9Ep/dTo37oh68+3bNSK3u15DCM5pxqOT+kW
oGkxPleQA2KkwCXE1vjRo1LN0cn8syyk/IzmosvAI2eZySqEJUH+Aer5IVUCmVQ5CjfRwCi3Hx5t
d302H49Qz7m9Dja74dJnWX62wqvT/Bh1cwewuosjwYnYfGoKI+ktAJrZr1SOdzQfAwr8sVJNnawR
UbDeFdWy6ZcQjzudHWRD+7ueK2ZUNcc1+KdyxmRpcZtxFgOtuw/L0pC6u+A5CUj3DzR6IIWSuiLU
CiLviIJmzt3mxWkkrCBjdZ2yRbE0Nrp2X/8NZPumkLXWFPyfvKCb+gVg7B0iB9YalA08S9RGFy62
WRHkiwcIFYnb+Zc+eCcUsK9UmR88E0ftSqOMYSdy7iaDYyWEBPv8YXs+CIsxL1HusQByin28eENy
inYKS1m+Kq7GTPRiLCMyM9gGc/tLksQmtxndXElbhOWOIeFj5iXGF5lNYqBiP25rLqjLjGal9rvX
M7jxHNPa8K/ACUxd8H9CP3M/71t9DwVZuTnA9gpkLSrldsMA5xwCGOsg6I+hC4TxkplqCLqP5AST
lcAADx6yseP6zIFu7zrvBIqQTj4RO6Db6t5900N3kvxqHBKt9xzBznHQ9vpYxly0dUF9WnBvEE52
4tL58VqqkzXYWKiOdre0yvCWndD2AEY/DxiIWwmzeJKhmY4fELlYx7JbFzzmdkZgtmnhqxuFYLOF
K71Q2ajoOZd2eM0XUQKuko9AXmNWKxWkZRMywZEnK9X32fVnp6sUy7hu/AEXu1zbN2zWTsCDh8Eg
b8nXrS6w8OHvRDCqjo4G/zJN54y9mRwvBeRe86Mlz+9tdcPzfvvN+xguC0Cpxpkf4grXWwTVHtNV
8CSANq+56INxDYJDOGT9cfNCQpyKyt5ATBATh2GvuGb7yBBMCpD0RMXOoIJvVIrtg5x2qLofOl/U
NWJ9GuQV1167bvs2MuMOlQATc7KoGtcYtBeiRdZee9Cm0+kjjWBVerRw5/dICAuewB19S1whlToU
1gCqTlBH1MR6JVxVV1u5Fs7V8KXIYX2F9ReyzSbNp4erb+j2JEZffZWNTrjZSFzd/XFY5w9X3wc8
RqwHKXYYyHOr5WEyCSrk2S5dwJZr8WWTAvMeReZ9Lw5JpREIL42X8druL3cAi2QA8hU7PIH5390k
KNB9+4ak3x7Kqk37+VCNzKhQciXjk1KT5vMGV6HuScAI98wF2D9B3mijILmKBxEn5QpHI8jQhPyW
BJAJiN5wFCFpqG7P7grUJskM0StE7wwVbAAQxnSpRhw2zOW1PFZu6x8jMWFDBVml3MPOSqUiy64W
hcB3wbEkSYt/34MmPXfu5QccQ21PSDKMdv99l1q3QK7IRkq92vJrfjdeWmyRg7G/o1wZppMKuBib
tXrtf8kATfAsffswo1i0XPgSqz2na+Jwo8M+TYWS39oxxKp4MV+94ja+qXim4XPDAJ/oRUSX7FYc
A3F99F6jD1a/xILQgbyAOSf/ZzyXS6mgL1BVgbSnWSOePqPDFvpwbDGvqdugOH+vxG6/Xvs8Fu5X
IY/2AaHRDo3Rb6XNoaW4+cvo57qXM+lFd8tEoW5hfMgNyE8UqJjOAmaxXdoIG+UKYylYyKz3Ymj2
pn15RSrnmANNnDj1LIRUzGfBcS0g+GAtZ3BOvEwT22iDRSM/CT+PLjkbMf95RC7hjhaOr19Sr5GL
dO4NFZxAjq3UsQ8kGvPgmClGNYdWJEE6TL57bqef1WN/MYYwku2HLsmbfGQ04VJPt57TS7hM8SIw
t9QvPPrpcOpf75oxot1SXBM/lKRiMQ90F3IQT4/vLKXqZvZdn/bwkmR0cnnBEpHz774VPCGxEK9P
fM7LY8bCpzTZgpty2w78lF7SCO/uPVVkR3Ej4P+4YhO3W/BMhlSBxPaHhFPGCsQB6juvwXq+XRhb
AwRcrttPODvwy1BtLmKVRWOYqTNxnzfm3AjZLJkoWwEu1M2kx/949OigIKwOG1e5PPaV1dYGkCsN
LhwLkwVU7QRwWVpdGh5WB6jMkHHRGmd/xa2qGgMVyRXg+4BX3L2103BmFzsGJgxTVUYwiHJY7gVG
NQA0tG18Owm4I2ALX7T/b8qb4K+OMYlfevbay9Uoedm2Fgj6DAJWDGnOn7JGoK8NUh4CFmwKaI/E
1y/YbqNgf6TEaL+/pC9+VAwGWVfb73RRyKLfHTYW+7AYN5wUV50x3DXN8D94C0lRzDE1+5zKxcfz
hPVUKStXT1g/5azlqrADs/lYHJOlD1nZEfRGw+f9PMa9rzk1mkTPopTWhFbNad79DwxiOTlfHR8R
q0XNxyUhTDFl4Gtx6WhQlsQ4NXM6ywisCNL4Jl/HCarlpnwKWQD7ydXLXNgCw80gk4k0+BK1/YXj
ywWiUAXWeVE0rCGvXGVV2hxCCpLPoEj+PqnH7QigR8Ig7EJ+WjOgEIq7vh//kdh1sXO+oTC51X7L
1lfeD+hh28rXPUFlNLSjujUdyVNF7EWd0wtY0jh2zPEpYoZV/2rb40SmKNVhWZruMAESN7vgJnnH
1BNKjZyD2A2c3m1P/cKGKcZ/BpTz3+LBMl+wu8z6H8+VswdSObfMCkHEyNlfJK8I5D671bjg9QXu
fj92yC+anEeaRbMs5A+juhAZIbHh5/e2ooT2t6FeA5UL85nm7NEsoDU3E5aMzMCE0bMYV/uPfMKf
ke1hOVpY2rxOdTfSEg/fffnKawHdIkMb/B0mQXrJB/zLPOZcnsMofMBMGJULaOrV9LjGablxiOi4
1gD65rHfDftB9SKi/XbmhlzHLBglwVI/BFsMrF7rH1CjMPNBbONDB+HJw5a4tRrJM8dR+BZpZC01
76XqjTz1gADZ5YNT2u2Scd+vRY+0qV2zNdb2WsNlPVLXTAenRmwzh5SdAVRtAp0EbLtl6kB0caBz
I0fkl3qbJZZQhIR9DEdkiutZd7PVuzSnTiu8ZfNr10CobsK5B1ZHykhJQUB5nrrxaJy9QfiIRqTO
95F50KZ/KANAKy61KJtPUd5eS1Eyf2K/bw0ZQPAJCviCaoEuqCUrmQZqP7H7WTqCT15C5i/pzW/b
Q3KITJurzsqrGxMv4zlnMHtzxEHV2uIT7+HtLNKh8w6I/3Wrw8lmofVTKT0hNjLkLgpzLgGWWnCT
LZWWIDMTxMfOtPnOdEpC4X29haO9Thhf150m092nkc/tUDmtwTksQyIyaHW8mCucxrgVlhkyKo1H
2+HJX3MJsKGD0AHR3bPH1pIv2VUsDomlXz7Mna/12NMjeD8OwdcG+XBaCZEAzxCkIFiOT/ap0HcA
hxvnFALpQoj9gq+bxFxPPxhSMoSypE2FNXDh7DrXKMmW78wO8O+oMCRiA5qLS68yoQVbcagloyFY
bM4nuEN43edbv1PmuFWBt382OVI+GmBe6+Pg/TslC5gzB7CEkWJq6JwXpXxVHybr1ZjqrFlIMgAQ
1TsTazfhKeJx/Y/Lqns4irwUT6tdE5uBIlSXLLHomwF8fV/1MFdZGtmjq+OHVsHnWWTQabL5zjZP
DwtBwDc2H3z2AgmGWqIIMsBSjrHF5mCViacvL3EgM7y++bM/4ELyrIQbBaoLc4B+7Y/n9YHCSel4
gzwKqQB98qBvuKsrUwmNoZDMS/35PDpY/DPWGZUo6Q0lixv2RTS92dqfpvGwPlyw8GsikaXoLsqX
pVJcvJgJQ9s0QIKb7oWTT/XqO3ZBp62I2hwv9PiamHWcf7khz0U2sw1l0Cz4OgLIM1zP+DUKGzW1
ja8wMo+KoW2aNesrmHFXODoEtMrCUUQsurx4PQ3EYaWrTpXcsM6RzHnYczytAQLpH0+ODGV+e3pR
cEEDUhf9u99XQoBFqZfZPU1EQLZybVC7aoycSVVxoAbVwLbK+jGgBfoOmEpU1HycSsYfVM1GnYGx
5+LiJlnif+c7019cUonuhuLm3hE8egi6tlmDmhYS2/U1PJBlfEWkT9Ym6ILKNNI79dAZ6C3Rz/gI
j80xVgeBDX6WYoWumh6vOemltoa00AYkFWyuHlzWGAiAE/2m4EUIfB031NqhMPYjohjI41OFs0Dp
JVAHPkZWCEM96m6gtmkAdrdz4u5lhnNmQTFcsTJwNdYXghc6l8SFjrIVhqNmys2nypCZ+fvrhq3K
DsULxTvp8R0e/h4SJsW+tLxEWvPh2kDTD1BxWFc43brPSAqdMDYNxtyDp3+lQcfxfVGN3q3gVSZd
0sR5JXq3/einXio6XL7KuWo1m3Jbvn/9B1GhOyZeGJcCZ/Kb6WGadcp70ZjToYHtibA+LDmNqayy
0uU7qWMqdNWN/M7SmA3HjrWLPmSy4mj5eLbgIwK2GiABykeQWyhr7Ezsk9xOHCf15lFglfzQHVH1
usXrKZ0x6glG3fUOTVByeLLOWLkWiHQyoRpSuAwWcr8MHAsZI9aH2KCXmwMbMhbN4QkwS/Vn69a3
FP5bNylddSS2KbuxWmiAmHjBehZdvwda4CuRZhZiM7JUCTEEjolOjZHnNrJAnJvIsSGfCOak3+9L
pFrbaxhaUSkFDHX1N7X9sFkUvvLht2m7EjTdl2IuzYdLegFPguU0aGUX6X06RhBJ40xGppO/g+dA
Qu+aMMr91Wl+P3PQHnCsUTojt2fyIdzlABLggMs0R9pkoCo4V6k2E4ayVYFBrZuS/mHnC090rySa
FAjy0sWheADtzIOAimMBWneq4uGzHw+VgYvb7p+8QQAn+QN48R+X1jPx7/SVzZvDgEOrzAC8D8l3
AfOC7NMpIbr17EbsHIwhYxucxFUwzHuAz0oHhCcVIzgc0nWo9k2081khOnl7315aLlVnw0ySHhWZ
C0nInRHit1YF+UEVHhCuRhrCMSdW7r7Y2biw9ksSF25oCzHS6TSj/52oMxIiy5KAX93MDQkW8Y7t
QaBiHPueJmJuJB5AS6flPK1cmwzuQW8eT66sI3RyIZgA+lLJ5QzxufS7Yct2jguEvNK5FQl++2wM
6smDBRXm/aF0tCIFDUKbOunjs/VHWb0Hw2xR2eiUGeGZUiSf1WDUI5ykyIFXlY2UR9SaNXpdPBqQ
qRGS6f+3LA3Ec/bEtC6qIpoM8prZo0rx/TeXbLSGY+ZRYgO17bdovDrHSF0R/5CRGhmevCHTwvqG
6mCpKeurIx0zSaYRJQQoJS1yMbETNpvkfBbhrfW61usqHChQmweKrHV4sQoyVPepJEjkDKb5XmRw
Mp3BhdsVThYjG1SHxDe8raEdpMmmNmipnu7XUyNpWaH/7zK9X2aE09y+m5wccy4wAN7LNAk2C6ZK
6j3lK5u84BVkO0YyFFlli4SpXpgquv3D94e+53lf+vgwaLKqreZhQ3EQnjW8HgbQ4xxH4yN459VC
E2wPaINW3HKWoAhmYduYd3niVTp+9tq8C/N85sNnLgFA36WwGwFJfTApAHXkWFn5rJlFk82DsFR5
o23TjdruwI9rc3cZlXO3LfxTzaJ9bHb1iAhywQeOlJmbeauUFiad3iNRKm5q1fRZ3OBZSheg5sUL
+Z8rvZBLb6l7M/nh4wB3QeuOXRdIgeoKXkODbD+vm7/ONf2dBjXKZp1D0FwNTylHkuii6Fb0lmUB
lfoypex5aTo1dORZ+h3peuPTl01KZbjz546Ytius1bDWI3AcWJWZYVtK/hNxFUCmh2Ea5CMSsUGY
m3DATK6YzmF85/rwyXxy+f8f2mDUTG0010mXTk/22yg8/uWGHtmahC4Amvku1L8qCX7GAPiqtCxf
vl+12wnmWn8igj9prlWt0S4/2MkO/9bSABwQeH1G5ore4Swh0t/hjWXmhdqL6feQOIh8ReCola3W
CI3nMhWbnGkDR8rEbXTJpe5zGjs/YkMChzx41Pi63B6tu3xuDDazYKKAjKpq/okzX4/HGXB/7ZQT
rQ5lECSeOts0ZWIQ6wi5xNDVXLrZeNgffWRDYdlEv3TP91zBz+A0P4NkdjN45fRd1KuGB6oJfbXC
EIjJRtTtl0WbVLmGv6ZgzKLx5q9OB0VWM8kFET3Uochdgy7R7j8ichblHaPAHg0WmDwoc9b/bZNZ
UvS5MSsfNhQqCftFcGKRezWweNWWQaPxAxuwQYljKOm6twuCIV9hYG6uAKbCV7Iv/V0rs99SSnnT
Tq8j07J9cu01XKXkD0l8GVk85F2atAZgj+4Zgw1JtqhArkwcjvSZQaIheSGssr7NXnwRcJ09OPBH
CF7Y6nefiAJaOLFPc/feTvRjoo33MyojU2FdqNx1jZpLztFtFIIzpRi+53OVakIWwqGbApP/SkoX
qjNz40JsBIfJGSOkYVXqg7mO78rXOPX208PlKR0i8JYTE4ugB8gu71j9+ESGirvq9Bpl69v3UuWM
n9ppbvnvj7yaIW6ZIsLI8fUCQA7EJ4kh1+ykMbKizdIplU6Wy9neOBNzryPq2j6xWlyE2RA2tq8J
UiVJS6N/biSA3aPwshwvdYupk7IAh7BZXpQ+L8PDCg/R1TgRwESuW6dzyVFSrf/MHRI58jGodrPg
Li+0cZ8KrcZ4My7hPqt0xbrDzBHBA9z07pEZz5GWjsUx743g1MlmndizIEKBeL1O/KPWX2ZYKHU5
ggrA8coCv0uPRnpzfyiZFYz0hvLaaoe0TZ15/ptacijGvdi9ZYcVgqmtdX9rkFiNtrGseigNeLuJ
CnIlCKwEsGor1moU8p1rim3VBFc5ZHf710pW2e90Yr2g/9jAvMnC5NYvZ+gg2noVYXZSiTAMaev3
x3sBGLRQ0vahlWwLaTCwTPfI3S1aS5ANjZOJuDWZS/gdO6pbcRkoZz7D9cPgSTbmASfzj/SFMoVr
Zpbj0J/0yXQeN8uMQn7FY2UoVH66PjedH8g4epU9fZ7nUGjkSmssBmh1h6yysJfuLOFe2dE2H1wQ
WGDWeJ9Itrep2+HIY9BvFwkLvO6jlr+7+CfCPgDA3cY0BeQIK2uB7H4eCAGu+5xR3WAOhzXKdrY5
IkrkCLq4EUEoN8k82LI3RpT4x9skSllAT6N9IpbETYw9Vr7Uz/hReZ53+rYbaSU+fp8/4U01TNrW
GzAybMyJuLPpBW8cCM2eZ6yA2bqIDYnsmapwvcfEqvKSmXmPDbvLe/X68W3X3Y3NyXakzksxroVt
yxFUPc+uOVgvwIyv3g5/s2EGqVnZ/2Lqltzrf5ebkaNqJo4Y0O3HR8ClVY1DAHs+ag+jGMbt16Tl
WJrrx2NhTXZj8VQ//QqltW1g2LOGQ4pYSn0SH54o1WtvZtxzFgvFs8BHzgqO7Tuy8q1nmo1qBKEQ
3mLLC2MNEvwTG4s1a7NHQafHXWK+FQYuQGCnD6EAfJcEM1L/VFw1YQyoQRGjgE/SFfB6n6tKdrN5
93v4mGAx1LBTLUiH5CfOoO2ODqL0DEuvFNWbs9nqcBzx6e/WFL76Ui0Te10CFhS4rfcLuVCtHEs5
wa8zn3bBMmdDJaAd2GC2ioPdRi5q0PN4xENKgoYABMTvhPV8LZhWqzjPx3+6c/uD09Zvb8Z/iBMC
/2n0kd8zgE3rOxezHGXPq0FbrgzbeQkcHdam1f869zaOlfzYHf4odnC+diLcI5EmQ6ccIox0hpZ2
Rky/gbxPlNs/CdYI8VryleOkYZg/jz6lQK22l/iUKT/h7lbJp9aroCnZQUbtn0JA4fCY8qxfWkPy
56Iye8q6xJ95JmnSoAge8f/TEs5YUr82SqVz4Yn1wO/bENrkryNvwEOo092Yt2ngTcc+nd4SRGMc
qmRfNkvwkO+638isJlJC8WlahBD3OcXHqpprJv72q62D/HesuBbgp2qOalqikvRf0CvEPD19ZVvh
NjkZ/wdJeCII3k/di4FeaDLZOaNc+RAT57acjgmnW35Ogn3Y7VkT4qBg/nGCZDEz2UAaPet9MtsO
Xz5lAo0kO/N6ujLmIAkPaXPDNB5208vEjK/qZdC11VyNR/h5j47+1bwy2gWxDblRwBxvX4zDLFba
qF8nfOoMfV2TE46ZHa7/RiAbK/VyrT7NLyTzu4O9PkxsX+mhkmiYn44GRQYYsHacno/FjNX7sAZD
dASFYl+/sMIPL3bXqdwo95BXC2a/S06LdEryp3nigwc3dlo0artqL4w1CM764zrWYIXUe8x9VPlr
jGvIfMCQwRtAIriUnA8M/vzaHCGZ8veJQpuiLd5+fYhh7QuwEH/oSX3c2L6s7LBePQnFWm4apUah
5oXmhSnE3eLfxr5RQQG029GJ/oQm1lMNDKHGAiTlbMz+QTdQ5S+0KistWyMSxDonLG8dopvYXCIT
cfYvE4e8N72VyussJw1+n1hxcEedSGqWQWAAz0Jw14Co9uw4IByWTHsC7bAdTvr0AYdsn8XWqLSI
vV6IMoypsqyp4FV+tFlnxOCVljTrbgMdcsyBN00foWjnO7Cdb/iAAu1NiwaEQfd1BLxvprT7xVKV
IFhu9Y9b1ujTmoHtcUa0Q/atryJIs+svJsSCGL2HgNHPrfO6LDDj78cVp7gPRG73qck3GEk1Rsct
rAk3NGH9oxbLMBi/jwn/EktGRCwqOAmKVwtj6HwO8ZEtgmwxuABWPzk2auqRvCK5V61pCrtQwqr5
Mhj+VplNhYD20HOK1IEsyHxuOtnCDqdYVGsECeX5LMYTWz3cI0rjR7i9lFPOhAxKn+uZ/kkh+9aT
n8z/gj1I45u+iFw5dBAWstNUkU13xE87RcXvartdFJEdp1SVKwBKHG5qFx4BQPk7zr6EY6UzQkjI
Dl4MCvHw3/RP3CU7+JWIcwOsKWP4ACLphztlkYhpDANG6S5k93XifcXoMoBXbxct4yiU14XkjeNv
QbFloe9kKTK0OrgOg73IJJZdEHfCeSH18vwyDCyifcJIfQ8DLw6dgMlSYhNgOVSX+qED+p+gd6N0
nhR6x8vMPGq3NkUMHyOgmYMPAcSnEsAY7LSGahZvDap+Wo2xSByAIMe32lswoI9K2tZL1i/OCRI5
5kRLQFQxb/fLdCJ4Zkq97mzUNsELEDfhCNkc25duq+u/EJtTNWM/7oVMRTgs/0Mg9DX6aSED/NGB
8DbTNq67yePl11AD7E+yD4V7e/LpZkQZ3RcaUsSMCIuawqR1TlXtBbAyTzVbcpRFYqjXPEDrX6uo
BNtEVqbD5/oMuDCYFP341qwI8Sk+26x6BxyJlVZUrOfzRNWdunO3WsVvs2Kev67kemH/geOErtIJ
uf9ESPWD0O8YfYfKe8zApB+0nycNjWHKAekD81OurJOq8ORNSxsr58J5vryQ7eJbM6jwqOeFQLx9
tUp0l1aKX5i92NwueRq0Br7sZlv/ojQvBmqe3lTh8UlJciOJ7VUPuZECU63DUuanU8qOfhzJNLG2
ulsKMfFQ2xTurQ7m694gOIZohad4RSd6lELLezEf8BbspKKX9cMbPpOUC5I9twtCIyUq5fc+WHEa
fNkrcSoQE6YYfZdCAGg0MqD5SbK3kQyIW8zt0gKX1dmKoPIG1ob6ai23BBG4p4XVBgsDdMvuE/Sr
iuCcH6aUtIsYt8+GQQwtd9xzh9tEUUgJrXSB86cOU6q8eyx9qHvQU4T1Sx56JY1Mm42yMwSRgoKF
lJaDrZ6xcZGcypx+NTNf/BzE7bzYCYLPlcy/lKzdp/pnt598bLzDVsKZIvZ8mfY0Qy2c/9MWK/9S
f62CGOjDatMSKoMuT6dUgjcTG6xgTlzrEYnfceruiY8WYhboIYhVYnJeKReS0v1EnNOEx6p3axYI
e1yKvJJ+uFwiouYCeP+mQr4wlmy2RtE1UdaOHyb59WMQqdOFj7Pwoc7HWIP6SoMdshmZW8ihzkqD
uA0SY5vwoqZQliB0pb4ZMs+TMGFgEr++n5Wx1ALTOVkuA5TwxXjoEW6G50nWm/Kt5s7SCN18wGXL
e3EUGDyMywqXYMHK7ulx+oo67ynwPaAdVrA8gRbLcVYZqxh6jOI71S1Ul4+SFvWhoEH4N1IxLYfo
VQPAH4rqGMjr7DcNFBEczYdUJuljD6LYKXGPDJYLBrG97ZPOthNrKxuMxoXK2t9oRb9Z5cwWHP1D
k6S3DWz29KU1tUsqC16emRVeSyOD9Q/WmfHteMN39+43265SUBer6BAv9cC4rSHgqCwXGwV2nM7O
AHIWMG1bQlRzlLTQgfpcFHm15hAY0RuC0gUkFVL0AQVR5Nm2p3fMaKna+vxFDvuhRN1+ZMlZQtD4
kIQOyzzp+qAybhAYEpprlE+6njer1NOJw1nRT0Svi7dh4HBdxxlLwMblW7LFVWvYqXuHBdJ6XUcV
c1n3/wT0whSVyz+UNX2xgnzGBtvCR9O/JqEQMA6O0offgU/P0HfIWGBOx1ltTJIu5Wz3Wm7D5iQw
rIaX+/uHJT6259VeBelOiX6ViobEXA41QVIBnYP6QKMqgFpV3db/aLu2DTWQrIMio2OZL5twgpBU
qcLV/mJ9N6P4Yn7/j/9syzYt8wk7zGTrb5AOKmnZ0slbFV5JoBTpVYMKB7sLorCHl3wFF7nqZFJS
+7cI+wLOUpXVRscWGw5gJe6Co6QGSRJYrKEa3xujPI4xW/ZP8vpJ7efE1kGOj2rmCHs/07ZORJ+t
kkvE4W4g5OnLTmed0vzDKGQAL1mPjctoVZ4KrrQjK1cNuxvEs5NTk/uHUNBneiSAx9g2jHun6x8H
gj98nbhvJRZ8bnaxlazz0eqhLwKjqm3WVgwEU6R2w0KqZEmcATIcB0VRKD68mDcsmS899rYnNgZB
yMNIc6oxsnOZv4atHjyqWnVdjvz1JVJfVj212RCqn9jeTAg3PiyW98QY73pr+TqX9usea9trzTPG
90gvPH8SLb78DnEIqKsaW+RHcoTQUQvPxYn+p+xDGT3CShqeOK/YE5oZx0QuaFhTa7kxFXuV58wD
IytkIZNnaBPS7Li+xssLu23jrgtqgLna91a7odz00uyN6kmSYt9wFlSkMvGeeSCEPmLthCUmHOT5
7J7lknwe1pLGMphZiuHSfTCb+QyFk/McqUkcA/wsOAc7XHyF7aTFq/8q4DySwC6xjmqcvjNQgPq0
AAxthr7E8zjHJNrUp05iAbWIXm8vROveSKWfYHPXRk7ldNwb3ZLEPCysNjP4qj4228WscCaUVM9g
SrXYcz9/DL/yxZdFY1JCooxQ/YdKpcZPDMnN0ph5WR5LZEkAiMYrz+/5QHEpUuqIGWHrBgTUOeRJ
TpgkLaP7r+VisSOka9NqTfiMXy3aAyJywXfPYnueZbGr/RypKhuib6pZGCPJWeNcOt5gsdEVZK1T
8I9jcjZeVTYr/ulOyN7Qfu3gnj3EOGhb3d0RKYqk5B0oFFDVDfg810mZp9GAg4G91Dlt0cPZLGmY
Xi/qaXLJUyEEpKG1Qm7KG7jbRyau7OmkDPLxoPFyun/UQW8t6W4OONpv8FDlU05Bgh/8R0GUFUJa
RyY1Uoq9GJGf+mUeqX/PjlDT2g23TFXpwxPquPUoldvJDny0Qn8LARrmR7oLE0S5e9l33FoRmeMR
miMz4p0X+RASTPL8gIVZOmXOsFtM3f0Kk7m+95oDEdElTBOFmttvcFWB6WAw6Jmqe03qYe3P+/I0
FZCS+pRw0QLjdhGjMs6rsiynS5XcqSVpDXcf6qf3GTxvt8xlGKjgVzkoBWhJk9bhMMtMf++bO7I9
EdpYT+emorhWJYByJxC/sxe/Py5SGcB+XQQW2ZnmtKDIhdLPqe3kzRPMuKe/x4ualFfJ39yYV70Z
amlNXHQy8n/lfR5+yDMjQVbhhfAttYqVOdNQRUgp+gpDuncqyjUCXaCKNIBH+yciQ47eeZK3754S
tlUJBRqaBbBQI7KAdgQSiSEJMafBKUnMIaErqSwTNR1cx4TLoWS2HK/aDHE1MHaim1bZjSHOvk76
N0HkHv1vzCctQyHgwfY/LYdcGV+Q+2VeIaj9nx3nbRCCoBpbSHknJWSuDDq37jT9yRWowUNndLDd
ISp/MO9nkJ19hFHeWawgf9DZ9wRVhl9uIaE6FVT9S206Y1Z6POfTlKrT/HJAzFW0NyVpe1avVsjB
w91TxqW8pWE4IlhI2XhwUi7zZpHlv+LzTEmDTwIink271kJ3pK2K2VXkKIklE2ujkWqjrdFKNcws
qelHXgmeqelyWB/5Ej5QQbzArTKH1lq4QD9ryWMDHFL+HGCeiXdqH8YLSM6j3DMnEZojW9waYCNf
Nqrma3WLuVGTa+KE9DUKkly9g7vfME6VUh3clF4e134fmqSfYzFvzLCkMIE/xKJ9+Hr6s0GKQFPx
sej7p+pJmOhBGaT9DqG9ilsS90KU1qRsk9usFvImFzKTqJer9QLdxmzYeOjvpjR8/4Ifnei5MxeL
f9HYzGt6L5wJ/DcdUIrv2KWaPqOq0Bzsb9PPQ0m/NGhAuWtqgfCYJFoOqll0hu2dsfTgqWYb6kR/
wSUIj/SoJkQUIDFYo4BsulzLedngt+OgZ/HNED/KkZxLTVog9INOJ5uWpJfKmw2wEr45E72f5XnV
5fgg0z2xf2NcMGLJdgUspPTMeKVjGN1cT9WXHGoitY7BSm0y9HSfM6DU6U9rjJLhbVdhHzpdjxK4
1lYsPMxc68OYafFvI1PrRDk9zY/pZ91W/JWukpzAuiumkKdj726Xrh+6rGmwLMYtKMJzVJY2J2dM
Hup+Q9ZMYkLj8l5URPUz4wwg82WYhgS7dtRJl9FknslH0r6EPfeNOtZPQ31rTlC83k071nNhd8AB
D5iwl1LFwl1vETMsCBF+eLQr6HoVUD2XTys44RxBaKseMNs/Kip1BGJFY+l8Qp7Hw7Ve1Ihty2Y7
/zCOfSb3H25Smu6wfcqXDfqpJl9pkNNCpiI7WTFKkTCCmSjlQr+9RxLLQEBK/wbuKittoBN5diOs
z97T8C4MvERLel+ZNOeOtrO6vZ9ZQso8n9bPuHh/IUPu/sN0Jhl4mYg1yOfVJg05CjK9G1oGYXog
ySUQgqiLCZo71nhbH4Y7voMWlIsA0r8ScMBFgEtIfNfOYhpcNE5gLvSdENDGnlWlGdzMGkiMn45Q
3aG7Q3iYCJIH+xhJkTODgXMPv8IpDq1dMlIuEqUd2Qye8jRgVxATDnx1HVmOOxJkVv2IVVDI6wSM
bepCwvByHMFWa8ApJ09lyGqu2mArrL2eHLNI9DUNGfeF1HZbZlglrjbh9Imjn/Owx6fX4O0elc8R
pP6dYDLFf2JnlBv1h4sFpx7nv0468viwTUdoRWjEuS50ukBgvrmixClQnvn45Gaw+HWmGdRD/CJn
BCG2tkcrcsCwGub2SYJRlBquW70oIXgRpKFwvAyPD+VJZHGYnNVO7xUzeYnMHQm8DLsqnRe7UpkA
YeXY9X/rdSx895USvoJfE/n+WyWrN3wHfnFi6qwCpnnY5iCdY34o6uCgkjkUqrDqgIogIuWm3YGM
UM+bQOsXMqA6E3AVMED2iQ9/p099C70xEIZ3UpP7on7XTx71+KbZIcyFl/ZCkLBBCI2PvS//A59i
35HSfxWilvirgeUL3w+k0oMa9yXpb6M6NV89e0YwWufTY8ARYggmoE62dWrh+8Qjxg4aV5/cnzvK
WPWFNTQlFaVIu94rJLk92IKhQzcZZGvdpdCQ8kBfaRXhwsXsJ/1ezHW/QvnncsEvQmEjn0+KQXZO
m0r9ZknsuBeV9GwB69C/6MBQ0o5nDb5QNTS8eqd0sw3hEtKBFsmFajHk3DoIK+mlVtf88Yh0/mF7
MOnmHT7RWWz2dSP46AIRBs1Qv2bDel5QmHzCRQ2ck6bKOU1/MiDZBRaQEPGrERi/1Jfcb25CST0s
B8wBUpii2Roj9f68xMszli42y7xmtq1FtYdB9ZfJrWwV3Q9+g0d9b3ZKzb/K24LYhCRPQLOkoEFs
940V/eYZK3IlcwYWNBjJGmETUcyGbbB/eN+G88fw2F1bWGqQ1wSp0ftAd/wDYXaZ6k43LdHXhKtJ
ElBBeptEhaTdA+GuiaalaHH7yLKQktPOy8X9HQco+K5wObrt3HbO7JfqG9IvemVgzGdsEVWsKbKt
zZCj/3Yv67NbUWiErtxYuIcL1m+TjufHGQKHbxdjpyzjikir6eV7RtHPk/13o/rfVdwoCvMO7OC1
95hTMw/H/1Uxr4xWCOqeH8GGBKxg48fFAfmrXU8PcuXN+uwyAop4/a4mX9BzXmODE4ScghU57yC+
gWd7ndPM51iYitzY7sBdwix64B0IQgDnc1rb5BtBppIQ8UDLDu97o+R8iUhLHLUWVb2/AMiqkWHl
QaEXD8ifdvz8lm1uEktcRXUnxzBTtWUvhsESN+0bdZwQ5YG3v1fhSuhIfJ1MScg1J/vn+trBZkGl
xnmRiTppbvEaPI+itr2P9AGylWbnRqLtsEFJM4sHnrOQZIOXssXFyFyxX6wPGFV2JqJjUQGp0qtq
WAtMGluaFOuIXSiGTXLfV7MgcqBL06Caeqi+cODrWrO/YDfco9D7NK6l8WQoZ6YfS4ifNBnEf8eZ
yM88F3ZACGKDR25z0GVJ1QAKZ/qHpx3ocRVgDaSu5F+xq1Rb5+TopMVeUiDNQdujYUzkcSAp9ud8
S5KfdTLNMvf1S5u1qdFSNAW5LRY4ucQvsZgnZUHwc7bgnWKaCSBLCLWOwuCCj6an85dFUSGvNuTN
8BNZ5J1hSjS8cUt//wjn9FLzs8D4swBHn/zKsLekufZ4Ed4pkjAHBPwkarc+F8tF+YCF1XqK7avR
DMKX78feX3NQ/khvChjOPN+l26wE6j5r38wZ0vuxT/lqX/fpg6qEU8SqYA3fSslwv9r1wr04iStj
DSUqu6l+JcoX73+I/QaH7nlOaICSuGmHWK+UrxmIi0LfFHEiCjKCebOTPco73x+yENFU+UU3dMHT
d0aG/C8lTT1qREPrFmk4DzcaaN9xDwKuuYdN4Enp8YyuJF60F7syLGJUw07UImUmmpTjkA3qpQkO
VmoXBlkNjdU5SxLIGqoddkpv8ryozK+WeD4HHn3KbrXYEHYGhYsfRO1xZd0jHPZTDMCNw6L9SF9a
sWgCN3G4TQclhy83NZnNvqDz+Sq5f6FO68j1vjdcdTa1Ynxik//orkCjR3m3U7G/JGLcd1mfEn57
MTXo5jFp5JNFS3CcBxtDHdOtm/pnlD3K8upvYu3S6fi/m7PeGSaV7eCpGgpG/kI5jtyYLnICv1AV
xdcy1B80s9aI/fi/6qnd3cyXiWKO7Xhq0EPL29u9eurqLYYN+dbVPlQh1knVoMNWbEQizJ93ywKS
zMLjAcdbamfA5Ryc1Lh7qwkcyQAmpIRK6BRYkEbPEK6xkGU0Uklq17dlt1mmPzF8ELLpmlEci2b0
yoaK8r9P6Z13pZ3WNB2vIL0B++koWtVG7ULm7AwYnnszbJRQOBvExZDYLu/eY/WxhohsoYNIs2qh
2RINQYBergaQ5qq7n2fTNZLvkkFYR5u8W+RZj7u48dUaXe1rq4/H/ngtbROIiAZUiTsxec+IaPWS
0eTV1Ab2bFVsKKo1869sTDvolmkZ1wpRVAP/hIkEJj3UMH6BkQuVkdwSxca9+ylSziVnzHWeBV6r
fMZ0ifcav99wAqwCob4KwPcP7bTU2NaNI+3PRGUuttMaLMQr7aoAw/T3iKYj7zGkBAdjzN2IDoOh
PbNT7o8d8YwBvXdUX1dylFUk3/qDWaLuKIX18iWsFHweK7KUUOHQg3ZE78eKORA4RSR+YMOSdic1
QkmPPFshOljMoxpYxPCX8o7Xrud6CGPFD+gYmaIYljZzOsE3gXujkQ6ZOyY0L30di1anxW87la+2
uhCWDOswERc+JXZh9B5lwEJ01IQ8O7SgWqKhIgMJWjk5A3Gr785V6L2Dg2DksxeqMU4QNPYKuK4D
nzlJx1DZLeD4r9GSAlRFow23xws1sPKGqB79vCuWD9Fc6CfD95bwlrKoqBaYraGAvl3YIaa+WJA4
xhNvc4FZ7k3DhcQ6Gv7GNXpx+b6HMw2xVX1tcleHcWnMRf/x4yhFLsqT1NwK4wod1BUXit1ZG0b4
et4nTVbnqmlUF/JGWmxbSrDxfLiydsOHNlrdCjSt1onBEVHtjB/B6Pqsb/kaKHMTbKVSEOJYOUW0
c+Nkklu4MCq/0DNcPZ9FAXKp6LTsM30oO7xGqOPyoT6A+F5HPNAQ5UlNIJ8t31WSegeqMHBojIXA
6aS0h9Z2TBpOhyBLgr7NppV3vq4iuQ1F5dZasGAmptsAmDEtvMr3qwJVlB6hBPCVMgTM4MmVa7kI
2jKd59OHAWXiIEowcrPYQqzG0Gf/NtbX1Ru4nf4J5z7Ujk2kZNcs3i2tu0RkFTnxkc/2fshxXiRp
1y93P0d53Zkx963hgYqLdwLbne9UvEQZvwm7N/x5/iA3OZVN53GH4ymP4ZO5a2D06Ni7P2okxd01
62L1bDIRIrcVwtfCF9lGPuPmXA9tv8lXDh3K2oK3S/6tbeZT+5QyIc3apUTM/6BHWJ41VsI7+jw+
jcNieMgenQATY9Z+nhmunM7LCXYLalnqP1q/PZ0N/0rSR/8XqRjUARmsm+OTdo182Tie0X/d0+8Q
rKHreBRaja6Z7mBGu8PfzDJ6Hl08espcREmWIXybBzbjmrAByxKcngQ/U6A35Yr/M5xswo/O+Tvq
rP5/8BB9c0zgB5OZZYUs2jFj7qRSB5mF+vOZ7oLhp0U+UwbiZll6TVl5AOij/53TVQKhH7eMKpOH
LtW3oxyTr3Ix8N3JzWFk+KFkWUkNugwL7VVKMqdYlxxBR+mGoJO5psJOiBZXlD4ylzPGE+MrLb14
xd4OpSKExmaUvJicXUjDBHoHycjAmvaxBQfY4gNs7LhT2rwYo7JLjJh6hKBeXYalCsInb9FDb5q6
z+z2nQ2DPZujLq80LyD884rKoPdGt/9jQm59wIEWm7z6EZEZsHWsQXeLar3SiRFICCHvm5laIVCF
rqwLO+G60XPazKn2ZOu/XDqmDUBgCCjCYTIj4SzRsLLdmqwely0y4j6EQKkj6O62S0Z4PfcSjwH+
ABdcYdKAC8mliv7mctoHHQC0JCneO5hmSAS8Em7ue76N/vlRUDHHiSompEOxOxYxTmuXebbnfyFf
eHLmNAYFIyLftQ3I15AmE1MjaHhIBOCw/3xJF7PoMQUHhHOija/lbp8oP9zOVIaK+4Rh9qlIMKBE
NYAfLGDXahiN1NmRTQzd0Mazzenfx1obkCbuGLgnBRej0TPUCjMXeB0mwRMK0ebRUY8T0dOkY6Q8
VZapTCptwdoI+m4YI8ZI7eoD+D0b3nUQGZ4OYvB+ziOoSQ71L3FqQ0Qd/CV85uGYscNnLp4jIag0
rI3+FV3w4DfCgbkPJPSahpdS5kEKKxgSBwuVfTZmXsCsQumUZ3Hh8CGbbXGeHJ0FEhjSyUkZEQt5
pGekCtnsLqUaUJKNfm8b9+d1CzP+5x8hFj5xPth5zC3f7q7MifItsbACohS71ASY4cERQCSfiNj8
pEQ/q/t9jOsdLgFmvTghTfG/pQQgRumHms6PgVuQu3kgyMEp3JdXgz1fGaKrLOZ3pKi/QjYV6QW9
r5HV9cGWlFbQzLrN6H+THv1I6g9G9H2SSw9/uveF8uIloveE/FlriyOxLGWkuH3Nv61K1rY+bgAy
mlR2/n0TNZKsH/zM6owFaGv5Ml9XypSeHJGZdTePXHZvoq6eELv9jH3O90q3NbBwQwww+z7mqenH
oOkBtd2efrZG69CfI8NPhcx5fb/4QtnKIzwn/N7hYaeaN1a0xFNrMTNFkk13wkHVxPnE/hdXaBUL
zdzjKWlvYVMfN7MhKfn0wNPuaXFsZTKtga3fid4PVnQskz5L/Ak35CVgE0KKVIkffHzn4QdYaVv/
tvbmCIp/4KJJl4cxrkvjl7eGiBI569g8ddDIDDzTQtt7ELUvO6LlA5ZAbwowYaxn9Z9kKzWjmE7h
dsz4fVqcfKIIp7tmydrV2D8XPXWv2goe97vIjS5MN7tOcmUsCICoCGkT5kqeP/yBO7b6vTxd6IN1
gK/ypBTZiIgaJ+047Q//gOAk61rThwzqkGuUDb76ngp/G37LZBSFAUUONu4SIOXSfcivwTj1GXBY
Cd30SC2iyltLWa6mADnJi8Dvetm4gsufhuaTdzSvAGCT3NfauRsutFB6kdR6IZpFUKRkjTYN6H/G
2VJqCvoM9qsmKZtJ3O5/HfplAw5Hbs2Il9YQrbLAQDJy6DdXl6O2h3N6XnwYzWNExL4Cd7PYzGPQ
Cyf23tcqkwikEqMmiwUWpJLFEiltziqF+ieWfK75wVFnLE6w09uNnNznT4oV8t5qBSafFAMVT46L
mS6jFYjnAsVbHDMMwYejO0YV84m5ZJ6UN2NTUAXGO5vJ4U+Iadv1HT4140vqcHeFahjCx7+8oDx8
5DLmvw6wnVHZ0ix2gdqMVAt5Rzp+zZv3vXK3Gd38ZJdua4urtbpYOKQGsK2XbjHNohuTNr+ZlGgV
Yl6+XJdbNzEMmhv63wwKukmF63842URWoVmTl2lamqwOkkekW9NCLLcO8HopwloFphGEKy3UZE94
fYBdLv7b4v5+WS9edFAVzfN83pm4+hERHHGm0rlZoc3RsDqVL8guNw2y3jLRD419Zwugq6UZz6pv
CfreuBRZRl/rLXdupSS0g+WrjnVcFqlRSZpa7Oj/3weApl7PWZ4j6+7oPO1ImIqm+HrgjgBJZlHe
80JCNBEfz67n0NsLIVyIuzlp034sX388uU/H23qrL93KgU6OntUMadXvuWgeFoFadFdTiBtUBnZh
wYMU0gBNAwAIYzBdop4RmHZ4MSEWkVRZ8VYZIsT54LtaAvS+FlZLAPzAomwY97N1cOvBzFTxDmg1
QMwTZyiMFUP1cThzfhzMmI82hPUvZn619ojOUmzYNhoVCqdXZIcul3xNTsbTiNtXnkTTqs9jCC3D
DpOzE+KR2CohhrN2Ql61ndShTUgSw6Uy7O/sVW5NRscPtKuCSVP6wI7y/6tx733ZR5Bwt7FLVtMI
S4a/rcaggVGogS9Di4LPAZeNyiAL9PU39eeIWeEs1hpzumD4TrBiugcqHNNa0hbwugItHW6WPKxe
drSkVWquq0LSTgWcApEc1RRElBPS32KdgyZQGvSmljMPE0XXeV00wKHxhKWJbH3DX029vw2ESWmg
RtIrq5OIcjCTTGlwmFult/gpScCgW84TVhQbJWkZxm1qryWEBo4OQsPqAamZqJTmmXm9axOtDh4V
eJqdQNe8WdurQnd5KNdKSxm9lXZax9ZiO6c8hNEPbdg8L76vlaOUUIpjpmjA9fvXmO5taLABPqrz
UUaEcZ68orTqrDOhpbpEwRZWOqGJ/u/qMEP+rRmFzf/wpBCl2OeU/NdjhoKwKnA3kt6altZJAdpp
AQitiYQESOl9wn+D9pdQ9TJYLKTMu3XDPtVhkCC9ThcwLopk06AnFiDPczsY2gSqspwUU/rtRPxx
LXz31Tb7wWo8h4NoLMcJgAfuHAIY6womnUTJ8sJWXYQUjgd5VDq3sLVL8x5YALmQfEA/gVVp6XTW
3HQ9zCNEwkct+q1l0hcjvEOYKofacO5XKnWBmrJGzeVroFIDeY9aaQP6EtSimWHk5/eFTxK8meec
61wa8ZE+KxnwQhFijnjVJLZLtMn3vijWGt9638nwIV1fvnJlJtWXG5QbpnTmZDRhxiH6MJxAfo46
nrI6BfLZKz7UKuSh+35K5plfsGZMMEzBOpZgryc+sQa2n0+L24jd7e3X2+fHblX1lgwoTTaDToZB
QyF4Q2qz0nb2EBnGbHHdO/6/N1atfPyrcsIuhBsRKjcUcm8tm0O4gu9Ju+4kPgJLmqu3QLocOnLj
hgPOAHfvfbGroY+pqCZ2DwunR4PywnOPAhvzo1es4CzE5Jw+tpp+ZGc1UOdBVVzMVSk8QKMyh+IW
mgxCQoFESiAozxl9m3LfHwyHlCOG7Ft8JMjmk17iSO7LJFTGoDNmTFb8A+tEzriN+HmMZfAEVcEZ
CSR4/D2z46cNdWrHlzWYAUPwUTojvLz2qO04IDCWajR3z5RcQerp6ELWlWTedEUITLCi4nOeFiOT
bW+Yhof5ADV1w7WXi4t89F4mPGiVFAdmZl7ocipZOjkLvnp9OOXKC6KQywlSe/w2eIKlPO3Iu7va
GAlCflaXOtCEf+IZXcdkb34D6mUJKQHkB/jsEyVA1Zo/Yi8XWv1piRhcmd6DwaElpCIeSxQJSy+u
2TU2QZHdcs3gHNvAJ0y7BIVn7NBBKuFGI5UNPBkM1PaSIlkMIOmysJ/7tFpDsIN/bCmQvt1FtIYO
qul98BwleVRXnFUu9WjgpXj0fKIiErYXi/W8wvpDaQ+JlrbEAVyuMFHZ5YfCEWQdHPjJkFxmJg/y
zQsn9BXpD/DJyP1xt3MYMVbnwdnp4Y8bD3O0QgphpQO+u2jWJjSZ6e+ssYojGsWYvO4F0djDTHyI
0aFSdUkKUnzc91q1SRtwyNvuBTeE8mAcRNDcNE1/EsSniV+wYj7y5mJl8Wb3L3s3SNr88KRk0vBt
0WvTEFhW88WWz/tUaF10SpCdC19oIynE+aHTiiFgyjS3HoNwF/40zWJeGmwhSYuMolEqskqrHeDh
9BxpeI2/+nCEaAMc+GKj5PIAaikP8+5IrQuUHBql/bCnY4eX6OlwSYx6Ly7IwYZrWScGZ3/prGZ2
3b8g8ET7oUo9bFv8wa54SdOFM9i7gFCPYOFX6B4aZYHXyvk21QoC6PA25aVQhDH2SGiNWRhigkwi
STXCtyH9N1UUM3tPIOTR8gelGXKP3lD1t8v8UHxGLHdUR36hJrytO0agxmoEdDmSSYu4xYcyjyYq
XG7id2sjo9K3YoszUo0GnCN1PeZQdEW/NrLL5M7UjE3Rd0I2qgNxLYyR42t9v4oJG7ENvo4be8aV
NYoNPC+pIAs0pi02MwsMD/IKJK2XiBn9RDnaA2QZJTyRn1/BPKIUMfE0KrVGJgJVhqAKPmNQQA3L
Bmh3lLaHxPypV5ZAloqXAQD856y/A4yMgHn9HZI9K/lFmtmjkjcf9cF2VWtHLEU2Q56YhQ2x1GMU
po1166f5OnUi676/D8cCLQaFIbckGPlKHzJFKd5ifq61KT2Ev6BU+7CeU+xZw/n/lGTroK5OjUb8
ipQUiICt5j2H1ookM3Edjx7d3KMBgT/w3t3FrNsf4Wf8D2VZ8lwXpHPjd5hdvjnE2YN3OgqMWLHo
g2AvVCWtZ0UWjnC/p+J5gLKjwA1cxom5Ys6ZV9r6b/0ssP1BT54aZ9+swAt94aWkyDW3Yjk2scJh
Hyjj4H0/sqvFK7HR6XcCcv73VKK/gtXq2J9w718ux27FfRaF1T5Lk2L1gBhWvw1lzHZLZfFU4pJU
OtYgd2lORnG/XnpH+Ha25MtsnKQRbRZT2wN98YN3s5afjkCTt7FjKxXGTPcdtnY7NaRhHcn/7kha
NpThGaJ1aCWxaTR8zM9iM4rEyPwTSsiaXl0FVW82dzZ1HWgCqwyfVsCgY/F2nYlAXS3rvuxhBQsR
z2W/98QFs0Rggp+Z0j4Bwxqe/anq8hzuf0mi04UWbw7HAiGhleHtdYAMhbDJQ2LOLl9wcTUx7kfC
UxlYtfrRJtBNOcE9n69pqlU67l9aQ/a4edcWymJAfnn73k/K3FdvxmXh+e1M9RHtm5IjFoAHyrjf
/hWn0G4ENgR/Iq0nfPfIrYMa3VxUdrUsgk3JW1h8S54A94s7j8MzOKoS7dcQdlluh05fzxktQVRj
Gt/6/1p52/4Fl6V5wIK0EILF3hJ+FKV/KeJL6yc7DOJnogAgJktYNLBHX1yBxpVm96cNdKqqUEiL
dtXQAq8yQwCk/1ot4M2efG40498YNjcvF6HYWQPmsN80vnq+I1s2BQV9F1kwIUEK4pPHURzs9VJq
vulY8gfrMA/B1JNl5ShqvTYQvzrb0hxNvpdVqXHSo4x5H4E2DyqDLbOC4MXEHcNp7vs0e7n95HXr
QfA7X/S+NJiTVs3n3oFcd+4w2MKa+pPDRgyIzUVroJBznnI5xe/ThqdP0dmvDVCn6IyQWLIollCf
d42lCqKwZ4raUjxQK3iCVAcOmEU2AedfPiaFxEJxKqV7lNqPtOVibI3+84pOdLy0vP1pGeEJ1lI+
glefIh0YjdjduTnNLb19LZcgFOfsE+JtL4Tjb7LFI9i0dNBTLpzVmM/EfqnKJijOOcBnq4fd1Zv3
35IdINO7r73fLbe9mhXPTb4uU9XkB/yQSJErpvbH8sfYhYrNrIEuz1nYfdj6+AFT7enQ9+pW2uWh
XsT+qDXpLLoweq2EgWB/J+5b+H+vMYW8mdyT9Pb5avjJww6flhKkVXLNxwJASFP+Ip7Nqx4fYBOu
wxWCoxKv1CipLPWzBVd4TOXZtEvQ8mKa39r6QsqfcqajnyP3/pBcfLPZJMePN+P/HNTjvTna2+iy
peg3n7haq8MBD7mM1KZkusD8xalSp74kVwikbxFWQAjMIZMrRUkq7Brj2Uu86TGEWezbZN8CLper
zIgTm8rN57U6diAyovBZSt+LBM+4flxkfYIcWsgqHaMK8TV9Jwuu2c5gVkprLJqqGFigsp9s3pW6
LP1wOMmGYpzwrKJwF/kQYR7Z4TDKTtNGbkGXeUCutxkEvxw7vUwMQa/jb+ew10uCtrsvS0U4ymnr
nZqCvKzXBiNgQVPFpQ+7Zgb3VvIIM+fqlvOVB/h/JwSItxdE5Q0DEB/OxBNwvqifbSOp8JrH/BvA
w0QLzvBci3fqTpy2iHHbKMwp1zsEagAgaQLFHmKV9Ov3pnpL3Ge8VkKJoWrHTc3hMYXAaXYvIDzN
x+P1A1smx2+H46FdfzhRPDpC5lggJ9YtFx60zvSESAsI6/5Kq1qXqL2JWkJvYfRKCMk0D930X9c1
5pO0ScNGTwQPnpwa1UX7UJZ/2rLUyKqP36CM9PhngzBgheWjqEFFKaNt0gWT2lZN+c2TJtuhP+C2
O0nKv6lf6xhQu9yeXNm73E7KjzhOo5+VX6DgzJ+IchInER91AsRoS0oy4lIljcpAwBxl4Rj2970Z
s42EUy/TLG3YaGe3qgRfCcH1isVOpP6/fLgCBp/IJrLOwvwcsRtm1fBrWsPbz8nFncoohyDMPbCo
6m+ZhIpksXENVSU/KoTAjca4TWBBiPx4Lq/aR5jkzoQQ/ioPEWIR3imb3Wd/e4OIWJj0bY6Oy+Df
OqJQCk7GWic6142ZmWGbCqLkMcpLNDQAKlYjj1inNb+0Erl8zTlql9OkARBfceBSu6SewAGLW0oz
pQmMW4nbiEqo7odvZ/J9RxgKikoCuN8m0TKB4tkucIviaBii/CqiBA9jqg0+XeWQ8uZInDVWENZJ
aczgOANGdlClHcuUrSDdUN/cllVJrTVgyfVAqiVW/kaFbQDbWOzq33q671HHWtoaQ6PwNc63ztmT
3gFGeGeobteHH4nP6xVDZ2zCzJUnpNKI7bIY82I1uSwJE2nTKzqOvZV7yU7QBjVGXuZGJ3G2pk/h
br7gP+9Y/vtXIeQzVah9aq6NUz4fnwvSIBfkcH18v19NDoqufvFi9VWv2pxfLX0AQEqV7wANLx8x
4f58F/QTWpBFVHN/BK0tixuW1GSd2duGNuT2O8bS/yRyjfDY7ofpULTtijendwezq7dRDdA5cfi+
molelAgjC1ij12U0X2YbWN0HOUBF/NsthCL72k6vmDsddxmUJe1NWeGBFjZGPt0YKbw5h4NVUbqd
kKleITc7DMnEfr9OsUOZROhD5T2CQ6+J4RWgF0J6HM8zIo0ADSy3XsYpFFULs/VfNny0tyWD2M5D
B6rJvVwDLHl7kMbhsh7E6/FjgjCtFeT0EgizU4XoijDHRiMTDYu66qK7zEef7PeKVQrh9C5vqTpi
aMxjSksSuAhmw8+eBX8JIPE7T6M83lcRK53DIfHSz850t4jXzSf3Olv9IbJP/SXQbDo6SvL7Nw/W
/tjCjr89xPCilaLsONnOM0M/ShSR9B1e/Q3Xzm+6A3NuotG+5TgGeH69k7Z6bOqo/gS817kyCxqZ
15UCloSjBt7XtZnoCkGraKrrsbGOX76reNhCMOdhLFoVoK1ON4bEF6dlnsSFbwyrLyzpn3rr+IPs
fKHDX6tAgBujQBCh5g3EbEpDGmXh+2aFkMHUPd8OhnI4V2o1l6Ys7WgBiS5YWQhHysNnPu1in4CY
K9tasuF1QhOxy9+jMwM7TnEQPQF/gUrR+4ZGbMSb7HHd1fZ1j5G0UJelgYwAcFpEeXLOA1fraA4R
QD4Dhf+egxh9vUriF7V93gVlHrx92SYTJxxsrUdhYs/mpTR12yJtjE/0VOY8mCSAwYx8fG4kU7ma
3z2ukkMQjQBhGSwDjmSWOocDfAh5/+HCAo8cuAkvilWzgcloMWmmq+xtllDrFWRMUV5O7vY5SKwd
FZGE+wj4hJ0vrrFlCrbIFPNzyPTunJx3Hkys/CWWuVT6PV2UMSJVWaHbI1mJ4dgPDN07WSMd+J23
JqogODU7/0uxpDZxwTBeHtBG2H8mSlKlHtHgUuHGGaFqKdoTqY0zyad1y8u3I9AovCfUqEOMWKE+
1VqPOKYVQqLNswUzuoI8wrBxcNGIWEEeaTKyajxnv8xSkPym2PIed8eNNyPdJpAQMWfRY7w8ihOv
GOZfGpX+SOq5Eqr6Y2htU3l/BOevyYF6+Oie5MQD6Uxsc45XY5MPkwbgI2aNqqpl0Z3h8yK4kIns
CvB/l3imVPTSlB1Ral9vlHhjnpl47ksAVT0j0OdfwmLheq2zTzTrSuxpfxtACwaLyoaG5lrWHLju
9ORuzYjTzBeFrIP4tqLVkbDy2PXPi5McoLPECGoRq9RiLel0GZUAtqqsiPok04pi0FeUZq/7WYYO
aTbP5mFHRaKIvcdTZ5k0CH+5QeX2AeZpUzjaROwFUCiS8cz0RScedaAsWVNx2HzYviCxjPpqCOT+
EDWv3ItJ2EJehali7EjdZJJG3FjVzizwTGAWSbtlFOEaf3LAU7WmieOCRPUOMw4UYlslyr/y/IGX
16Zq3QEW1rh1oisb7IWza3eqMCmkVlHrz/1DEkCMcjNJ53d+MrZcDqslX4cEg68gp4TrVC9l2gT4
06vRawVecCn7omZrb3pYWa7uutZU7BMabFAbLasskQBgnGYw/oYAIp67zfJfLPdHaHhf1tkzrgyf
oj4LBRrbrXN20UwZ7n6+D31N5V6HTDFDfj/dY82itsUEPY2R309p1odGyd1At/HwXC8aoIWsOH5N
faNKGjX1/8mml3e1UD3981Yz6TzuydFAjZmt75BJ6eJv4QyjFIra0pX0ienZmvJgaM4g1AEOBAwu
PnCKwAaNx1rH5wdiFMp0QjnuzWT0M68uy0P/KSDpg/Al7lTbDUNEtlTCfQ9sxDKek0uAnbLvUbiG
MNImsCoFrbAir5Xcl/xRdw/AZVyW6IHZiMdzGhNIHasqyerqXSF89ch7r5rZDAkq4rEdlNaEpGtQ
2XWrQzqsDJGe7Sz7lFmEDxKHbbslMb5HsQ1m5Wv5s+xbbqFfMql6LGKCjV99ooBy7ny1QUwviWDJ
Sib0KpF0Rm4xEjkLS73+ECxRYXU+joOS2C85xjL23D7rSb82SyXM7zRqtyiKYvrK01OV12PpN9Wn
dYpjFpmuA63zqwJYBPS8JWiJTPVgWdLysF1wUOriwWD6M2vJQFct29Q1T+fisFabfQVSYE6qnAhK
9NewVYoFGTDGN6VIdrs5jrs4uJqxajqj2IUFUiIZH9XP8O/kDWbzWOoOuM6S9YSuRDAVeXkrxsOc
cB4FAsDA0r8sxj6VykvXMo/FdcyQSHu+AHGxdtiUQaVyT6uctNXgj1J3fkq4ueqYNvTdOR16FN5L
EuWEpZmGl46MhScCbG0OE8eH6E9HTptQd0n+1+/n5QX05XMNKA3y65VGyrlyxwJZ5jAw//RdYahR
wS0sinCsjgFo09v38D0GrwSawgMRSfG94R1UH0rf0D6lgzyhfurK051jpaletQ4zgkh8x/wfksZJ
3ZP0qtmZqfCUrQ1lW/BNxZMDorBZ2hr6bUHvYp5dgQDRZfivHvNdS0EYPrhKGYU42qrD0CvarK5l
kLkR5IWN6JvLbGY/gTUjeqpcEmHneJfebxICDPLwcujfCyzxKZfXeT4SsKdp/Cl4yZQNJbFPSUp0
Lv5AVSKy/PwPvsMjoR7oh61RGti596OjN9ZZRy/rH8p5T2bjM5+fjNnExH699jiNVPrrbNxphVVN
IyM6gpTqTfKrRDMcIIHTvJm4tTfYk/nKtCLzsHpJnazGzaPhQRfh4KsR2YlcI5u45H/L2a3E/YVJ
KdS/BzPvX/F3P4R3lBXdMVFHOKxOApSbEJCck9myND6MZyXAFDcA5lt7TJnfQdPMTM90l4FdXwQn
2T+gtjriVMQLNGEHaZe3ENRYEnUviYYAAienIMLIRWYc2B8Zcbz2iNNg5OuDf/kUoLpUHWlWlXXW
vNr7xIQo4fL3YHN3qq9+FkWGCeZfVub/k1t/pg9LboBkyc4CgaJ1zB+rO9B+8WWx1lJfrl31zvMF
0c+fenTm0kTHXMb+Vo2zI3Gs7RcvGltFcrLipsWWmcw9pOI+rfFAsD9wr2/MJuZyrsJo5DiZVgQX
2RyWFKYA3y4yb/p22uGvWtGXAVINscJCtsXfjqqelxNqWgciEbavVARUhRrue9c0jPV5D0xS+Yy1
FilSG3u/L9F/NOKMtXo1VXDu05+LElYEgeEUETNSnOfx65eJfWQPRluDjPD7ljK+A4m+59ClP+TZ
p+AzHPe94hIrt1GJpFQ6BhFxNkqAdFVIRCY7GqEeMW7jAXhQW3m9lrZSJZWTLtVJ/J9mfBpW97iw
ZCH2G17Y5UJkl/dWqQy5be3g+jpP3BC1D1dHN+R5WErXguDTJcrsMsHtoeszXkzYepJtHznNCB50
36+aeGgBro1AvKCbJ1bQE7O54tE8eXSqkUkxlst7C260/iyp0YDj5NoVeOncvuOcBpqPpQOLkPNZ
LQwPG/BeAWXyzL2WVvoDlzH4r6SJNiL45vfQC+ULbH+9YFC1vy7OxwyyRQFxrk/vEqyn2Ffoh3Y5
1RngqGBqZs+tkRgPvdXCmvQu0thlL938f1aJIvX2+9ejrGRbth73S5H1NabkoMuKYJV21lLUV2u0
oByz7PAq5N50IfaROzuV/psrBsxTixkgEZkd2WxKlUETJMW3SMBMMeEqLl6vRQfpnTTXf2Ai+SLr
U796C3IVv5Zb1N/BZhBd7vJWl8u/V+R4cTs8g8H8W1XOuhZAcP+2PgML8CiMu+3Gued6DoglKe1h
Rlvdw9+mFtYhUAzyg0wH+Pn0j4Ub9o7oDM7giK5UUG4YEMS3LA8hXXrzYik9T3GjcPp/pbiYMbo8
Xq2H8b/0FSG7XFO/UAk/mbHC9ZWk1QehYONGGaDW12qv06qoHgULZ7u1BBkXXR2v7xgwwZn2bqg3
1dR+KuNa3tSga0/HU3u+ZnnlGQlbtizuDPdM2HDLMZpYZ9Sy2sXxJrqb0PaGZwRDo4bk2BkVsp/J
JBdLnW2Q9UYl22OQzRP76P6PjJPSYthf6G4LSqPcg+KK9uGxgonRPmJsS69DqKsozPPde+eAFNd9
1IHh+UoElCRzj6pulW92AivjuE6xJraDwsT2T0d+SfxiZSHrW+g2Ez2mDWg6T46qoNwt1JGkCjRA
ejTsid9Mp2VLFZy4twMPh8nAGhlxN1qXOyhF2CukiJsQgw9LqKjotUrFhDlxePbGm6tOIfoQ6pDC
7kdfruLBSe5iM262pBLp8vJMSH1afgadp3M5sFyoBDQ2Rwt0mKeqchpcVTUVbq+cVFd+8Pf52HHC
TRFeKGA5QDIOts244CNsBnAsSNSXjOA9tonB6IjRC6bU1b1ixl50SAJoU1sPJkE6jm2UjK6ubs0w
nvCbvyaXkeGK8501jyQkQAJ5bldsI6MfD70slCh68OiXAsBJOdzeJhQ7xomQJd3La/fC5P29hAfg
J0VKnEoEpfr0hRJO1M2ZKBOVLDpmRbSQrpx2dLxFzXRHRVKzSuUOSaG8tr1rmMDDdSqxaYWhpPd+
w+0c1LtjZSP/+keRcd7YFx5D29I/TwQx3DjP73IBRY9qPedRRqNNQlom/krp5LgpvYE4W2e/XpPm
v2Fxrk/R/H56+x6ZIvpXOzM0bBiOOSM8PAfx65OzThTxWtEyaL5qz6o7tYJz4UYf9zLD3nPqs9I4
OM9Qc8rM38FZQFaGO4nLZtHxzx8556He2g4eaofCQMhrUbQsoV6LqTUmu5xgV89AgxQku63xmq+z
2Py0ZtKB3RXan6ZmChIg05a6MU6B29cGFXz6LCjzsehDwVxtSCV3y30hfXUVkNw8x8KM/6YZOiIc
Pj/eTagCgzkK4RBClLixdABTuDoNnOr4HZa3pZU7cja6Yd8DKosxyxbTx9tJ4Q8+zFjZKhzHvCQ/
RXRT+DWz2k2f8//q0yR9vzFVuh68PyeoylR6gFg3HhRoHNokQ2qpoW7ZIESQAPXnNh6yHxkpk+NX
BWUjttO+sU52RwOopTdlHVuOQzqH4gqRQ7CF6wCs8dWGTcu+Lj+dm8Wt/Wj6yLfJkr0hHgDvGVcu
MNHzi11gKeV6rVwo42C/M4Y7p66zvI+6dU//WzqgMSEARgRn8MFm1j0kUBYcCGnAvwwjCS54DQCE
p5lDKQgfsxc6AaAam3+z0lCWeMvO3zvaUkOIau5cJLpU5EkVeIb6i+uAoggFhgc3bpbjeC/4VCry
1zRQdY4wbot7zj4S8EV4v7/baCh86kXKqL1iDX7vefwkY4Id3xMdc9b97InpnV+nmoA+YPNjALWA
DXYmxViwIELl+6ICVgAjE34YAFj6PREqxreGY3XmXBX9XLhTlzZIgbj4JHpFBtxiRq7s8+FmYNsN
dYVSy9NVL+ClUWCLL5Js/IJM6XSIgBJM5xZu2b8afOPTdBYdRVflQPjnO9ZXsUWxja6OVqowh6x8
H4IVp2rBSQW1WOgjIz0OptES56crDk/Z3lSwENuhMW6LBKQZYaRmaU0sU956/ODTwXNU9OsOdpqB
sbGuGzxmprrfsw3TQhV/Iu5/711/gilsXrGv4GiR9bigex3yTEZzcjdNUemJ9VdnaAQPdjoZ34Y1
8A8GFR154wxj7pEofWH+Fzm4UExZFcHvJDCPhL4walia8jE4gBjUq7mOX7pBqCbGDZGg3/9gADki
hmV7RGaD3xa4ERZHuUGC51DQQF/Rl+6uesdoEdmXhoJG1dcPVmbgpT6759QI+aHFKoFBo33NZJ20
70gLQPygGvDg9qGa+LE89r0qPZVF8gzifhIr6PFVYhl3cKwRXQNIIRIPe0DxECxYwzrmNXJC1N8v
cxFGXG/ZWy4WSVkxBAHCmNldbb2p1etfcd+aynz7nWqXLgkTOu+bWqWgtt9F+j9mK3RSy2T3qW2a
S7Oy8Jjq/F+psgaJr0CNrN4gc6FE3rI6kf9GFCRCFIwDH+5jOysSrzECD6ZigLDZK1/KwOfyPerY
Jo1i07eobi9MQzAVMD2GogxCQPqObPsSs5sO/OZTSZL2wwQU1WoiIwoKEbz/OJUMNaSHhQHsDGpb
OfFa9mKDVG5mBx9zccGeaC7skbXtM3dkTozHiD5XjZhfkRk8Zodv2MSrKR4P9hc4QA1xdOt/dT8x
jJbj0q6XgbREqqqXnR6W7lXnQ4nGpBDrmOUjVZaHXfxbPXOnJCSA6C6+3oaoeGzvU7OdL7YejXKJ
KGmAXf44qTrFfu9Cf/vYM0t9zDBHi2XTVUZtH2DNVmdLLlYCsjECxBHmXCc472Grp4nkBm3+92Bm
ZFKX/mqqIQyypHI31AD/K/pEHdDpj4TE1Sx/K1MyYz3ESvDOxF0yw0oL0u0XlXeRVjHw3/Oxbwm2
L6AgrbNEL3Arxaeyqm5Rk0V72qNMjTwM+boHiJ5/IrqV/Yrfua1SQH+k5Xy+9rmXFkTjKQLm2ehi
LlE+drt8/wjw+MkBUrtvjTnMl7EJgfIV4Xs1+m8s/V1NeCsR0Fvq+3CTLx1EZV/NaYuRDRQMDspi
kIjrsmg9PY6wuzAAlqH1ECaPHbDn8LyuA0jEE07adT52RNefyrm3OkydN0yD3HwrPlrj+NhRzZpl
gug0e8ajTWWb9tH/1qThWUGgdgF31NN1rR7mCtyIexOAlzbXapZHNQW8knsaoPlf305SKClWmIs8
fhgRWI2pgwWTHvvhuffn1yoegRI+BkAbphNKBWXvN6Vl6+h5/6myjgYQCoUGzRu4JzkLhL78e1z+
IuPqik9skn2FFlMJc6cx6ga8t72gV4PxuqDXg9PUbZyo8ttka4sZKgpOdvTOopcBovR7YwWmeYs0
1ew7skstZvOarjxgM5HlkiIQ7B8Idg1dz+kfm+EIGa8zSFqMzdX32hmgWbA3Pu+0HiocqzoXVSP1
oyB//KKM25hyN4IPfge/qdecTIWNHfp8HqzSsIsI3tLBa49EXTIG6MxPtinaBIS/FnN9Yi7a112f
aS9CZNd1ez+gO5Ev0WHMgRCz1G9f9XRG1xxiYqGhnAcPl+UjWkMZbw2EpOlfcV7E4H+2+UYDwqPD
qfkq6dMlVMzca1nIxFKnthybezcAwzuTCxJbfdiOGZIW5MxAA40t8OgfvUmd1AYTcwhaiKcMQbOU
JI33BQEh0o5ZrSLZq8vMYPw68hvHBhokK5I2kY7aiuuZQ9FzaonhbZzB+U98MdOO+W4oeH+lXO+c
CdJbzevr1f+T+N6FFQz7udiCq25fN++PrvUXJxpt1C688iOGGMIAA2aLoNcWF3RupK605/2HaVZZ
e5jt+zRxu9Dn5fZdYtzAOAOP7w4OQAqQVZZ+0FowQhGxUVLhoK/juRYFETLk0PxRHQ/HI8+AhWMA
8Q7sexBhC7hAxsOc/HnRoQVPSWd3yy1WqY2S5JLatS4ZgT9qDl+Zq3YSfNokDS5fBEL5+Mcf2+5p
zFeJmRaVJWyGJyDXmwdVNThufoCWYcm2l8F0+cidJIL3SF5q3V22gzZ+3zAsaH0OBap6c/sy0Npn
BQ0OeYLlKNxq/FClyIMR4jOhEOQmwtVBxw39N7/uNRZ7XBKUzFTyXMxROKIqYdOBpsBLGb+xz+JI
5CoSfKJmOczTVl3uYy1j04OzIA8wIyqAT2wQOOrNO7lakC2ChFOfvmyvO4n7GjaOC21THYsrGqm4
1v0Xjc61tcXJKmmsPmyukq3KLFOx+8nAYCIRr0+2HwsiTu+BPIy6ZCgQLOwrnzXXk/VfPq5ZBqM2
KSJkNP8wd9JcUO7RWr+mirt8THSvoaHU+g2JVjNwnFybrgsdsGj4Z6gtdubdT9ac0r4kMrxct+dT
RTMtW7eRKrpZEPKADbLRWlEJ3q88MTifHWdC7aI9n3Ac8j+8ke2TEV2AO29O0ml/brrGjZN4tLa3
ScxqlSUZTTjTtOkQt4p0jZMCGdtZP9YYXwbOkHfTn7W6zG1wM747cevhD/hOh6eVx7gIres3Sfv9
jCH4/ftAv663Jhn+0MV8JQovqhc9iLqfb+ZUEdI9FT9YAPotSXUuvmUmUTYiXYkn8X5+4mYZf5na
RqbHh61Y2kyutv28Q4m9Kp3uIYTlIRNy+a9cEBaBZkBXLeyLwAWT4Fh+//1S+0GajlUVHyxz4lL0
uCPoP2qk+SOXUm+Y81UH7rSBGKq3nURfUTtYXUPA2ga8ukkiBMo1ydQFvKJJxrpzJ+C7FlufIlhb
LwZ9ybc9gLAEybbtOLoOmVCul7VfiF+A7EmqfLq4BlJ6RDQF+T/lTHkoexIVdz4rFq2+UJMjB8R9
oOG2cAQGNeOTShWV3rD5E+naCUYKju9JanuAyME+5HcrxyCuvai/fY5daz+bCpRQr30P6iiNnaWt
XcPykiWfm32Ze7UYuvZRC5Xw+/VUyX8VDdMWvUkHCx7UnAVqbBsvNRiRFh6TBnbmypNnQ1/bxlkV
Xgu2C7LnikJYJzkEqYsAjth+mlRRLDA+6A7f3BdujI3nt/lyJY+MpRSLOpN4pUw6ZS2DdOWSYW4W
ctlE52ByyNVNjoxwJmKFtt/1MxOVP2EXVg55LazQ2BrZITTA/ostxUurVYw9MD0DpHHKFVcIt/Jz
HyQxZszuVBQVRnOspuNTGXJsg/DEP6/69nNKPdD3KtBZMhM3MG8h6PAQwm5xL1nWg6KylPVSLvDw
TI37wCFR0tzbf0Ys7PvIRMjAsOOqb1kLdS47cB/IZxtkt3ty0ntF1+9KiXczH3LIExFuM0jcet8r
KhNzGN93lRDBxNB7kPWv/UlUFcaSUr9G5vVeYGvTXg8i1q/PoaDiso3GmBOMNrGqVtViVMhbxdZX
Hr1pnI+y9Itv+UjbJwOxEPa8I13Tgjo1YD8J0xz8QHO0ISHOMF1PWfaMsOuBvHiB3yFHVlTkWaSj
ZFJLRbatiWHHAXQLd8zxe6Y45fWT2jIuf1VHklovKiCxKhreIJOlETYNdz8Sw4laHivjSrxmqbnz
hvcOOaZkyxzxExpd2kt7SyKktn1SYpS/62DHLVsaKWvmh5CGuBqYUHugzFTlGitNcIoC13f1IEgv
GbqhmIyyb+25kwVO9NsllR20/m+9dFYcknfkgsBnCsb7bX9I4h81hUtviuvpQ8aYUOUfi2nVQAab
X93DcZ38T1ib9N1j0wAIV0z0b/sYS/HGULsF3V+JE+BCNAW0Is1E9IgV6HNpw8RvR/aceirptOxV
C1Y8bNz/+JUvODiOJWS78hAHiCsDRQ/j0Tr5OsB817xWao81BZvyCwt+MVi/cdkscsNL38PC8HpB
pLHojQU0ay/d+gneYd8cQ8CCf7cUwI7qgw9WMICVtew3s2rawvpOFAsmf7nFdMsGBzJCNpQf6riq
DjYajosTlCH+bKvXfKk+4Wg8YhgiOFncSwbP5OmYYCaokoIcDHWrQwWc4CjRIhnMAkGihTEuWJk1
sN+emCAyH1EeTEzowb7X/CjUoWeYAKTk7BnmCJ35+no6JnWdhmvvbn0ASo3W8l7RPyYPM2+/nYnP
B5B0y0rVrQOcSsxz2vk4EtzScxCMVvTnPlf4mgi5+t1MzuWcRGQ3vJp7gYgO736qvyE3B+tnEV/c
SfqKHN/bCe+sSJ4AaLjB9We9GB9C0eUEuhZvClGrCT7RjzMfiAX/8fmnAAs6qPuG1rt0t1tMNoEJ
/C58iBwbDTkgR9OOYQwrxzvhjs5k2b2aznZNvjk4vwIx5j347ZUy0HCrunjSEPfNK7Jredke+AcD
z1B3usC+zTrOuHm8ruPn97jCiBxgXst85/4ks0jRjMdXYdEhQsXW0Ygvzllgc30Yw3jRDDDJ2xql
xPnVuc6lTuT2U2u87VHF4AYUZzjeW6CPj6EOJq518KvjU2Mdk6/QS4bNhhS3IrdEutdDqvpd3l+G
1w9Yq9YiwpAQjwETjH9s0baj7lQc5dJ+phSRGdp04OYwemD0LTooraaS4rVbXSgYFGOMuk5F0rcK
Fzcyd/YgyquKX0GDQ+GJuZYjJo/+/ksz86xhX/U9pOTetgadQl140V/sqXmEOsxSHNvkymW8n8KA
cO/4WfskCTQh3OgZUDViGsx/b8a5h0+nIXeCf2Qkz3z++sOVYt+MKv569Dg45QNXI6bMWDAkUkH1
sEm1FOhIsteC7fPkm1DjiI7gQd4miSzX7vS4CV9EW3Ql5Egz0y+70BsVAi5miTIISWTQ77Z9/wsm
kLvMT6cZlShBY/7VoNNF2zH7DAr1k+E5EAzGNDeytheI5c5JT3HCRUdEauRzh7jAAg+ETDtv0Ise
bR0TtgYMVlfwSxDGCaXjHWlve40QDosZc2KTbsIBMCLwPgYw6tx+45Danlyl9PYK3J5UkpSdqJ5n
/t6CpUp0LS3PxDPhxJabW3H/SwP/tmFSRYDaRIAHtYnBj+PwbnidM2ILL8HQESmBob+6GryfvF1Q
3EeqjyA5FbkdG8BeNy1w/Y+yD91p46VCYJkVPLv9Tk2WI+LRfV7WJkmCIMa1m9DututUF5K8/4W5
w+tU0XoJ0ND+4sgKMVwCDUWtdXvLJ56Cb+wET++RqbhlCZ4l6Jg0gKiFEX9iiMHv3u08tdbImQ5C
MykglAumYtkomMtpKXCobYU7XMT1M3mHSQs4i8Opxjve0GZOWjnsiVCTob0/8Rqzhe5y4vPpvym0
5FZBF945nGEcNIMsT+UomFcrjZqHWLCMhvkT+vnzNbhTn+CgmihXkukUzK0k6UP04lPaN0AYE9Os
lu2QOPEos1mi1Nr4FMvw8SGBxL9KfIV9IaIGcwvrpF3Qd1a4gLvTAHjLD4V90SaDQ8paqROWjKEV
MBGoptM4oHm1/noeGWj1fquft3fRv9BCZmxQo5nXT/yLoq2dZpKiY5eXkthgL9GLZST9UJjfsZRP
tvCYCsFBiEeE1fEKrDT8KZ8fSFDFQacRXYbESchB7buJ6vVmJmgNZ1QYM1mLaXwHihNvMMiP8Ok/
v7aQu2OIEXfnPL5uJsaRbDNMVawDh18qVByeq5bWbDhSP5u/n4a82Re99aDYt5vKQFl38zn2jKUM
FgVJm6Fg4csYsdtje/LgKE+9SabgZtR2Zmoqnz3orVnCv7aZNVrKzO2HqDc7EuZvra0Mau3IQVj/
biTI+l1i4OR5jy4YN/C9Gcp5tPLB0ciAh5mYZCG1zxcEBZxsGEtZvcUei/+ZkMWuWh2va74roBvc
Mh9p+WeRUqGZxcNPLd89pFo0QZyC/9GX23xrVLAvX7xAitprRqQ0sfkGjTBr164E6a3I7jgvlGrL
bTHArBExbGawMAGjotJMTLZyqtJANs8FAkQw76lXL3B72CJYrMeu01130SWN8EF06ioxy7wLHwDs
XZ9Xxu9VteQLAMLjpJYZoKrsbR1Ik+0uVaYgDLP+oqfmo1RfJVVNnpXKiRAIO9bdkV1xIxRooQST
5C1I6rMhI/qsVBANXhypwyHUNrU0RV3KHJXuwC1/T0iQhzLPd4q7fd7xWc0dZ3IzjAUWbwoYvCUm
X1LMvPqmeZa8i+8rSDRxO+R92j3HF1Eu8mRlNKuYZb2t4v9UOPcvKNWwd6Yf/ovIePt3LxoQvwYX
J6pVJWoRQNyvbxaV3KMFiOGG+LufoNdxDSw3MQepSHBZtduftVYlxEErRG7i7F7abyNwHI8br/Go
mc+/qcV4xKDcKEDl1EtM6W3wGy8omKZbNLtTRgxWMYCjg7djWrpdxvYbEXrxBKvOqGiOP7Akoz7H
E98j2lRcU3fe3PbnR4jLFHPdVXVxBqDXKZ+S5c2awEeUtxnq1zs7zJBr1w0GcdJG4hLeMXlxmBIH
/DohCzCLv64jnC1OR9gTrpifNSLGvhuPUSysWb6uWnp4gfNPGaDQqsWCq3H4W3eEelYb1n5cjNPo
06mGegjP1eeFPE6D+T9i4v5oRJ8xDoDJtFWJT0XVlqwjxAO0LL/oT/X4U1ykVdneOJXU141UksuF
1l3driTU0wJq6a1TxrpB2Fit7HgnC4HSV8IQ9YdOJtdV1plwMyVgOD5R4obcbsyOrYEnx8u8Qpjc
kBFEPjaQUz4jfFoXjj9QKrhxOIU1QT0vKADHyZVd0KV62QTm0K87R9a6OCeF9Cx8v06EsjTOHL2u
uvM8w+8LEMKJzZIyDTn71MMP/rKRjTJU1wJMUwdJK/ojuRUDzTuI5mvPZ+B7divkZZZHx6yWpXBF
vV6wI7s9NJOAlC/lmr+cYV4qx2eCAe9r3UokTbRg8N2Y82qT7iVjSlwhCapm+QaZbYe77ZNKcvUv
9L0EZCgxmApvBh/UpBFdKDa25WgheIlhGWSPXs14YmhRdN33DkqBrZaytrYRbWeKHwT0A8hJEjgR
caQsJW9oLBzVAiB8xji8fFFTLTuu68eeea/9ugn3VhcyO+wT7jhplgGxB4BZC1vzbgOtDm9RTLFR
XcYyQBNoopPKH+1hgeWDRUuyPgoN3Vatsk6z9kihV+BxpK2JjxAJPn20hZN8BZ50ZA8eHrAUDSCR
W0BC7+lcXDH93MUBEdlv7BKrEHV8l94qVZ1Kxb6nbxbiJmviscW2f0umnyL2mn3u+VrtL+BNb1Se
PDLO+9ALBqZ+wCoWvLSj4uhIQ545XjpTDWMC+HQJZvnK/pcl4TVPWZoCoYz/y9abHRf/SdIiETr2
cCpXh0aitxbVilaDUaisReu7iqp3OjfBrj7JRVHzB0SsPYrVth5kRAVoYz2L+nrrjwtWndo6gQrj
zjAGc/RjyzRyk9+LGzuiGb8liHFhYNFTDH484jVnAZ3jQRxa6IFphF6DXwXTpJpcZvou6PAoIByA
9m/yHDduExad77EiQmG56ndTtN1ge2xh9PbsI86WFS3x0i0oQGr35cYR/oQVdWLeoz1SNduvSBN0
x4CEPIXBOYqGt1dzlGNR/uSqG11K7CV+WaGN6Gbp6kkDljjV4iVtT6Ppp18Bj2n2zzSKU6TNmn9f
F86QgPrFvB0TVTCVtPDPdQ5B43OqTybT7RFWbrj6lOdPyCEa6NR2wxF1HSS7viF1M6fmi27kSsX7
QdzU7F6Kr5wiNXbfVub+ozVjDOHhmzMGOzkGV3cUYMnx9/MKDWvuA2YUugUIz7ISDhsw1Sxr+NFT
Sw6G1iBM4b1tnp/EuQWgkyYI/XOE7h2d+Pa+XTVwjNOsvh9ZwFdeV4CgH+9DwdD3jM1SMAfjWVlE
2cMBDmAhS7rLkIIJtvEqGv07P0tMFsgixtXgPkd9DNwOq/TUaPbnEDfkmIgWhKGS6U3NlNtzL3co
T7G6pPr19W5jdVbrzZFoPqv/gGxwMHfCjt+j65Iel3zBgsMguOqJzcsgM3RzZ1YXfqP1tSvvK8Lw
rL7UK62H+JvCAIKtnxWD8C14Xa/qFOCfm+jsICFhWh459WqyrNc4sg3OH6SdERt4CzFxH3NObzy9
cHK+GElWnV4pf6N4M9pY5WXrH04DmTzw1J/XLa3bNu7O9zprNgHw0cI5HzPxC32+twkClC9GK7WU
2fkWRH4o7eBKKmDloEWVAan+m/AJHwwuxlwB2hWnjfWnz5u29hBuVk/p3OPgJPHWj777b82TH6HL
5EWjhTnyfDL1pmSg4Rp0UNfvK3rLXXVbRhGLusV0PDjVmIoVw2M9xldTcie4Msi9dyn3YlH+lRbH
nL9FVAMCnYCsRx5uAlAp1yw0eWPvGlk+uSif4Rvaa4B/szfbWhhDUuQjN+wFdsPQBn1pWIZX5Wlz
/WvWNmw1L+NSDPzoBLpcUwlHhHv9Fhd2OsLnE5wTG2+kUAWytswNjJBq7ztpMSRysTVfmA/cpX4V
pXsBXcqaRCGWU0z625KbVEjgc+KDK1R0m6NSkPGAgC17w9iL1vsfE8IIWlJq2o7bHeFY7jKHy8S9
XagV1wCbJ/iVszqWzpkLeonB+1bpYU9blBe5SyKknXgRfm7qXzIyhOvXNBf9RrSD6F9n3TXTyrbP
NW6StQEKwnS4EXp891VK7Dr92m7llg+u34UP0mjpeXxrsEg58KNO0xFkT1tRTLuKF7sX2vBe8vjB
0WlYYiJPBIt73QdHpfmF/h0GX38pV5lgrrXRbH0db+mRQW5HTLG0W328ieADHeE4qhbrl3f4Bux3
4LXFq5rB43CZfwmN9GdBlByafmDyYKO6hY/WBtEJiaxva3LgNfkGpqQd3j+f0v1gu9RvZ//EC7aN
5AjQQqt2xJbMGEH6Wf86pPg1TB/Vptco9pp3x1nxohoQddb1YY7tCP6w18BhmxMdufyJKzjo2+NN
0YEfl6PQ6jb+6ue/NA+t9IYxFlF6EV+q8UjVrZIPBj4a4EEwjz9Uw4pDOf0e2UqU+1+I3m0RUoI5
1Y7zJtr+Gl/ms7dJjHEqk4B127L0g0HqkkFSfcNrWSNQd3WZXf5CUlqr2Rb9AtNOtsx237Ki2wzN
i2cTWM0SSfAa+Yvrgz+5rUsHuWQYqb6p9QLksjBSCYYNjDsneI7GBLM8a8zVB6Fs99wFSI4v2I7e
D9KvAUEy1p/0j8YTBBra6guxdv5p4WCem16r7nrpuP5x1CDzyd8nPSdcSpKhwxJXzvY4c3XyxVAE
9OXDkfrZ8uAYEklQCkHEIFgPmXrKQQNPGnYtytAtonVv0DTTONtVOdPmzS55UTVn0mYhCeEINt2X
GC70qHhlR/6wx7f49DXF9V+1IVC0C9vCnbm1rdycvJsKWurVD3EMGun5cmC4LXpCGZ1O+IWBM4fE
IZEPA5KmnYTWkvyL9zt38FllryaM14zPpSR9EIHvy+iu+OVyE7uVHyY22tDEelwlqYHNfuZ4pCrV
iJ5Zd6DJ1IWBdstsSaVxdkqbcx62NiCCIET/Ze1jgFpyP60ZUIdqmytZsEFJohZbflL28ANT83Br
DkBaI+3WaWlPxk2/fC4kbPhQXwKQX1Vc74M2Mpnj1lMYEbBMQPpEUF/5nY69aH+08VMTbsA5nV3J
fxzdHONKTxPx52VyfYao+3fjN8yNvS0/vt8X2euoXi2aR482OYo7dOG5zTMWR1d9uEeFcAvrbsrp
I7i7kfUoO2EWJwxLOaeY3tT75rZeIm58DYTFaTjTrlORa5kpx4DLPSM3kSgi/x+UQx8LOCBKDZhH
V6jYlGjjPe7Bi2YktLHPJHkSar1KHBB5yKO2C6mBS3JXm6otq2cRg708RhRRwXw54gbr0DIIlIMa
Ys+xb2doh1tkHy0O0OOUVnN5mzwjIo+kxwpvyWPzr+cPiLUbR8rZs7JfCZdQ1ikCVdy3S583NaqK
7yfiYx2drY2/eC2drhr+u3v27Hqwl7FMmH69lgZ2YLQuH9rUaPWdhbydrxyrYOpmeYnedmum7y0a
4fLdL3oKpXTdtFWG7Kc9E9/btiIkOOz+q+WEueanb95Qm52BYBDcpORFmVMeBzPI7+UwwVwOxXpU
HRIZtpUD6hYRC75oEDyF0JmAirMdh04V5DrcpK04892Xz5YTMNHFSRbzSaiLD8pt5c7T99jBAArp
JpXxMqyQDdk+taKw433NKrmwtdYeEGOq7GoSH5dg/XXqop+qwwnkuWzWPXrLaBA3oJaOCLx7ImSh
ty+tPn1Ti3PxrPWfaG/sbQXP+mtMPsiyOanPWb9YwVcHjOFjXN3QZDeWgZlvTekWD/kMVYXCTyYQ
5zp9sfLdVpiIw5sYTBYv2FrNgY8WIdUrDmMmlqPjjfGIVHGPV+tnY4DmSamkE4+1Vv+G4Q8JKl7G
YBh82b0V/9x5qVcSS2sqqXgq2yX5eVKvCrwpz3gCwBVS4su4r6PUnguK/Fxiw4nRrsedN587j6yf
sut0RCU2Tdb+zLAE5+1jKNoKQrqnuQtniZiql8V1u7TcSSyQat0J/8grbqjAIxRCTltBFUXQaB31
C7IoGJbG1pEHvYhVv1IssB/G4EGeR5BjYVjwUvegixxr9jK/JyMfWpxIYfIlNUP1+920JgyNkaEh
KeSGvcWK8ITFrHWq3y8GaiNdUsExtyvK6WoB6Ibkvdpz5gqZitohJcFSHuDExcT3/V7vZmneAq/d
/xu+qlb2hUC02ajVVIelyEDUjxb46esyyPIpnngEJq42NAmmbTXJjJX7Pj3HDNmUnQVgI904faQb
vbzVaFIZxQ8fJozAj+EuNQbo1/TS/Fju0Zbwr6C9wGyzarUb5sYbQTZnDou347e6Idx6riXFMicO
KwI1M1c/7pgvxW5zuXxQ6JxUoNui6zBnM9BSzPPQv9/7HTdsl1/R7AVxXsTzPs3gextPgS0mTaS+
tHylM9rNPwQkpjCfaeaNTBdXjN/tgCuaeYOiX3KXHMS7fsrisbBf5e3lZMvRARk08/AGO2P9aEjv
ZRw6Cl4aQzrNWz2r1vbsFtTaresWtlcfGhhWu5J4tQWM5CIYQP4xTQU8cuwRtyGqg4t41lSvObw9
FkLkFatTUg+exoVTrBV76jFP0hGuQxcvyxnAQl63ATr4FfTHKr7KSWUJvTda7zFFOnJBpfezPZvF
hK82OzpvGKYwu4kbnE42e0M90QqBMb638btLMTk1/3VX0/8tIVFvATai4DaNo/CF9U0PbVCi6yXT
HS6cw58uzRrRHJncPW05idv6jXENlIfG207wey1pIG2Ywhzv3ZLENfsSS1/tROgByA5sbKm31O6K
W7C7KoXFTmNZNMAkfJLBhrY4JfbgxKNV9eJ9me/KzYuMZBJlzjEuoXXhVtkieIqUwppt7OuU9pQR
eOm3h/jY3SW7PhHayQGV2h9h0lRHr0nZDFeW7JL4pNwbTvnUhjVh+xeDLLuoL5l1PbrA3YVjc38Z
nOxnSODHvIqg4g01xEj3TzCACvJxCTASLSiHuS6I7gB5Oht2Y5Gq8jvwFdydx86oUZThiP36DPXf
7wGJi2MZHKLS0LnuN0ulK3ssOH7pnd2IUmN5jgFV60Px5ikZ5KKbYNWBxxIIceFmd98qkdZiGzpY
0qtpPOx3Iw0eUvjv6Oyh5/HBfiheD/22ZhPYIIU3hkVAaRBsRxhR0FI5yOtdmj+8CEoy26WgTQFw
rBsY0IOFyv1iJumMAaO+dDlnRIY0OB/1WnUffwERLcOUCEqgWpS7uQw0iKqhX4KhA1v85QcOl9yr
Ovjpl7vkPy352iFYZxKjTWKpq1mPLajQwlxAHofsNAYhFOZapjqoZKaHkerIbZykXf6NZBq6uHLS
6xDuy1MAzUaDBmRlctdrzo+2Vo3Me34ethkShidAkAlAKpMYqAUTS5FdgKMsxS91csdHE4zemjPy
k3xMzBaknutfomc3uhWfYEzyAz9n1T0zyd4XYpP+hLM2zxWB+Q3JP3/EmptuQEzW7H2zkCxuss2J
SJZlk/FVvAcF/44KBuT6pFV2KrSVf+xTP3M+Vxy4XXZ4u3b1rUra7dP8U26UDKuAm1R/BR44EX6D
v12NxjUY9bQOGyaO8D85KIm/KHBkq3P0gaHjXdYQXK6fiSaXpBRlT2IVH9lRpqZE8mkrv/GnRmSA
dWXSXQN+gKcwPTIehguirLlFr4QzFvsLM5oWfT0l4GIKZ7jhRRzrpYEOOsRFFJPTkweNUmVQzUMd
RPWsh5elLcSnhqcKJOxDFYI+yqO66toLQCbODpW2wU8tVkZFAUNoiLvITs/vWaXGbHvdIQT7sfWk
n3MYBFrUeIoZvO7dpn3XgBVfat8n51d0IBw/RsmHxnHY61IIALVCPZLOcnwjXNWv1vKEm0N2Vvjo
PKOhzqefPFuS1zh0YpL7UmkWhrxlo9vdkl7lS9yf88/xAQtS8jZ2j9zeKgVUNDdkvcGIytlK4o5F
1mhd3TmfpCnpvyJB7BS0bczvWhSEdxVb1mydBfQcVaYGnhWvq17eUnK1dcJuycKi734HvMgQmdZh
XzbRMQHvbFYIGFyF4ySxfM1bf43ljqLauossWb5zt7DL6kOveb2/y73KqXjHTbbhn/2AbwWB25lV
eAAM3KGCNn7MTwzTElukB/cse5rDtM2EfbB238HQAj+m1tvKz9/ZNAsJQ3iK+LORmxwOoBWUdS5Z
YuM0rxdmdHf6ubxtMLv9NXEbMyNs89upsLp/uAdak9DmZusW7T+PyJS72bYtzVoNHAdLxaGvVmnM
SIeU3+QDQzcxJgmfJO7v9DCSTM0Zk5CPSf9cBUIW9LWg3xrgMtSy3eaTHqX3KP8zs2o61dwXYW3F
M5UB5zhXKul/yR3K/I+sbH0i4Cfa+yd9eb5c/FqwqTajZ/5AbZFO6S+b7Jj2CcLP7OPv6U/6Gj/g
TWXYs9WLC3XFGUegOsxjhG0mDBDxpAR6mT1EYsuvEDizatKDQ6FxIF1lV547+54/kDm3gC+SbeNb
RYKZz/RmHQuVJ/PqY038EgDEQJYjfP5rCpFVn6HTqzVQL5FyGMuRta9dKN6MaKhuCa2KQTDmmODe
eJgatKXVZSQWFE2Z35/Acw8sXDPeZtONIHaU0aPJW2amTaGjeFtVpTr5Yt64aFdjTheLy1LEXPGR
ZCgsUoQhkVH1UWAaeGWele+45EWZbnkojBgVODOmR5Ca2amHZuGkFh9wxmI1ewrtgYUYv6GwPFJl
Hnl2l6kX7F/dBnywiWJDYL+j9kkAB3vbi6TKkJgMXwQjYzjqUKgfuiMoS7UUPBfx1fWGja9BQwEA
T3yMYsjeuYd1+8+a6NMX3unGcoot1rGOTxMWBQupm/mpfdJ6+8dS+qeP8MchXFSIgZ4oL/z8m5e6
zMnQbSssnHTlzz1gqn7tZ2i7LZxIfziqG6apDMIiXcBG3IoiUHSTefXwlHmvQ+0HopDWBepqV68Y
Kri1BYxyJ64r/uqgdmrd2kRjHhBBzntbg+gWvTVCw/AWfZtlI9ku1wA6epQdQuX5t8JsWH17t1Db
sz9fywd1ajyXJmriUjNWHtjCECCZWDJ1ezZYK8lr15y4py04vuqspB+TarAF8kOVn3VSEbee4sdV
NAiLr0L6ixinOn28lqMfANn5eAg4QgaBjAQ9La0K6QYAPLcbqdrBvakGdeIqJcHxVhRmtPEUY5wo
Wtu58QMV67CXYYvCP5aUwauVSLS0yTqM2DCmF3mX3hte/TrdYMeixfFx6+W75UQVW3i1L+rpqBin
vch7391+X/gl++KhXRGzUsSv+xSL0XFO5ODwUBQu61jthpoIZ2xdzFDfxfG6V8qn23W3diDRGe4/
jvk50g1MdNygpycxJrD9DMN2yOrDqg4rLI04j0GnFkwoAn/jQmhKgOUCiqDtOXhPa1q71cdAJeb2
ViMKfJM3qda+Ake/5HZx3pO7+vg6p7Wr2bpCpAcvZiH1WNNvJ2JfnYho2oBBSJzDl/hpq8j02CXe
ajBGgFNeJVddXUcc2CX4ynxxC4bUnbi4NRLFi4VHYZoyDgYfKi/JQiJRqIGzl8LuGR+ojAD2N5np
8izfOO7sp0F7cKfPDlZJAlqMpDbuqRL6CbLUk3UGRODK+F/gNGoECl92EfceWZwlqz5K1G1Oj3gR
x7JdkYYqTBj0dT0E3Q1eW6tb19m44vEzgI9vG/bF0QrODFdkHfWRZjxkNXJfpPkVrlHStjLpmXZU
GIn9VYwS2QoeB7Prtdc4nD7j+B7GRPQALU818C7uTnq5diqWg/UhtDQyH1v0JJaohCJDYReYwswg
872R9Zzfhh+EYxx37PK7YFXozosh/MaxnEBWihXP+35p3F9ZAsrfCmioOgtWa4lspXshPk0emUD7
WvgufK7QDT+fNS2zY0Xx/L6MBRJ9bQqEyEJs7EZtJHjHTLSCkPDgtKBNfpO9elUx6nDUpVSXTEpQ
DAxapJMT9DBpJ18QGB7TzF5OI309xeuybDpmq5U/sjVNmmkWxKY7i+6Gd1JdGyaUtwI6TXqPqpuA
Rnh4kvrc9ZQ6aB2WBpZyMIyTZvDl274Rvt5eAtDT3e7P1ZjcsOBQs1taXjAYM9IXCqiz8jr+OMaS
8xd1tfE4ajwx9NVHAqfhTvtzExwlaj/9+RwyOBHqdFgbZ/6mPndTN/Mj1XhgsaZY9IPdS7FzQom7
GW7YJBH4O2UeibM/6wgIjqVNt07IlpJG5zf7bafX+fEhobUb5e3cXHhcfMiaj31jwnULWfGPc4KF
8q3wyj8StcJdManDrguuKZTbC7iJ0e+hVxN61/R5LcawSonvFZzZhQEyUzucVceO+cLECKqRUGi0
jKdNqAeO8GPPIfBVT+NtHTYcyNC44XteYyhUPAS7um0A/u2SeSrtygwTPNccsF5lnSwb/csd5+kT
N3ta1sHjzps0UMy5FMCFsKipwfreFU9rZN5ESvOha9iMZauXiHaogfZtXAfBprItU/mgFe5qE7be
Rohf713C6JhhYRzqIF5FND+HWjV9b+NPKQcg62jtAy2HEMHxAGUxJB8a94OAWnB1Skz1wX98dZXq
jIdLQ40u308XLWVl2Nv5CiFHnGk63EJyioqqkmgBxvbotO1J0T2RK7m/m00oZxOxsDM5AV/vXvCM
vA9cOcmeauMP/8hWH/dNpRZ9LbgWgPQ7u0j79/mksxdLifIdPgJB/pDsqItfQqotZ/swgqOllnzm
/PraCHo7nwFL27L+FxNI8p8+fDwzB1n+8+A+ABgYyxjEfrn/iPvhmnBnlUPFO5ovXksnh615VQ8n
KHGKPMDHaHhFhDOHxFu7igYCjbqTmX8yA/3rIoUZ650u1vJjySyvufacQqMmDZlCgNduiQHO3CTp
8ISplGmG+ChQm6t528+xiofhQhozjj26EoPdGgUoXFOhPUXLodO2Cfln42jAVzweMYBCkjyLyDRQ
jtCDn85vWUdXMr9yKesp7YQN2C66Hzg/+xVe5MPG1TT6FAqTq5WcGjBPdAvfWq7RlAnVMOhijn3B
dJZMLUk/dRbCxwmfpyoYVrqyk+/BEKhk2hZAMZWCAGoGDLOy0m7tFGta+EoauPsvQIFLnGTH+YVX
q4h8vV5zepmcgKLb61v2yHYbqhe5rgKTCmQpEAh6/Wu3ud8b3TmKljwhxOd2gvExW3WBf3AnFUwK
D+JBQakDUqKs90Hvt95BdbCBDelThN8jmElqpknec4htHOdJKdrmOrD3IFSIHrwFLEkvqS9EWuCX
aYim2sObyEwAgAVUUYqLt5yFg3LpVh/S3RrMFD2bPk06cX1uNnO3Vdj2UkDX8A0A/bXIrG9Yg7G0
Tb536SpZ4HezQvpMPxivM6JE00t732MqNNBPDrZbGwO8Yq3RiqrBVos2KANW7Fqjx2CHsZp5ZFFA
NeLRJvtDKDt/m8kMq/4j7lBzNQcvHi0wcJVT5f+mR49ogDLHGChIdmiAn26UBvOnrN0tIW57LSM4
QMeSYrDmT7gNTAm1IrKBJNYKz63lCqpbTfh2TM4rUyTuoV9z+3PysGTw3Zgg4tozbzRj/DoE91pS
C+AVmW2FKik3SjSkPgnpXJGdyGMCa4pG/Q6E1Joaquqmck630Y+w2osWSS5+p0kVy6bd78ukQ+h6
WWZa/kMlNl1gUqo1JDgbvTCudMsFKLj4SMyxKSt+WLE2cflQfwIl5tLLQcuaVdSuH3nzRiirzx4y
YG5pY0kuM6/7oFMXm83wA8mhqHoCgZVAn+yGVvJ4PRk16cFhnSWksOjELwbki2DTXftKwNwlx0A0
/nPLFGCmO/4CL5qdOJD4ySOpaMSUr7SK+HQI/1raipSwfQoyt9kGCLJkgvKxf/6QoH5HT6+iSQ5W
Vd4qi+gm/nkJoxU6IIGaqAITH+noXhah8G7kh68DJU9BRwxRm4VDqX8W1BogPr+W3xi8nRJztbGG
8h2qZj9mxaaW5FRPi6z1G0nRkUOoCurtC+Xm+/6YdbNOa59jcAIbEQRv1GV/SQU9lrtY+v9wgvic
I0uvV5m5gcYu2+fhxoyLMT6F4y/3BDvZ2armeeFb3F7vDLnJ6gqvfVobdqBdC0bEwPIpAVuHsWcI
e/UMPHFrXJmAgUD2L6QjmWfsvIItSuJbLreG0QIPFZV8Fiho8WQaTLT3VLohyOp2dCq2XwDB6KDN
c5eq4AbrXfL7qU/9BkwlnGNtsjyJqGXCsaN6e7YPowhBonhp7VXvxp/G/ZEBAcVHWzoPpWsdIhCS
adxJhMA/pgYZ6XGr/1wk+h7AGDkBZCNonYphHx0YTfJhTP7HjnGk1IH2nxGKkcIMf+y6XCBPjo96
IoNBotz1RxBGaraOaeqvaS9t0EslOfRTMOY/m7l9o+Nn95Yagvqr0hodxC82RfD3L30VH7x+f6eq
O5MMOA9FGx7BpgbjqU9TT+vs8/5It46G5Ol0ZRVaupJS/HssHsS3xypw48af+dalSo+lkYUhNRqP
kucB43p4z7O6137lbNwTp/6kl64tEXpaSlZMXlHPeVZRlGz/W4Wx8zCh2FGa7kmHvcxPjzlxjd38
vy4J8yFIMBsTmgJ64Er0EFwStfn8YA3uFCprWkHH6SdwMKoD7KE8iI/QRh5MAf+BWmRdzqC+PVyI
WUxzpBuQnjuFdeIyDT+rgMXzR+4OsFZn9iLiTzBP1U/SsbRaZHZKaRDxRxO2K5yEWJN+mBofsS8+
ULUZH2xLI0bu3Qfpnh1WnXxq90sEbd+OSa5K8Ip9FOuMZMzioPwFnaN1acarzDvW7y+ODxSxKEau
Bl+xa0S0hHO0yU6pgHBziaonCnxYtia8VIobH5ObhEXkatW53U7l95MqwzBSwKfBvCZsvqSTgapI
Qxf+HOjQoyOhh+zyHLQZqQ4sFppGZ+BVkDcy48nbn6FvU3rZtnhnVx06C77NoLP7HT3rJIEr0YMg
cVE0v4ilxKxm1jNb3fAfnOzzEEBWrl0KM9pYkRLAobJ0HGwxm1T/Pw5ZIIu0d+51RcUyfQ/5zzEg
PMam1+6l0xhesUZZgu8c9sgyuN/BlRSHTJOeubzGZG0bu2PI1ckIRv7r2TOzz8tMP/L55I914mGl
lXGjxLSS26f9HdG3dxO7F028TTa7LI3a8gJ2m9QbMABvj0YAsJtajIPIxwpmcUx2y1j7IpTRxgLw
MWeL+LD1iLen6qx7FXMnMnfbTu3BeiCW79kwiKqQJnZitUxHp1nSTGJsZmQXYfzBX3FodnkFQPS5
GrCY7r6rXVMhbG39cLdPbgTOwYeKOdwqqFwsNvmib3ZT+riRuVTK2i8SZfVN1Qv6mVLGhBN0d//1
N7Mh0AWRC03JH7vh+RXYyPYducJAEegt9oCKkMmFC18GNwmFLtweIy+jkFtCDfsjeR4/AkCR1+oH
bkNw8OOQZqZxmIlq+ushl1SJ+MOTaUYdlebEhosDk/YU/YRR1Qw6tuvTHjIrUMhRGrsazD8kdDBA
KGQcHthUsaiT1W6w/sACOTLuXAL51wkazULg6YQKm1TcWuxt/T0esvHrAR5vseXEBXt96U/gudZu
a1rr7kwbttoARNu2RjkKebgBrVQ4ZX7SrpOJ9eYxKE/8trD8AaAqLfkpRlLb4hR1kG6Xwv4wA1xP
XRK8Z+r5l3xSSZiNrDG+xoCU8KeXrO5OVdvB1UjL+ICqLbBW3mnhSECVQaNQ4vrtrFxSOJYqGW/P
GuLCAE9d//XsU019UJT9HbYyTGSWkyFuJB6cpOAWjYrhnhXW+ugRSuBIPQIZM5p96e7+K1MUA5Yr
vt6eytsc+SuiGXYl+/NAsRb/E6EOnOtqSfWVK7lL8I7kaBM2wTUbCpvDM6GgXUllNA6YZ7zvkEfh
cbmLUO3T2lPxGVo2b9yHTakZio/jb+vYf8PUY6dAzvyhqV0R485K3zPjolamuqSXrPBNH94KH4FZ
eW24qVa4DR+uz4YDyJ1CoMaz9Qm9fpyMO7ItH6C0fq3t3zq6PY9wVd2phrU/WoP9Ev1rOOQlNRtn
IIJb72BmSMrIKiM8E12J1soVN+UQYhS7h3kxNdRx/6EVth+FPPODP65xZPiCIfYvLsoDm1QB4bLF
8WhsClossOyfkogtLW0LHeQLqeclBNmXrihEspMlecQpUZ8nBn27dAQwF+xkqtBbiHAq2j01RJA/
lowSraIN0N4tSPrPx3Q2q6E649dcBCQn51d3Cb0EOlSMzOVFTw0V6gFo+7sxWiYT4ANIV296rzHe
7nKWaWeWs6Pj7yHiQoZwO1UIc1C6enq4cS9ofNozjfGwqe6owQoa8Wkl9L3ly4macLOuSvA4a9AQ
qwV2PTat5tg79JqLSUUFmLT1dnbw9nfeYkCHVQplTi+hClBY9YMxfIeH/woJUsQV+SrMbC9n8MUb
2k/DwwixEye3XVGjX9GYL/uZ9QqdbzYKIICorI7ASo843DlxxsIQH1Dt6yyUZ8pH1ywOjmvPaaai
puOTS3xvPg7FrSWmttqw8NGL2t9ANV91sRXyCpgTu8lS53Nngw8syrchDXyP1xJui9Wnlal6kHYP
TMD+CVyyaPDjpDQ5UIrSxF8uYsvDXtaV+Op+u5O9P+dsLfUe//CB2HP/SqvWjNikUkD9QUB+XfMS
Q9zPcod6BNBtnX42i2mRQKDM6rm9EKxZv2v9TM9CwhvDQz6VxC2qPwI0ipKz2XL8ubNYd5QDNPVH
sXY0pdcDMtaSKJYFSWnsP4tyyZFHc6yaz1U7LbKT8+VvDqaPcflfbmKsu1SY4SCpaR07AUJq7FNU
ZEQ9jl6LLZ6b69juPr7X2FkrdUhgOFWeHFnAMXs52vxNLX91LJz1ht6XNjWoJSXdSPmPnCyBPsb4
nLUn5T0/pMeGVdgtWmBH2xlm7jrbxxTWsvJHpjFNOmjpNiGMsqwjg5D5qb/N/eTo0gAr8G58s3AA
IU5oBCDAYXUobh5wrFuxZuBMH3OpmZ1pFrCN1owkl0FD/bK2VvLahbpRj4um6uKg1duIOzxtqq8T
n5Sr6Q4KDlXiP3n3NScMtsWJlsXtFW5h5bBVIhAZiZdBilgC9COyAAmawTJXihxvfBHQ265w6cWT
JH4t7/za9vowujrNPJtX9jAMdxW8Wl3Z7ETmrrLQiONLlvdARGIeosezTwLXul5qxYoG2kTEXe7d
SRettvi6UwMPJaOJ+LIo/d9JhYrGlrPpIkkGbyFbUxGvurJaUhXG61mz9Pz6q5R32BejHLIgc/EI
ndEOKGzF7PP4RX75nsosxspzB4t8IzsC/e3uY8Et/b+DRV90AxD1RSnV8VxsjnJ5fHUl7468Kg68
kksW80xcKRwEurmOTm2Oawy6SkPhlM0aeSgQjQmDTbPp20twpdddEsrFaZpVFpXAAYoYtwD2jy+5
MPSuUCm4gJodTMnQEX/8+OGVZmIaAIMqd00UPRb71+2JUoJk17+CjpueunvkIaMS6Vfer7t6uIgH
3r6X15ej2OEBxpSFNpuGfU6v2DG4gIbRyeddUWj7A4AuTR3CqvfahkZ/3YsqoBp9GHCm/45UfFPf
7+L6cQNu2pGroZsSPPb6ORtFJsyfgj+OIv3Zg9uUo4/mzvUhvXyLk2dVzCxVUaYxO3oyfb0B1v5h
/r1No5OrIXtDW4/WDQ7Fy/AoDG50BgGZhP5U8L6BrlyIiNkhFGLqqAw3JlDkqtEgfHJkqndgm56/
mZK8k+L9PUUNrqVsyFKB0nw/hspFP9ZCS3ncKl+Bf3YjGn7iawArthFvWwQjalX1HjFi39d0gXwX
zzzwsUM/1n6Fz2R/mnxZlLqGuItjw3MHhMjumjbPpUMGKKpbVgbQJIjz+pzyWAVTYQR4ulzrG10r
quXoti9pprxU+U2oQejD/SxhYxT1EoF+St3IayqAo/oL8w8Cw7DIPL1zOCGwfMfue+RAl8TJVKan
OHgDvY8zaBJDKsJqBNE90/Bj148No47qU8YnZRDjEnTxxziSaWYJVJN6xNfaBtSxXpto3DfvDl/A
Th/rlaVBNnSIodz3/tfgIxc1+3O83cmsnwcCVxx3iMRRgf/mhgjdnNqbRt2niioql5chUff6dG+t
GXzPygIgLIJU5wiJ5XgeWQuAnBJXXFPoKuT+V8U0I2D5MfBWyJ5ES2ZZdZ8Y1DhTBp0YKjQmoKln
n3CYjjQ4KUN88ZsWpNVL5Iqw9bmNQOUX2M1KbT5BHxbYTdNCo3EVobJDHg1/ZgtHG1kTpJ0ZMZxH
UldXy0Iq0mt8Rjpx1eE1V48kKj0Fa9A8NVESuvMp0RupVW3O7HDG9HRg0NZwN4XycIr77DIvMgba
/uaH5dSy28lU6w1UHNytYaGQGbbxeXkhfMHYyEbStGTpRjPFI9kJzuUXRWvmfwF1v/mxF9dekUQP
3n352Pzc0OYsGaXC4kAGdphTFHaV52aGnRgMSZelsBIZqi6/2hJ6p5GiDK1SBr2xglopxgARRp42
yVVeOfsquyiz/sj/r7G3Jo5OzVcL73LIER/P8JLiw9Ysi7ggqtTeAtfQUf5SMBbny6CnXMw9ypTL
lFlEcHsUQxvFy+0K71sUjFx9X+T24uJxFot2/BbHGK1vfsuB2WBJhWIJNbwPFCNHRen60hoCnS9j
gpLtPdz2MhdSJqW8OZ4aZhHpyFKifTgivhwItzlICdDhuoYFml8Z16jdSXb02ajUSwXdnIPdJ2NG
oSu5ktLAZcpOYtWeTK4KkRZR6zimCdKhp0ZyYom3hHB5Kwj8NW+pL2ZzRINUFSPEu/7P18u5P+ZC
b7G9RtvnVYej0symulKwTYdZBPFJmZiBW7YrJlzaW87nfDx76AnoSnqB2jgSS0PMzRnL0VnIWSQ7
lDhVrupjUKoTqY09dNQsSKIFfG33gz8Whph1oAH6D71C8Ra35KrSDbAt81/PjE/654QBcSzjbiMv
YAlAp5HTXm/LH6ggrGZPIe/q0i18n+25deY0wrN2owBSbo5f1QNIev7rwA759FM6ETHgF3UI6Bb2
c0/vZn6OUOW7AWfH3DRzxdah/vuCl9cDsEYWW4Exi7mxhCFT/3iyBz8qE3GeLec4VtEaL5n7hPqS
433ApUirvAMMUVqchru+jmxq7QOp/rkOFOZIi3lF5L0s7v+YDrIPXWpGq4eYkN9vXLWQgCEe87V5
/V8AzAHz2vjNyghlmuIvDEavYwvK54xW722NziX9J5kW/zn+Ygp042nWA9sd7lF447LkQCFzsPzI
+vxKG2bE+6DvMmkrmtN0As+X6BAeGuOlRzqUJZhrXdLqI1rlnJ29KLlCL6J9oy9grLdnEr1IgEe/
4ya+Q6RDFAwZ+Y7lq3Z2dSfxAfaDb1FRAgA9JqbcbW5f41RXpeinAu8PY1hwC9/fbgSFsc3Jl7Fi
2GbN/yanXamktRaGo/XNSYOVZdKAJLR0bERyr6JcQ/IgrZj5NYNFQk1yC8wVnraI2q2dIqQ0bkTB
TL+RGAqYjrGqOBBfrrGuitYj3EXM9ntQ9MevZhL5AXHoSvt0GO+8nl4ol5KUjDDw6WH/XA7kzn5N
SbAho+EqLs9cAAxrhaKtuxWKnovetvDjZEKx00y8KlchoCObFzLTdoRNxrI/7bauJBrIB9saCULd
8gam3mikWELXAjYSXG92kW+AvIcarcDYG0Bvv/SwKR/QEBgWCtEBl6HxXoYikl9EGaUcqsNFMPlC
4f5W7VU9yX0ePQcBpV/zQDMn9IU7qJX728Ev7+QVXxFni3Z3a7TMuAhEMheGbm/Se2pdVzxupkGe
bDr5HT3yNoPTIS8m2LXuJhfBjdfmP/eoc8rw8AD4ezo48RR5VJc9sPsTL1NjU5LxvgCofFsUmM/X
NBD0r8B6OUZpkYsOvZ1UY4JD6Y2z68G2QafGqlYZmzA3OPyFyqPIsTN53tip+W/MTYNM6iIStUVy
++AnWepPDdFcPDXqotZJTdYshARgQOI9Xod9oQgwzmpibXetJfiwuJ/zz6AKn6nTFLx+fWZUNTB1
HwcPf8VEg6SRSfeayWTQ9hXSHVUp2C0jDpTX9AvHgtCxVFBedAD2UUk8skJUXMDxdB74F52gBv+M
bP0sxNAVjUA6PGlO3+VX5sa4tSoZ/i5ONwJm3Lrl+tGGCS/c731jO3Gt8o8ngOfqiMj9jMQat/vc
71jtwODNIyCOMCbKj0E9LRYsieHd2hlAu+IQ7021TnFPRHAmRVfCAcU/UmjZU/DiHlYqJ23g5PyB
h7RHA4o530NSyA2S5GcekDddRL2ABRV+9M3v0zDdNh9js5BkGkeu3MRaxlhaRfUzuiPMBuCO3PXs
X25uRvIz05p5cUkmoiYmN6ouu7h+nu/53T7fr2QLW4kqooaKmyfYR91iC07W+zTJ2WGxkl2pmnDe
yeoL416+dQa3R7KEZUMmTCji+Np5NMq4cdUWi5XOjHlaJGYQpQ2cZ/uIP3iNvbXprPpxxH7EhI3C
98G0q1SZA8SQ9f57Y4icje/Iv0QTO1aiK25vYRupFx5TZ+U6yc34Kxw/XvP4RfbI1v64MQRZWuKx
IlcEOwvTeI4Xxvd7wxknrhJkTBMkMdx1QipWkDr8+ZY1CKWPHZYLA7D8yioSZvnI+viVnk1H+mG9
MaS9NDBDr1xzHNAY8P5KMtHQlVZTtVNQCLGzM2Xri3QY3jVCuZgzkpuH+ugCAeK3cKVR07Vwu77M
LtDa4ksjFiEUe+IsvWDUjTy/DKRKZ0AVEe8PfvhSAXZ+2cFi/8TFsm0SHBD8PZdD2VwQoMjbW3kb
cZ5/Lkvfy4qxirbCFwpQYZyd9CM38BT2OKGRqvnLxOtwUFO+Lkl/v5/DQ6P9Qr+Spgk2oRaJAyMI
1arzH8qSueVvnRm8g09+1XZ2WMEuwfUXWKlL4P0jnLtDXfuVZwVSrXvpGo098ScA+qlaqFN3bNsm
FkOZ12sn8PF25vBlX3iCxRw4J+hX/RsuyoYWvgEiusVEe24b0p3O7tJL905nrkDWjjFDRtzSXUQm
VsifchAM9Bx7pR7AmNEXrleFV2xyTG07csftTE4s6VRza0AKOu6NmULrFyrRfZ157FnmJ0exK8be
NLXdMWVVWeau9ZI/L3fk/zUS74/GpENXDH921m6npxYjGuws4LYXM4kPZSnpZkHNC00lqI4IPoDI
ELsM+ciV3M8l2dzmam6FHc+7loj34FgzP2XOQlDD/OseeUC35UH1rLNpsdoTURbAiYvoxGjKHtIP
1tNucdQOxYZCFtchmaZULvPTNj8F+lOjd61hNVLkXiuCUtriuPKb/0nXZ6JphUgQCpqzOnDZWJ7E
ALOoD+B9HH0urwjrc6NVU6Xz4vDziKLK79PNh992zdJdtRHO7uX++Hm3H3jISS2otIko5BLRGth5
SaEDhCK0Rbd0XX8hZt+Y8pIhxymZ6zbBpr9aJET5GiEO6ps6yJFADrpkgUsdrgt86t6Ys5n0VCVD
Hz0dTiLyB8asw9AYcJMtFYQoXcrApmZo7Xj10H5miDEaWaS3ATONmAALlhzDrEgglRAWjQW4CZls
xO7gnaie9roEFXIn7Yf9o8rDPAXIqKhC25Ll7firYRBNyW8St98847TJ96oB9jTUUFRxH72YsmbB
wz0PH3l0qLjTLWredaHT/54ohGxWJZvCO3y5N8/eSAhRDYOCC3fiAPw33CvlQIPa36pUOE6ViN0Q
IVPk/VwJRGDcbahcDndjEprhg7K3GoinwcvzbpyGavADDfp5n3k2xnYAvFY2huqOuaePclXwWdLj
nUijncNFCoOeJ13faJbPntPZFzNSN357Q4eTG6TLl/f6j+V24m1z7X4gJcoDvrtBpKnpFKqoM864
0fSjvV/emc+6Aab40tB1RdKKv5Fe5TNc+uKlUwmlpkvRP/spVJ2SWvlvKmvOkljcOis10T1MarwF
L06e67NouSbvtSpQei+EKi7AqcQ1j34wfGZfk8t0pjPTQGP/3di4wspKnQrDOBrgZbs+dr2OznZX
rKajkiJ7izlRUPPByZAVJimqV+Fx5Q/673+kLJED6EeOzii7RowmJejenDRpRjtCdI3qWQfMDp7W
Uzb5mt8kdvKgQSsxoDluBOD0v0mzp/WRHYEIuIfp7k6DkZNRDH9TXl41e1aGEslrs0Sy0rHMh6Ut
7374c3vDVK7dkkrlCNGHB0V2wOEI1btZyLAq6R9F63f05SW+zyehSb1cxE/DR8u4uLpfdEy/HTIV
S0UDtRFTc4j0eFGjrsBtz2y1LJOnelq+PYuMfXSRYBXGD/VN8rlJ6cujMurJVCJHP/vvVvf8FQzU
ZfhEvRmiZzFouV4hotmCVL92QramLkukPYx/LSFtAdJIu68XAcNN6q4fZBMEvNiD1rwUzNSgMgie
q28DwngUrZwSfRd0hgZB49s1YdmAzNrlX+ckNULpXs/revWKqZLxsyJ118XMR/cFYDacNbrFB+jE
K0FFIag6fqDAs4zosy//WiZDx35cdEKBQOU6adF6MbXy6viv4Mh5jLYIeXX8NDXYMx48LX3eN1wD
MD9AmRk3Kvxaxgwddsj1s+VpGHmw/kBG0mzCLGrU3PlG9sfs8VhOSrHTXcDuPzZFgreJcdXfyQJC
VY/dC2jB4JvpRVZ1QI7tM+sVfVDLavxGzz9TyKN4ua0m0XN0/mMAJDsGftDwUoOpQ4ctOp+wRrX0
JLUXFdUnUU5NQNKiAKGvSnLWY4++lSvhDQunXsvhGs6tlq2mWxwHKPAnDFx45k2g52CZtwG3kwWA
DHJEExYeYam5Lt46U/H/8hMEADHoMGDK1H44om6CiL25H9CwE+eaTGb1fqVxdoQGpaMQmo5K+rin
gMT0PehYR+N6GmRr/BHsQWnbMsA+nvzALLkhE5UihF5m+N5PQv/2FH9Je+ApyMVRKs0mL1YYKJMt
Y7Q39qtmLMiXHyll+0JInYuq9XNoWpAVVQtm4uM2YOmqy62qDZmks2YozWeYcPIO1J1PgtlFBzht
KHsFFbyW+O++iYpK7nsEEoaT/kON9r8FlMM9a42r4wJlMyry/pqIt2NzbrMne9dUDFB0LwLMuyQB
XFxEj2O24NmqiDy/8ntHA/jeF7df7ZKuY/ISQYKiZy+ZsARXXlFIfXgF5ssYQ3ac0RRiupC+YUc5
e/OgW1f8oInxEtK7vQFkEWGHGlXEqEZfeJMOmU2GUQxfS9EwBqqOo+V9OkYcc+O6r4JqJzDaIMhG
Sy0jKUq1QQOhA31zYR+fNH09e1s2SM6NC8H1lZ3cf7lmWkPo8rXr3k5Vo/TluTZ8YqXZ13pJeeI6
PyF9qATQP7kwbK6+qJnXoGQrkMVQdirxEbQ2rHlvCorwLRAmahZJzGm6WBNojI+1xvT3G74ltUih
m6rmib00JOyzMxFv0WwXBgctO/K7uQSgRzmnMT8Ant9yVONmWqlJE20T7FPy98x9T2bz9Nq7SSlm
nZsD5cXa6tEJS3dP2d2vAM/G0ZThNYj/8iwYJXs4V+xSw67f/S49hBO2xI3geYSmukKXqdVNf1b3
0E7d/zCJVYtMoXZhwFwZrBBdEE0WwRi0Vb/7R2Ps4aqjR/9X19i9+TcyUkQFR6oBHiv1j08itgtJ
cgaPgu/n2EsreRo9iL+QH6ZDFN8kgeKWGQz81XMvBPiOBFnWigaOkWBJ6SL4n4S5mte7jzoI3Jv1
ZOAu5XGM6E3tm4SQuqTjXZ97O3bI75H0LYYy6FgnyQ91nYzNKbLXI9LRGRqeZzDJVZAJtmUVhwMf
GXV1c763GxQIHqPsVRj9SIrFUljFuSj+aubq8mf1miiUftlrDWGqoUclgbRcJhtkyLatCSqEf8KY
Aywh3QQFEBoq5pGFaIk3Y/+tgwQ9VZR4W5NkDFT7sSTnTVmqsm4bW3Uhxq52TQQXrgrR9pCQTnRF
dEf8o2EBMPEjsAw/+LHeuStJLb8Z5DAOhZ0lGDq07eU6JMMa+ADFzr3szzLrTBZbhlGMhxSweJq8
KYI74ZLHct9ZZr03PIyUYkW1xTWLPHBSXI7FY74c3SaHVeD3yOJfSnxvHs9ASZuMpaLGphzmQLvh
uCNNFsjt1IT/7hVZt6jhUoEpx+jQFsYfm6u2OZtb621ndOY0sFvIAZiGxcoj9uSiTNpjjh63OvR4
jgRBi/yQ0Bb9HvdfwtJrv4agDvOtV1vMYvNaohh0+ShrmjpC6/TIBr12FEzg3GL9KM9KDnCKWWve
fCB7mhKkXTZ6L2e4SmRyR+R4zrv6FEe4h5v1SscWJI3IHVbrs73oqPqLwkTRd8n7fU0RFrfaks4v
Dqi77mBZgcF6Oj61u33YmmEGWdnpnbTiOTOX1OhIX1+PQUoZa2V8gLU1NvtLqMJMTfuyl61MJ93q
e4V8xtdjPBdHlvRFaZUcc5HBlTnyZLULNZ3xKE0alPvcSYMescesZ1th4VF+Imf9PKxRsLCbMEkt
dFCzbd0w4jpGoXhnd1iYkzu6a4b8igiYiM6VAbNu4OPEq9Fmg6cp//9h9gb4pa6YSJcS2gxNy/Cn
tPkUbNkqLEExTA4v6yWYSuLUxvQtYDXYm4k3NFfyJUwdGR5wTM7qWE87mLMSR47iK+DOjYC45ChW
hoq2BFl9GLGvDqQOKBvQyao4kGZdl5IQejqi48MmRZNEB3hpDWdbuOS8vRFPEKaX/wcONYALj1ur
UYtQVrCQrNf4d8uHknoixdCLorUAqP5C6ID9PMKPsKQvTEIQy6ElGHiBV5Qdj9SBimycefxwxB3u
k0E6XrVAuepm/lLN7qcRle1wDJw2iXBRtnlbg8uwZwsX1P5jJZaT4bxrN7RzuesdAzrjvSCkOQeZ
kT2JAQsMdhEL2JgIIR+cvYFH/DsZfWAR9N92aeiYnDJUSRJsI4459AA4ARmBCqr6dgjXG31tNgWb
L/7GDMJPv3jzlpxXNI8VOjqxzt5zYXRvkSl/OPl4QoNmczaNRZGcntCgWYvdx3z2AvJk2sQMQqTx
CIiE1vrAuz2F9pRRIuj8zXDvWCQHMR5WzhvztH0IRrlIJm7CB+bRXsU/FmNPWzLpGhatpnXvvrZk
aXPhoDFxOebt5d6nWJMjSmSBayC/wi03ttQNIcTeuB1Cvf9ZIwJLPZzTCUp8HTA75QBTOERbV8eI
PJkjAmmNOf6bQBZB7aVjkdzkJzI9Sz4MXw0NIAUfvouoIQf8+9k1Rkb8Kb0nWG4KAfTHID3fkzXc
QiV0/ugKbQAhWCQ3jzfRBkPFaOe57gsyTiX17HWj/035gKDYvm5htFk9u7Q43dftjaX4/2ByVRBh
HrZXfO89YB+mCSJcU7cQ3DIo2wAAUBVODsOrG9iftLf9hAOhl3bflRXxo2slhSyWZ/WQcok+z/qm
cEGIjszqJRHQSEkW9H81KXHPnfaRNpSJR/up/5AR9ao9q2pG12DkwWc89h2pPcq1xBkK2ww4P751
XYNzDw+sC51XlxOgdA8HSvu8PdfbPGioO/OgKhD84CNDI+9l8HKhODe/i5QGQYeoZnsK/OnMZK0h
3KyDP1866yh4PdhaJp599Sxy79dbOkU5vy8a6HrqW87SAHU8c2I5q3oz3o2PH36InVtw92tWpsUM
Fz5YAnqYU3AHiFEYkac05dL5sjHa3LimWlyu4aknmrQTGj/Uh3m6IJCzxQv4eBqYmHuBtOXrXICs
wAWLALia7QI5KbC4+roUeOaxzBSKysdXmYBU6Gy2ON0y9I0cAuXXX7jqmgL1KNWe/oHKiUvI3GGl
7RE3lABaO6BmWk79zbvZsIekG+bi9bijR2vr5lx/UzUxgH4ujJVfETsi6lVkhdtGPkLZ0eb8YGBC
H6A/bXXraOb91s8hBH3qU7vRLIM5B90N3p1R2LTPKgRtCFnhIDG5gNLC+9nWx838e/D+hFESxU8d
ncMUXk3u7qpkHIshiFMEQzWJx2oxlMp/HzaoTOdfVwiQV2iNdEcXGh30ci2bs9ek5DHBwbZYIwgI
/ENULdTVeTDwLpnN+7jzziv49fFLr9WblNKfp2bpLmlvuH1ZhHJ34W2qqL9eX1Dc8++Q2CvewcpN
bIX7hELbbqlCi5nCqKgnUIv9Y/KrIPMLCvU+gy0fEqjQkSSbsOQFZ0Z8C2GTFssgPAlrkuXrgmgW
VDsXwViNVok810eCuYjug5htNB6GGwrXfuFgOq1eX95QP0tiObWplMqrjWdTyX4lSPMkuyRwPcq4
XMBLKTNymzYe745e2Q2ZRBTVd8JZURIJ0sNOgfvlhMvTmgvmS7cUQAElx00c92RZAuIJkKcFRgZj
tUV5D3IooEonoxalBKAULoFxA4AOAJ6TRQQfcnIgtpehwthSIpXGtgu0e9TIF56LWoMvbqjeHjTt
IBNPvlQPklMYtYCmiIs2rD+5NSElZlpcrQxdit37BPFXwuHQlkwhw/hbpb45LPuTFm0mt6Up2IXN
XjSiWo9nlK3HJO7h8d1Pz1koQyTFP833JNOKilsWIpTmNuOzZTDux60CcKshRD5PBNELGbaMDU1D
BeJ/C22m/kDkk7aVsgD+axRg5cjOC1Wd7lCNRLp3ct3ca5LEUobiJcEwalmy4oby8MKFHWEkQCoF
GnTNvYynL8kWEcVx1SsoC430fCsOZUk2cNAIW4R9dU7h5JrgPIQvJD2PFNzngBqLkAcSAD2+LEN3
YGJbVYeTweWhG720ZpzxqN4iMac3X5g+368m1pc2ivT1UhgRZvYDfD1AfGZ05BVyTOyMeEZhSI2e
Ape6z0RJRzq96zNZ+l+BxWuhYCsUc0punKzPp5FYMLaDxBGy6HP+5aClLYVRbUoomtWl4LcnDRe2
fAaWKlv0ngWMEYrJN/8y8UB0g8puB9JNE+GZ85MSWFCwqWgnkXi8A4U7uUT6MDQ18SUgjFvUw1Q+
dED5RFGeFkpdsrcmAMOv0LBEqw9FerW0xmAfkdiOFiWS7vIQJDve7O5T4OWmNJpF3RUHMk3Tstu5
EM98svpqmLxH4TT9YRaG05N7QZ+AN3qGqFLA52kIihvnOBDe5gIfCegnqbn9gcEL6vO2qtwlzOg9
/Y47eyzOfaMmrFQ94y5ZypQDbhndlwHxexOTNXUf86l91qhS/gBfkmFDhCwcbBrSMPHo1ekrZvDj
eQgA2lm1SSZfQ3Thc5UHB7O6wGtqw8x3Tp00+0SELeGXupotCrngO7DKfxC7BN27URDmB7m9Mp+t
rmQN8RFU3n+273E8eFNlcRx0lYsN71eDYDJNj7Zhi3I3DG6vA72MVVeShZ4dwdbbTKMkMORTuE7+
5ofKiXFxOUHCQzTJep32xlGTlcHu1FCi3FeYMF1yolxCRHD9K9AzvCDg6M5tDNRyk2ypPdTDEs+K
bSdEJSz9CtbjL80SZNAi8YAispQje5V5rvhM5Fpvey28OQyURcRQSyZyFyc2NFQaif12qkbRxQ1p
ieC4EemDt4r3JlRgkBBiOcmOnwIicqg/uregpOmTp7x+FUew6hIUuNW/nDfY7kgd1A48wQTpj3bD
rcdIOcoFPvLGqtW/lSb97qeRkN1mEn1FZnj9i7P+dhVp4dOpKPTBfHGEi6ePZiqHNi7pZ3k6WC67
6g+aPJQE9rs4OpErLRmIVkN/NSLZfwRmRMnAsjqAKSOc3F7bORLIoquh6uHOAao2vf/4yIvIRdwn
3t4Ni0/pC3gJyA6eYtNZy7PguW8fWIjcU+Q36iJ/2jUBa/tvzsX6rr81v5r1TFEJkC2wvP5zVDIj
MYF8vlKbp06CUa633Xyt7sqwvHIE40ZiBM0PBwkclZ550g53RLx3vMcUddtgm42ofx4KA97DAjH9
Wo6uf0qisGBvSPAWHeaYMjAISy+EEED99DFZqBN26i5/nN5HLnKaS9IBU1XuynYO9aP+Hog/nTV7
qJxIXUkjy2Vklr+EmUrLeYDJKQ2Ea/V67B2+S1hHnCtrfGjhe77Bd7vOrHhlciM2MYqn3bt2LWOr
dlnGu9NohcVhcvyxxefb1TByqSfLpnDLLJx3oxkYWZSOeTGrdsYmPKnP861bEjKQTXK1znfKM6uN
h2e3ScATEsS0jt7PEJnvxj0UWtvv/R8nmNR8frm+eklGev4gVg4adkV/kW2Q4ikbmD0szvEzcVXj
cltmWL0p6X2FiuaI5XnC+VFdJoY6lBAoThBhB1hxSWfeTUJ3DYS5h/HgsBcjdjSgfnSV/8ugZv/c
mYQ4Z3nZevw1r5UPyztDVgSZdNYK2qHq2J7i7H329mY+xJv8rZM2uefl2t9aMdndQamjpJkwtOOR
DBZVdGU3cMruMYFjps8aeKSCbblRhGPK2RHEVF75Y7WOeVugfz1RLjjg3gSNFibl6K1DyBi2b7zt
v1WmE7h6MUs/4iY3UthQEiowxOttwFnyvaHbl1Qlvv22OYOsrP4rtty6sRHmIUOcOsX2Lu2CTov3
ZG8c+ObPZUpMx45krPrEmViz2p66MJOEoba3+QMRQglBHeD6T7OCNGxO5CFjXej/pV6D57QUJhuj
qdJqjh9+e8nJk4V+Ybzkuy83ZBCannubthLADut6bgRY/muzXrtxDkQYX2FsApTFlR3RQXhiMgtY
5BdjSqmZ00JCR76Gp2sMvU4rBNgQtfBYqe25eu0ho3t3zdt3hP9WifH35DFOLrHJ1k2EwyzgdDr+
QYkmaJbw8VbtAYFsXq4eYoM+90v0ta2qvQoHaeuizXFcKq6G3LAlXt9BPIEfakhob/FZcUazS1Pp
l3nNYDGLpynsaqi5FSgcGE6aNQqdiHZd6m8X97Z01aoVYRruke/jvxgsIOJgP55GOACKwT9BUPKa
FZl2q9u8wbxJl0xgmJhUBg78AvN2HgD4kG/vlCenpRZ4t0VC4Wm5kNLqeUTOz/MJMsC//KwOdiPz
SijDp0gKVmH1sQ4/WYosEp3CVhWbBrLuFe7bcSds0SulAWDlP+YEgE/8++y0K1x2dUYykGEgZphh
swQvJOGssIbYtjIT5eKHfhT14OdiuEP5wjEZtO0+INsuvf3Z5GTgLjk6q5t1Unr+lp8p36u4orJU
qFBjnolcCtr4ydO2W2kMhOAw8seiHH2c/FLri1D+G2m35GqPOTex/suGz3c64MBicDx1KzgFmolX
EpdGnpOdvO8wKx97FVTuS3a643G11+Tt7l5tNn1tOVbDVuLo2iOt7lMIEeHUb46xe/7B1huAxvoA
n3FST/X60SFTzr1CRUvtzonxauI6S9HcxxJhXVJ5ZRXT39gk98hPcn6u4Rmv3EZoNL2h6CSTh6UI
FBqg8hahcimuGeV4As5rTY2jejww8RnNDUXnRDOGWiLbMFjjLaOe7KJ3K+ZxtqksP7eg0GzS/W1f
dRRz6JUf2wRljVBr7zQWMTR7fnQGTB4GxTo8oUQ3UuJxkY5aO3oAD0x2QdBBFWDEcxs/iHWAAiRX
NNPWmnxXtmfqhrxu5ghBenue0OytcYlDwOBGJSciFPiazo0kY2UEwQfwwLXx3hgArCSiGAemoE7a
yjsfIuhwKy3poLlyX/gPL0G/enWb85lk64Uj92BcP4TnZ88/nCAXQCEHH2/QxPxCB5sPUjRs/52q
YY9Bziq4aA06MbMNbA7AWQKapRbPRIqZsnJiAXiUq9Q8A74VuCclV6m0K+tLLscRVaUotQG/YCpV
7CAsOfQxeW3lNS6h8013U7gOnVdWmXY5gCYx8uSyUA0b2+g2r19Fy/h7DgEbLIX/PG72x6mUIZNJ
SVdBwTm3VBfLuBBmQaX3Nt/yZwm6+UWrDihMZRsWGZFtjljHKjViKhhBnKRWyCBizunejBcxQvYa
4nzkvKaRxlnuj0rY9VRsN25Pmf92bjfEDPG1azShl5DHNvtlXaFGtx5z8ZzJIZVYPSzC7RlXdFIz
Y0qRd99Qw7c5fYmGhaDuQxTo+kwnC5ScxRfSackZxKniPoEjB47GOkhIGd5I5kxodD/48pcZgMHh
yyohlWluHHDE1YSHNNPXJI3MGzkLDy4awOCT0S/sNoJSG1Ydr3HWPGanU9JQIB0Esbj0njncV1en
FnUpgZCgYX0El9Vu2FAIEfAVqhqf6InThoeR4+bG7TDxhBe2pwyggbrIzRzhwfNCueCeSlSjI3fD
CZWyTlbmwY1HZC5KdVl3McAYen8xtGiMZhGCrWkLeIxfzdvE1ffFk1S3JHYHYI2E7XEgKiP/cYCY
LdfD3T89jY31PrbY3REJpaPg88H5kqbB5uvQpOT6V8rKVvnT/q42bODEPf7IVx9hh2gcYi7DiY26
dsl+a0pHRSHwZOqUl+xKWmG/9Z3CFVeYR0Upgo9joQNCT2BR1y80PaIGAsPEXkS40gzLh8BbW7ih
6UgGse6h4Nds1nxkq/TkPS2Mk4AoDnLeICdmdjc/pzn1lvKXxARSr2lqp4l9/wMprm6k3w94acUl
Dh+39W/nQFdUs9pJAsRs8giLC9JfC87i07Jhh6Wpsq9bkRa8wtwCepjM3+NaI5OicU9MLuVsmqqB
Ok5cvQGRgBYi07bTpL7t8Y8AoBCoGTgkG3pRYHvVgE2IJobXYtvW/eaEgD7NFK5gerAr2RmXB2G1
4jJOWmFSMrwo91tM2wyIR5ldnD/leRP1N/zh/zmJy2bE1ViRP5/71m3h8o3FSJBQmX/uUWD2UTK0
ccTD5yBFZJb4ZVrkV34Ectcy73lseYICEX15ylq6JJ0f+7ZIAfKpT81unwHMsSBoMPNhhkuK2+Te
oTHmCZohr51CiSwDLFsVuKAeuU9Nvlvw6L0KgTowPULrCSPDWlGT/pvnlRwi0xMibaypCsjNzXq8
154lqSThmaRzEmBhg5wcSiqc/6CUuIoXQ2tVcJM2cPuiExthLQKBxTUvYwsIVgVhIeHwz7SQcvXK
yIX7DfRTNMW6xvQ4Mvk26sX4G7eggBVTt6fIYURqE9cuqTshnzw4qJtEeZNH+dNSS8ajp3M9s+UU
CqiNSopNqjI8wg6f8grNoM9hjH03zdczk+T2mFy0vUrutAbRK82+r/0kxBdUxOcOiT+BRUaWX6a9
mcluxgIE0jXRBoQ8pU5kmGCxgWQeBsiSSP3jHOHOgig+nQDokrmkTlI2peTCecDZCZN0aXr/f7nI
xQFpeOjmCLQMlp0HSwNJXBlLNp4W/bs857tZU80x712qvctUU/2TAgnaeCGYMGcw0RweHUf8VBxE
zLDe33IWaPanFaGXfE4IEpBpIsi96LooTNiLui0E9sd4ZCdpvodqrmQEq/XiksEw/Nad0ZNUkfuH
KDLir9vFHKx280q9JCyqzxF+7fxgaBtFTEYJEQolHDtChEFF8vjPbomp4MBmpm/cBMXH13FNQ1jV
pOzTeu18uuJNHcSQCx+9pKGPDVKWY0YlTs1abqaKDOjTgkwHkyIhqNPwZb3ahdio/ogy2fzIEklP
ZXFtb0lxFGtO/Q2n/OR+Ub/hOLJd0Vg+tr1JezaEUwm27j0uK6NKXI75SSl7d4dNEsR6aRjxVZOG
kaHDZd5OxatFp/R5e/Bpjf0d8P/1Sbome5DCR9yYdR97mVFDK/3sWzc70CPN11PE7FkmZjrFwU7x
QP16Bb/1Vjk417IbLagWNYI/uZYaMqFQBLqKAtsR2SCPGu2+HdlNetkPSGCOaWe4M0u2KBMVxLZ1
I+e+hhW2NLx28DZknzL+QBoRMSmMVJVtbIQERY2s8W1KTZ4jxMsQS/WDSR3PHDry8tRGhaaBX160
pfEYVB6NRsOwXh1HRu6dJYHVfnBlqq4kYvs0QuArRAdX3S7f4b9zLWpnciswPDZ/GZzyxyWG3AM2
SUjA+6RrI+srrO89fycEzPLeLiOuwwsKfRJZAJsH6kumexrZw9Ue8CMSM/GO4KQlbiIuaDLjuAIf
9Sw24iy1FBW8RLRPlcDuI/v5aDaWHslLUQitv+dsyDVPFRzWVtfHz9y/OFsjNazqj7gZuKVSGbfR
fqVJ0fKV0Ep5a6fd+sqqW1uV9yRiGjoP6cK/m38GVPgLKQKDHoD8moA9TAzZetcT+4RQHpCfQlap
UsZa62u4J+xJE2MoyyMOrgaMZ3ftRkdKxN+aR9nMXKO5y9vVLrCzlpMHO+E//HMEuaxEfbRRHDy3
Lh0YBFsIvT9K2dsOcrqSRebKwBABW6Jj6cyWA6rSgmWW8fpbjw0RzrNCCmgEU55WnOS7/rh2y8sa
TZ/5WugH2/HyZAewWwgQUy5hOQLpRYI2VgOpytmJMES3UKKGU3Sb9Xl+++F0sOdMxe/s/Cv+REZj
C67fXJYnfrvh2Vls88qAVj5PklumejLuMzK5Z4fcCvOlcaCeoX9sd94LQqV1OAxgV5EvmSkEom7v
novcjMGlqvhdgy6u9nHa1ZUWOPUDQ1U536l2KTPAK0MYy2cvlnhWTI4+I1+6knPS8seT3R0LugMR
cpDqNEz1ETjfwHL1sno7X99HqY4bfp9xr3vWFcG4k6mmNLYIZlixZOEu33Z8TL8AUcj+NyC7vIHY
T+IxN0TMd82oOyCIS4lOzvhKyi3rYJ+z9xtHyzGGrf0GPmlDBpuceoRW7w18EQIU0i5Hhu4FLwW+
TnomJmsu9f6opva34AwqjkbfW1dyXe1FY0jX90HpKmFFZpg3dlQTy1HesQYJfiXZtEbLk5V+fzvS
XGxHKeqh7ao/hfo9baUYQ4pPOskSkUrcNmckGTau2wbKTw6MReyFs86ymoExbTVtxq6y947++/0T
0jXDv2fP0srE1GX7+coyYcJKnQLcPyqzAb/ic+4tNLXUppiXi/KVTkJzXtZYJwXLHCy2mCdzyH82
Jv7O7TORiMwcaye0oiUpAvRrG3uB+XJiLDdmbyQFzHH7dcPO4KxoRG/9EvChAcTjhtnj/8ecpXCL
mbuBEMNOlGPpKDuMst9Q8TgejXLHM7ftFmYeNWyS58WDMvtKgctgjmunn0bd20W1zWDGkrbO7Oew
vUKseW3Olt0eoSxYJP6BUrOSU9IgzPDYylyYtJwiYK3OP+ZnVa+sgaNWuZwpm4eSItDxsAdW+g4Z
lcGB/1FZgbGa5O8kNprtuP1cn40UE096/E27w+V2zbr79XSI6d2US2Xkpj1eMGw+FiBGPjxTRwZz
E+Amn+a3foQqNjwa377tNORqRZWLFjQ5dLGzrNZNrjmFwnhBJQikFDSq5pnAm3ga6z69wnDh4T++
cvAuHE8BGngSnV98mkZkDsVCO0J5QyyiT+/KBvUMt9Gnax1fBRnlshdpBu4wECT8nQrcsYDCOIh6
el0uaTOo8yv643fBDx36MpfYfJI3YKccp47EjRiYOdlYhcwBqfWw00rFhlEt1kfEtaezxPFC91qG
6yySRS45SKqagd7UJWeFiuj9XKv1QrJEavUYiD/ee7NgLcL9d2rbG64GalkPZ3DJEKvC1fN1dSqj
pc6rNmTj9j6sD1n03flsZ0/7ds5R9ibDhb0AtPszxPUv0k3NyUa9G6bm1qTk9jx/nAeGOL3FQAej
KlrlQRcIlG71ZfpmXx5qCo3KN2IDVd8uJeAHJs1NSDuZvXvwUiP1AvdNP0nVnMioEgswNnyllAZE
/6HlVGizFseUfsy+FmQw0PUpxVAvtY7DuYFlCAd6wBGXK8JHjDodsUMH4xMHhe206JpAkqFRilP4
aOENj9RtWG/BBR5Y81ZOy6yz1A91hYwAAMynunPn1OvasqxZuwuwqXDNB56T4yoTv4YZgqliK341
g0IGSv3lQl3BmuQASty0MMg1rayZVmwsC2Qo6J14YpDMRTsOfDCmrLzqcy//EDnFNwPR9i7TYakA
tDQrNxaVkzqTs4uw797IhIk9User5F5pWApKhXUa1jCrLQUrKJjmVfyW9nKj0QJchY9u8bD4cbQw
ftAN8XY1mOAqB6pMNkiCigQ0ieEQGQS+yRv/FHaA2Ajkc6h7fRjmH72J2lh2hmlNaFNYB2ZeMSnS
lRpiEkKvDm8ayN5EkFUzzPvVlbjDy4fMg8QZJo8HWNF39YtgUFQNwTXEFKrxrmxnkBHHyTGzpAh+
QuWLYICS3HvSq8575zvoeQEKX/Nr+Ukr9rbrCEZ89ZZokdZ4y7cfl3MTxwkfY0SIogvo+AJZ93hO
YFQQhEP/Rf08IBu7VJCqEdalplumiimH9m3TzzzLTaNBzo7gLrs/QpuNOhJ+kuKu4nJMMEQ6hyr7
8Ohztm2k0Ezie9OglWe3G/tLp8WCk/50CeCnM2c05v/HxCO8AM3wUK+DRylV+zJe/O67Z4P9bmxz
C9wudZHSSlvA3S1CVVwt++/fNvjNd9rdHMi/AfgIJdAtAregqnC9XvICBUXPOJRO9Yd5LFEQiTle
QSi8FTsHanXBoKWsvLqibwt0qd3hvhkoNZYQGLHVQxpen6KqJLgph54l3q5u5cagEdguUjDwrI2C
RvSWGFN2DlM+u/TjxIV9q+o1T3CIkevGo34aexPo+SDuCH82GrBqSuWxBb3QB0AeraRYUWqqMiUh
dNbotEz/Hd4WP7D3o29hVxUmZTRFR9d2WrPwXPIZ5lTBNahmNwW8oaNaCgSRq4Wr3RhsDj98CUO4
G0fQp5qiKxQHvEG2i9Ls/DN2BW0VjM058DAqLExQDaFRPw5DdSsInnUTcxp13Lu6VEXoHgRIcryA
3OvwFI6bFI22zaVQQxV1nNyclAT0iuSH7MN/7p+LTZ0n79sYWmJGJT4wmw/9BurO5byOO047QsIE
z2msBKoeGEZHOPdIEQ8iiFfTjlE1zpd+NtEiWE4dQGZ43L8ce4EB7/HticCTPf61cp3rWOvCm8RP
BftZADFjK213DiFyVD7qTSRdJFBzUZ8832h8jjPhv29li/F/Ed11fy8CtaMwSRpCxTrGzG+TmxHH
AZaGZ8TgiRBFFchIhE5ZJREGmz63E4x0x0Ccq9NW41ojYJhzvScLkVs+5mI1GAAIMUkUJLTD8CIW
phtsTnCOra8GSMS3iYAUCagzaS5wG0GAEaIgxbtrDgXsKKQaqkUW8VPwDky24266NmkQfhlyDvF3
MR09agDIWNK6jaDDi/wqlKoEZDDBvTLekwugazSwD215ScQoqBEw2FKc9cp4KZwLeiHmVCNUy0RW
e8jx1ivTaJdcPDz9EYswjG0hinZyxnjeRrdnynpgDePoaT/wMp7TnpWJa7awirK0mKZ20pi6tl9j
6sOr2VH40mzXbocJ+k66IvU01pABpSPYgkt2dwl1XWT1cVqdiMeSWK85ou43mtHtvU1S8wIuMh/f
4H/mlvFH+iCJM21pM1xcrshqEK/lFZDTolS+Ix98KX+cktatLM8ml7shc8HHiMIgqA72decOKnis
C2SDir69UnV5ujsoZNFiK1fUecGPxaEZdjDA/ubm910rUOVGr1f5mG4QBWEp2x88n6JGx1QhZF/d
MOTK2I0PJJymjmpU67kgGapq4wyX07c43AR/74V6cFeRcBIKQgXg4n8Pahg830npplOSfOTAgKN9
OwiHyiwXuzXEWAXg78I4Q9JUl22tUs9CIyiBTA6viMc5mReqi2NCk1oavDuh9rLCmlhcTNGQT8wU
kXaKIJzX+Oki52VFmxAWXUKQidQ9uQLi3KPpxdyWa85CPrFCToofkyxSdVdFK4CEc8CoJKlG9A7y
qFLceb0soB0a9YpWGg51PeWPSa7jV/An5/F7gXneJH115Vqpl5fJJDIuggd3/3aqdBUZwq1+fSmq
ojxhYukcxFX1VGZ69HTUZsGt/Zppea+UF8kw5Jn1j7aOS/K8zhu/VdPWuzXOcWdxI5TqkEzim/ph
/Pg9N9ZjjCkla/6HTVv2quJlTewEJeeAa5KyUyPK96whM8wpPHRWWQcjOd65RZJc1ifoEiiNmL41
7YVvVqOC8iJvhXbvhqjsyzb8ByX44DKZScPMI7LEb4n5U9AOjrrFutV7oOB45uw25qdRgxT6IVsB
/jbqoNNc+He2WDBCiVfTThNCp4e3oW0YlyNMn4WZGrdyVtCq+piz/r1Hf3vmex9THZ8OZqF2ojTV
3IfdUDmsUZ++4+WMjGaJhtyArNR84B5Sk8EhH8H/wSzlzeOcQuGKYc7C+ZfBNPBQP06EjX0Q6/pU
OmLf8oc6OUoTCvY8c630QeYEeQwueEJLn0GJzaGQEhSnb/qS/Un2of1D3sUsnBsL4aNGyNgeN8vW
1nxljwsaLJOWTZaK4ZrabbplBOj8RmSJ2mIFX/4Zte8w85P8St8U+ooLYVpAzn6K1pXD3XyN9irj
AiIWDt+p3ZVGrxZwnjjCwnJ55nB0BhN58TB5OlTA4AJuC4PvMlKQaVt5aq7lgolkdXHMt0jAVil+
/1kUDTUuTxVJa1QvH7ZO+g/R20em/QCYKEKFVghyvI/+MZGh42B7ueWeAHd/PiAboawmpUDZXtgQ
8Inxxmv4QvOnNpdSIQuHEUJPIcgR3g2wZvLpEOZekfZW/6ogVD1ud9/1BYVtG/fnka13TgV2lu0f
459pNy5jH463VTA+duMSBeWk5YF8HnpR/sLbMmu4jIojjSXZU5gjnid6cHWAMvx5G5fNM/xZ7z/j
d+vB1xqP8rKUApastZFmUqfGva3SUy8zByQn3mT1ZU+x6IwHPp/u4GKxsQHYIGKczlxtxiP/pPq/
q6m/M8ymrI5ISdi59MGyj2hsRxGEgMrvXT+UNbSyaNmmZxOBul2lL5t89DzueiUflj/ILMMtkqEQ
m2Lc9axeDQnWzwAuPh7PV4rHvEddual4Ymtlp39ayFKxMEg1Jrld+pk8ActnukJSEBJNtIbCteDs
MjlJ5KXJdOou63ZizfZZH2n8wW1xJ//Ji3Y2PZYcklyGsKGlWLoUawHgctEQjWDXLYDmeZiV7Trg
WO84VVExpr9ey/pyKcvo/rAjMvgOo7aV5EYRfOPPVCiR+zJuno+UJnRF3KGy5giXnnLvo2ODIxKP
1wFLfInS9zPEWt83tcffrB1G5fZM8t5tUSGRB9P0jVtQoAFQtqAvHPm5Huf/FJkxEnWnIUsJfO+L
XqGJ+ldzMQ5yKS9/LM+4D0C150Y5NassY2pP3Hc2Haxydf7LdclbrnsGoULbrq2Plpc6dcJ1eOTr
kCgMZgS1HCBZEV2Ws4/s2UpKlPyYZPgiygn1oh1J5TADB8y8XVmQHgR0w2zG4M+uFJkvom5qrhCC
MGGTJIuWx8BZaaMMCk2BC2KxLqrkwGe3jYkG0XIh3bl0rLb3Q+pvZXWhXJFI/LaaEOvSLCMahAmv
O9IZBZWWM63hQx2Zmmr6C0zd1Rq4riUN6r5sYGjiScnshDo8EbFnEo1YmGXH3hg5WUQRSxDSu0ti
V259EH54qfrgsljiLfu9VjvjjX9of+iXqYATBqeMQfLG+w5u8yLKOSgeRBrbond1q28du54mygV4
nrRomI/hJpwJs9woxSbWkGHR6i7cUXwD8Z71LKz8FNykIuyo3HY0I8/4u3yOgdCLn5c+Og9Xl1KC
rT62c+xD6wCsZt3GJtl/HMYHuwVQWHV46w2Qbom5X7v1V5s4/TPf30r7aKUQSN56vg/XyxA2IZoC
uRtp7mzoIc1ieTgN8TpcbuPj5Ifis0fX+wq8FgA44L0Rgg9hbLFvLTm0T+uv9EBjKagElD+/0jaI
xM6BVtodQtXKm/en61+aUjg1kZ0SNZlBrQp0+gQxfT+JE3Boyg9Oz6ONOYl8ugDBjzxObv1UypOl
mzFj3tZgjCxb5mbEI6k2ZoJHuJy4Qd8kKnvyI5DRCl0mHqocqIdP6B+3pdNtbQeL1rpJPWUDJibb
wt7p6S0AmJ7n6tujw9rLHUGbR2qRljiyXP/9YY11DOZrw6ReHEyVaj2lskU/r6j0EVRK1ypM+Wvs
n3MneLW8kwJd0zl7mmqEmegfusAdNEmZdMDtNJVK78H/TU1v+WhcdPmhcl1E3+frKkYdYy/fh9F/
cvi7mW5UyPTftQGHtzbTNrPUKXMDESCphHVHOxOpIKnNsBO8nPxMSwWFIA+9ExjqfYm9Lw3rCWXs
txrBUBh/dpXXHVAG0DYv7AR3XC2AAg3alkdDAeIl1OFaYcwiRi75q/Vry0jqT93+2ELa93liHMjm
FSo7DNT5yU7bebg57MPQ1aBY4lvn3v5WPAPqGNRCt1rc9RGr41WeXxpsemVz9iOmJJvwCRqjxBdd
kXe63Uczy/81BeeiOLclvzMG5tUwvULlD2BvGKoUiMgBepQwRmwpD2PMz43raFGoHsl6M2UoatTf
sWbYlTIRSh4tQ8dRp9ZNhD/93yuih2uHJsaF0NLc7uLa2rJMQPIe7wo0nMRqdqdm3+kHI5pEilIX
cQuId4vGYoxfhqfW/fXHhkwepK4VUXyP5UOkFbRkD5vMHZMlYHLrndfaLkjgF62wUtmFHvxIMufb
ltD62cJulboWREilscrCpRnDa5vUKr6Chk1aP6tFd58JL3FF4m07LtIxHkcJOcrev5mcsdlzPBmj
R1PDGMu0mYpyf4dLsFpKz1hYVSmNvtk1Ahawj3yCUa6xU+nyocxZLVaBH3H5qPEn9J1xL2rfGmsz
XlW1SponhVnNS5jGNogSRbP48H+cIkEhtZ6d9dKXJ763VF7C9VlLqSlpRxyOgFk51rqWwEEvsiPX
Gt+s3IMAwn1j7MBKf7vBDCjWVG4ETcFysyWkmEcJbrQ2neV2vyEcbE9fF3BW66QJOoWtXs70oJKB
qOHokYACPe82y578YTWz+RlT95qZQTgYSUNacsv423+1Gf75EPvk1owQLlwiGexYE1T8MfumezUC
nCUKybsaXThdQmB5bjNtb+0QrbkY53D3GuMdjtXJpCyyPT5IidcQmS1SzzYFCsus9HAEPFiVcja8
qkdszeQOXvZ736F7vNnF37lEZQgX6+1YD6/MVItOdy5mFPhURlljyH2V/RQ8CD/ZEg6t7a/XLOvS
wa9DrZ39+1w3ugknMeS3TawYBDABPrwnFrIsL15cdGTcfPp5JgL/D4YGuU03J9Bvx3L+52mtnZHF
FfmSIr2b5pN6OgSGB0iuCKU+ce6Dxktw79ZboWDcOPI8E8go9nTzgRYytCyRMD5nFkS4PA3e26jL
e/SxJXsQvRiSYIIfRuP+3JSKis9FnExjfX7XAD8s0Z52ZEiLTPFr++u7eZP4w4fBxFgW8ESx3CMz
U5KdPM6Yl62toa5xoLaqw2sscGerD6NK6BFGVMoLUnefBUdAYpfw9zVY+9IGXMUTqbMSAY9DodQE
7NJddXkzB++j9gsfx1c5GqpXTCAYr5LenRRvoiQlVQaO16Z0DQlDY30+kA51J33l4OJhfDmCEfLF
YzDU0bXHRBJtvBJ4nq3w0LPBfk3Q3KgVJLMt1wSoeUqEcode8Ozq/mhYXL8SYgjS/Y67AJ2MJDYw
LLxilZMcpdoAYKxO0GOA03/tReicshHOMiqBg5sHMShkce6Og/kNdGL+s/WGmN/UXkg3G6AQTJuo
/+EfCTP17BzSgloM4wh0ZuRs6FtgtW3IcZKSg4NEASuESNi2XtHuU71GXUUY/80nW+cHOhyJxSEZ
cCJPCehXHswRBFOWum5QP0t5XoZXHZNoYZPi4IuyTEcAHtM4YZD9kwrzzDFH7N3Ij1guP5Zz224+
KPHhMPvNzcnTSBP/JZJZ+/D07dZEGcWZFaXqyAenAcdM5D9s4AFgbJFfoK+z314ECl6+WWpiOCfr
HrqsBKoqZ7grjxISRxeFsh9UprGMh9/fwIWMDWxVQJVDvK2nZFi52jlZAVbPKxAlckAIS4ur4vxo
zgTzrHs9GB10c9V/8nlimofPnq1gP6abJzmyAL8aQcCOSn1aPELExqIIUfYQF9jmdJ4iKXhWwolG
1hhrn/0hp4YnslHCnC7KXnUN/Ha89Bgn93to5a9a1MfA2L4g668n/8aEk8RYlResJa22jaXFzP9Q
5rh0uX2RSg/xhLepl4zxir3+gdYEsQ+FzULzbap9aIWTmTH3QJ3naJ9DmeIxJ8Bf2SjShCROa1w7
IC4H6fqBCNnBGQ3YpRgrWvAEvIXOCNZGT9/+aN9dsjI78bhBOUCnNdYzz3IZqF/PmpVuPrE9yi/B
z0DD7zOl4+Bkn1twPs0D9Pf4Q6HX/UH5MkUqwTkweDOVGvtgSxn6I4j4krCz6Kye1mwH5keDswrc
E527fOaYHyX5BbVBvtyGK01jzhVsCp6bF6Z51TNdwTHhUi/TQgjcasuUljorn/xveWOOseyZqoUq
8BT+205yWCzWH+IghUVEuiJGn2cNLLecLXi6mv23Ravfaxy/96YogYoEe3060ucR79pQrIPdqtQM
chRr611ZkN8+r00aT0wEPMjHSG2P3nBy+4lvB6Ceny7SPPg0dzhhMaqV2Wbbt59sopBYv+j2ZiD/
noBgqWrGfaFvnxaQj6jK6x2mMH/noWAD9jPISxjKcXPpbiFfhqohMGCQsTj5B5MSAW6cVkHyiGPU
ULR1uBTZG9Lp5eSWolT6a8aQINBiVrg54EgSC1Vhp+L3BZeWWoSmbAoJJ7gy3eLRzIeWBIVrdhGI
APZiUO2KC1Tu4H6z2qnNHamfCNsRvzW0CoxDpf4ExIo1dmeGnoXmE9yk1kng2P8HU/J2JqpHabtk
Jrcmv4wAmEui/B/WlI6ELJAEUPCR+u33U/MlTGCF0uZqVmfXsqjOf5SXOyYWDmJlJIQizdzzIDs1
LESUqeyEKk18hdTcYRB9bRUgaRkU5mphwJkorxWJjh6jUUDnn1M/z1ReS4BhPaJSfoVb5oQjkZG1
ZCgEAH2ZTTPH8h6fzmOfvf5ODv5x+CONIGnsUrfeG+XBNFT5YXI3E2i/6tEx3qIg+ymubuSYWTJf
3gtFm0ZKo7OigxNeXJ9qhwqBFTnTl/hjN5xNZ9pgJoBgCkLzZsikNYn4sm6pqKQSM3+9mG8llmA6
xJUNRi9r9q3W/SnSzcnfFSzs6rMZOQx+lR5hNKaBz3KqxNUtF6yo+UNw/lZKdoi/+Upxfcf8xhE+
gtZBKk/EWwp6xNBnxM+v+vCCMuTE7/m46b5SWY97z+aOC/n5neug4QJriMkrsEMtCfEjeA/4Unju
CmxlU5z/i2BrCUNkot0IRICbUCkm2hbDlSP0m6g40sjZ3MCAla9COGF7pQCM9rpa3CgPJQIkw7Ca
qrre70rG26YBV71tXQAVFcpxftLNcLZ9nHCckA3Ly6I8fnCWgOL5Npnv6JPqTtKETb/Rw0QaQvv4
wmWKhEXR2ILR4L1C+Aub5K5ocdblW2no5h7wc3VWVMs5k/Y5rciBy3iN780CaJkbtqpW1MFkO0AY
uCgezORFV+sXiUDlRPVHrC0pANI8njk9MM2QIf3j1VumnGi6zohySB+a5tbW/OvMsKorz5OWKxCH
B0Gh5xx3RmdTPtetSoYZ8/plZ1eOMhR0wN8Sew1xFXAHo03jfyM8cNEMmn695QLAId7uQioIg3h8
LszjfEK3IscjLBdwm6LtNZai/z+HfvBj0uB44xlnxEehIyER8ZSlMl+LtPKFaENkfpMuWFnd0Kt1
s4rRVr0ZZY2yre0TjuISbuy6b8T3tDd5y1GilA5yxhtu4qkqJ/g+1ex18H915LIsGKm8Oqgxs/0e
RYQGuxcw8BwZHHl9EGIiMu1b3zuKrrZqKpQL5Gzymb9G9AUuRh49J0GhmvZiKpmr138aT78EO4aX
cdxbIHWWgm0idohSYZ1j0KOPX90J5AFNvuwdKvJsgXpnhfDIWlXAb0J5ukLx6Lo137UICW1PExZC
QpfUfV3T0NGtDk5EKnQd0kRmOAjW0Q2ilNZnzz9i4a3f7Q5k+bsfdt14otaliOZ3+4Krq3Oq47bB
8QXCzRwatrIDqXRqSBC0/oyExBFgdWK7PVGNrk2/IUnAZvFzCXUuo5KRdgS5Ue5+XGkkaHm2Cbt2
9x9sAH+hq2w02D9+edPjYfPJobHR/7SQJ8Xt/MFz9T6yVZG0RMypfbExTBuroG4RIedweV+wgdPd
gKCLeODgbmZPsK0lCEniSUeRjGenkxb3sOKGGT1T/3Z6njm+Pe1Emr02fzPcMmYM3gSLxd3Wvbo2
haOYbWJvGJD4BOo23ZdwHmnRPBFWwj6G4JRSNLYMkxsOXlA+GV6/s4a8UkUas2+etQGCbeSDxjSk
dLpzLSr5Wr9xmHw72wUmUpqIzk4RTUdgPioOSbocUDJPyeuXtmds24r44ppBmkUK9e9ADt6j1yKi
1+RyngkdFVbUHbRcDwu8vbZdtdl7V/Ra/a4R6iShElLtp749ToCjEqKbboaiQdWYDEuF5M8lsLgB
mjgS/xdUC6zF+3IIScsww3WIOedac+XedSMpY8dPIPLHFZ53trqk05jXx3RO4ykuFXTfj3S3EIWB
kp6lWop6swyNlM82tc4euKXgYCAsfoxRURLyrM5aQoM3MyXL4Nvv9O/aIZFGlTbuS4Zy+mBJpfLK
wj3LDD+AWkolvNhgmjxMLPGKKw9S0xC6SN+HGY4/+oOyKDQqZ62dMzssq6+nPN7D8C3gAE9e9Kxv
jDOFwxfIwQ2c1VXTIYiTIdbloZJWDItkCQvF7yOZy54UF7Dh+oIm7GIIylt3VN1fENJEg71vT3pZ
nxe256h5aG37YO/pTP2kYKlwyG25rBug87HKPN4UdqiKWVwbGNRWeXfXBFeuwnmQV2OJ5oczcuYW
q0jNrtrpLgz2H5pfojnGM8glYkZjxatxg71TO78vUNdwHWaYHODqr0SNsf5zBROrE1iUzbwtW6uL
3eqhuQT2tWOtq/DsSufSdGVNP6/FjIZF3vi+yHaVrs0ZESCL51kaOgShmRSAJLQT7OR3OZC9P+RN
70P/HfOe+QQTVRjMZID92NdaaFIyTfiJivKlLDorj8FomNh2SR5+BZ5MVQhcWSoxaPugafHbSxAK
QK2rdNmOQvrj/8VNBaP1ycnyhAHOiaksnNMOblG0BQU72HOIdsFwuMKuxgIDxKgWGo1EPrweYUDm
1cmien3ofGlNv8mhShg/PDth6p+rf66mMDvD8jJw4MxNO4noWR/M5Odls0GuV7PgJs1jDlWUasNx
7BqNs0kyB6LyjJf3lkHn9lymWQmGRGXlmmm4wpIIHMeLYUIRu8C5Yg6EpUb1Bbd3uJDEcK00dZnx
r7M5prWFittw2AzkDPzbHELnnZxWIcSYr0TuPtSNWREBL03bfnPdi8NLGRVnTxARO6bSWaTqZ04X
+eRl2ncJdSEmjfp2rkgv29dGjbWhoNgDbzQzGD0pWvHLukZZRTIJMtLKPwEeYUdVNHqTO7AsszfR
ZxCxqdbQAYsr4Nnn6mBKD2OB7S2eov3o9fjOTD6csg380ssZYCHqww+8zoTef14eQQ640fzqwQPl
vYEYcHhDxscfJIcZsj5FK0Ik3IRmW190A6Stj6OLwo2mIQEH+PI4JuOwaNzshwdGFEzk6gc8CECP
8NThHhAtZ9pas5u3l5iOxrNEbYF3uzfyRsPq7yjuh8FqmpZIQ9qxvn5bno3B5e1B4hFREjdDy13p
6CwFoD3+shVR4POm3wbG2mvvkLNNYJMtY5znOqqw0K8EnNrtqx0JB21hVHp+2x0OLPYOeWw+6NQD
HTnGB7L6NJsDcYK9+GXvCYfn61lsq4Pa3z473iZnayQEvsDGdUM5M/qiCKV9sVJCF6yJq4xDw1RE
4kSuwEULzcjMPthAvKqOX+a9ZcMXypgKAYygQCyJtpdc65LXR1PUZoLjPIE8BkGXqxxozKBAO7e5
6vmdIAbGrK4ktmyhaIbuP4uslxTanHXDejc39y9i+qSk0o3sbuvqyosQkXnHNMOArP5g7NBCe4nU
Ejm3XgKxk1Vi8YnwcTnOumh2hiwX3s24ER5qlDgQtPLDGaTeLbn2g1tjw/POzPII/pqal9HkQeMh
L53vclE/HAp1Q1zFV6wMExC9wia4sBeeX+hH6UOg38jsL/5GwWuEgxGxiUEIaI8jZ6/c+QvM63BK
lEgzf86jl3nNUd7qC7qqmfvZPw8qA/l2kjJagIZzYAgO+7zRl51vn36Jq8BkmQomxHlCeeXcBrGZ
UAR4nBUL2U+6GRWaBI+SWSYk5sLaqpv1ydaWtmbOy9ZnwguIq8E5hHPRnOodJ7/kdpPSlM9Mkycl
lpRUBg8+Sg+DPH7OZfH4kD0q1OV6ErxJJ9EI7nzAJ42shxXZy40QnIEid9RYshrX+tXRfMo0Htxa
KsVt6CeOQdn6bgwp/ijco61N7qWKT/glq19MwKbZA8LBGNE5sxoLNEusgHqGhy6AxrqpKtH/Dtbl
dk6hakJzPE5rho5nObbm1zqxwDpiqISZ97vTpnI3su4uqXOdIBqAfPJ0GhcvJGskMmVT+uhHYu+6
2Dy9bE1CLa6ufF7t2qtJo/8W4YKnd36O7RXu+cvUHgCa5fDrozGYE6KF7gX6djX5lyZDlO+6oIjV
HXd56IHwNLGWXYjpDUhBnAiN8lUGlcJ9tMjm72tc9vdvsnKxOvnM6cbaE91VLHybtGxcK6EOgVfR
faOAnsfVQy6KyPyFhDRhhz3FshGk5wikze7o5XYtQbUNKLbTMca6aV1ilIKt0jPVdWFOeHpVmB8B
KCKPs+Cv3u4MnWBuBin/5OJ4r2d7Cv+dpPlcCxnRzaVyi7+ehuulUjOXTTRCAHWZq/4jWnsh3wA7
P7g5mUMolWnzmbzloa6kLlnEvj8yBb86YNs6aOj/cZGwDR5GJTL/sVg9iw9qDnEBSCc1gpZ6HyTb
lbxbH9eyPSD1XEMOagLKp3cmZmusyJeZA5PAY3ceODKS2q3rruarHBryv275CQqBLZjbwY4w/m4v
hxiYTOMBwv4WOPl7kkBihHrlO1coYQh03DZnsGjwYleDH8vGo69QvwRbPXxbv6ZLNHNo0P9t7TdU
VszfglR+ZFRwcp/D7Q+gwPaIX6LXHtixqNVznyr0weGyEqq2WdjJlp3nRzKMe4U6bPNr9GWad6Gy
p9PwA1WDLVdB/N0X8pNjd17W8C9VGY/aNXyyNDWlDwdn93q1JBHcrvs7lMxv4oRDELUTKszlVAua
AV9vJm41tUp9t9pq8XmKlJK9Pl0cByrjE9e9/GmpLwcSHP1n0MJTkI9yF2O6eEXQapi461rZkNLw
34WegHB42KbODDDR8tE5RT+Ue+DCfZDEpdNoBWtVDnknNd3Fx6rG5IcOox61iy/91i3T4se3gS+A
73pVwQEpK5eQaOgTSj8f+JKB2by9q6atAdJxBME9JQw7Pkj6rGAMZ0tw0FXZ+J+548Y3bYHCKm+W
aJXWfbBHuyPx+TJbal9ZLKJDFCceKtFt8yymH4X7LtpFYF9mLjSj8ytJMZpFf025DNttL6pGmzJv
U0fs5uSTIMD6OVYVPhM6I4IeXu8cUIldt74qbwtQ4tGo7Wjw01K7xZEN2+mAaAPWca1pKPfm++uG
UBHiDwkewjzmW7f8MIgyWHcX3M51IlDfd+2IjOnkH9yR0gTPzjMbofpLuQhvavg4abG+GDMDO0f4
wsItLMl1pZ8rNX24qgSkm+E/F2gnMnsaNl8ZIlDlxZxO8jfZMsCxrkWImakJ+YDZWhXYjuvuvOte
DRPnbi3Nhsse9Aff8hxj2HtRQ9NynNmfO1UesD/SxX72+As5L4ouWcU9p/7mDWh8OrfkvR/6iKza
KOpTG5yUshnDq8O6Q+kA5TLsf4xxOV6ht8CHG+yqBt3BGXqog8UX0SNEZTGxMju6XlEVTuMXINjH
uowNl9wFAcFgQC59dQtfkuKR38JfW3XeRBUKULnBaZMOpue6MDLHHRn+faQvx4GDcjvIexm92jz9
OUEiL3ZIy8lq2pj+34mdA4cQvAcml+98cibkoVh1wbmNwNrfPwto2XzJphYL52IAYWhT8/yIWH/+
yegpcPIHQ9M5pMZe27zlQZGZHjRyAvvso5eoxacDY7gdLoJea/4Bmu1ScpSgSP1HQQFi+qSztQ2s
fVAUmcCL9kaM/T3Masmqg66lmhCTiBK7pnNuG09C/mQyBXmat09NfdyrfQZqAEZZI7hH0XDhxiq5
sQtieFWNAxQe8ULtCbIFjCM671NyLvMChYIMPiPgWLD6u91oC8+sI/AHo7VSLXz5o7BLvgP2nG9t
axquHO4frLipRKG48exhXFJ0fdXea3ADLoUWIAK0t38ZVdZws91dMth+frvjYn5XBtaWieLH4fpM
87krMbmRbkcYrWOB8MD4kz3iJEZZkmPr7FvtZ3nvrT4tXO4+9YTAwq5Po6JnWtBkgPKodrxTzgjK
OvfnCKyKKZ2tyni6jafgSlT7rKPSO0kaTCI4E9BWs1Utu8le8wbXrjDCUk9eGtPc/XSIRkPqlnoa
VTANUBXjXIMo0UcpYCTwMB+cypcSSceAeYKqIcxxW14r+FUUFpyidhpgx2vddxw2lxYb6ty8nZ1K
xB0PuYN8d7y3SVNMqqdioPJBFyPD8GlrPIUG781nmlOCXJynQPIzUJyBe6+e/+uPw0VaEYXEL5tM
tuWrVY6QxFW1zQ96ugpPZ/iRxzwINSkuE2DQE1Bp0bEAU2QX32f7h3GQUQVMOfTSXBWXSvdFDCRk
JRbKLUgjWJBVbS7Jfir8MOZ/Sv5w3YjMX5Ohm6P3Ch2ZRdnscEBvJ986HA7sIel6sOy1dxZpdS41
jkMQ4THJ92LxLqke14Sbe/6wstH4K+jB8ULn6Jukm42oMo+Dexu6DmqOn24JyjJR7qzVWmiVe6Wl
UYCw1ZzFALFVQndPNihUFkiHVN+fYMIBd3Kc04TPVTxwuu84d8dWrM1LCQD9B2qghKE3JRFcilcB
kxpuDcIGKzqfKQNKCtpWFynosiVJHaZJAhnGN1P2ONt3YBFuQgvQIIpTZFz0X/eMfRIKWwpUtRzC
QV2uJBjn1mbkujVX5HiK22+F409PsENf88H9CmZEPr7eA31mWfzVmYXji9VY+XS4yvvN1MZPx+pH
MpHX5qHySuzZTBqAElt0v+y6v9uKc3yv3pGUxEiAlUufwJ3NWJmbuoRKijy5LXSmJyJz5GaDZfy3
uji1LwUrHfQDwnbOqisVoywVTBE698VcO9MP+RT8xUl5pzmzZ18eedOP37o3FUUOf4gWoxH9qqcj
PzWx+tuBql48Tym6UdQfhVsUzEFuHU75WTG2CxvluW0M2gEYaGDUUrr6Ff9171dl8+tnfkV/eaQh
5L5lVThKibL0MvHjvlxl6rhhUmUqo5tRXIYDpUG3n1YSQJd4cw62dDf+9X2eoami6yUdziUQoHPM
UkrRh1blc7Dnk+sBFCtoTCebeSIBrvk+MDiMNp2zmnFCiVXIoFKubt7Xroi63stJxdS3WH0GzC/j
OjwH0NB5uoeoL2wP6bHyWJwSF12jLPu4DhKQ0o08bixKl9Hc9khqhvUPr6Gy3lsUM7hgtIjcA/MJ
urE413DEoMSHvw6McyEPCK/hv80g1ivltKt50A3xM6AZ7LKmy9pvQCaySQ1Jw8Vt9NSBGYsNnKho
O4cMkW+nAYek6v7Bw7d30CjQXePrUjDjEwNMHZWCMIS/xEpVsekrw/cSjtzfT++jE22pJ141Y5iN
JvpI11O19yCssV5LXkFg3R9R4xuviR/MP0xOqr58mcVsEAWtSzoDSiXEZuojv+upsFUWNhBo81Bh
0h2X/E+590aJlp+2L4RvdCNBZLyCb8cK//YAWATvaubP9n2UOaEgau92+CZUwD/3bHqrmwwfxKtX
DTO9iYNIqxOQDNL4gUmZPBqrTL0pdola10dWPw9oFMs49AlUgzxCXFnWggzheZG0e1vadIpooz6K
/L4yJK1ScKZsShdeN5VlTNOhxhvhd2ePkb0UqzioCXnwVikMngSR0pA5rICRKkK1okXwSz8/Q0WP
ijD5ePNBPKrID1i4w4XodfaSMDoMzv+FQMYd31v4GA6gKFK0FRIdKEGkw5i4xeP2FhWZQ3EWXTYB
gbzPpDsppfc6/yLmXT/z/+CHqP1mzPJQl6MVEKkQ1/mJE+wBbg1eIOr/ejuZ9aS7JoyLQKHHrGEy
86Ca20FSfnILKhQo+v1xAdb1Z6gXNMsUi7HVi0T5oBSiG/jtyQlpVA56TkrGzWhqscxAIsZzlPnC
NMGX+TnqsFICAAQFQ5lqvPO5AYa9HyWzQvvszCl8E7wRGbyS866XYm865p6ZAwSR1ZzUj5GerrFQ
eo6Vobpa/hwYml8YqQYEnwFWGzE2elgnKt3bZaREcvXKEMemjN8iZZRbI4DvwsVNgCzyCRWjEXYA
ktnuzFlYgl+DxVoBzOUrwnKirUvgl4XHEszmUGflEYHuK5VEUF+OLOSZr8HxuckFiz0sHRQZwP0+
4sVHN/F9aXWEzHeiSPRo1aQuqrQGx6qTXhh7cG+emYudHuORFyM+vGv+boZ3jU2y+omdEXHJGg54
JweoKULvHFt1gabvnRwGuf/c8wMF4fouv6J3+z88dKF6eFhteFf1kUxmmrvL3Jz+CXXfqf6nGW13
PjchB26QV03Rq2WhOetVRY6YU/O/a5Ll8AnDV9q/eL1dhrv/DtFBKOeURdsToGv3vvDhUJvCl0Xf
bJ0GEhpQYon7yZCg/ofdAC523cvhx+mbTs4gtXSwnS6klTl+0LhOBHnY8HtEZq3maVkQF5xPQ7Cn
ZM5sTGGomlybnGTZpfFPuN1pI5xYX5Kk8rbbq2dVYLc0X5sv3dSua5upgly0hfErllk2aKqiU7DL
nUioIS+DqfEKAgpQTHtuKD/D206doGGq4+bGFPAW7eWkAklZ0rFyU3Z8HqiUhnOBp/8Ye6AUHi42
i2s5Zaliffkj/D8g9/kAcoHCf46OuPDqcYL9nrbJHGsVQUahrQ5o8Z+V3bT1v4NzPi4CZ/u79q3o
Axit94lk1rjHvIyDkK2cef/Grfu341wOdVN9LCdyxn2ZMpJBrAikVH4modCaOuInhmLq7gug6Agr
qkbyE0UMRBR6SrH64RUYur3wSqpdYyOR8YtDHbVi0iSDOxe51BTaPpoxvJUdEWaAPC3/loSd0vC+
2wqU81bROrW6Q0Seo6Jm/Fpv23iBnYp+jdN2as7eU8oHRkK43m8HgdQM8uZ9lOSmlwvDx+ks/qRK
POTwZ9ppjaFAHVygko2PtSqpRRYRM10EZ7CGUUq2dBB2I1R2DkoRoWEvH/ye7au2Gn624qh4hrxU
sMZe7l4pmlN/ta874aZ1bw20ymwSl0FQH6393CmCeY/xwcHPTdVWj+8lwTml98mfys0oAemPSuwu
IPSBj8lAK9vLNUZ0ddL5uEPjpg6pnvadu5vM0qqT7igcrnulfKVt+oz/uuz8YzFCSVkdeaQKD78u
MmDXlin9FlMROHLz7eH45UdcYqmZ/FpPIWNkENqFk/iEwezk9HqwkyHsal5ITjsB3M6nY8sLSUOM
1fFx2KtZ8PHE+j03qyuqkYlKq+aLX+8EuhckiJ5KFB4GbPmQJdP/NDwhAM6nX4kHuRocbN9Qq/j/
lLB9ZUMoHaSfs7ZrPIh169zDIrD8NT0/2+g4PvJUsWtI0mgv9YbkxL9Ozu8Jy7Va/n/5oj6n8HlO
e7zq99vkGtd5viSnvZ8tbo+siqpZAo3b9ak8qJerNzZgxtLfNMHbZBVOy2ckGJOhXC13pZ9gma2H
8WuYBsiZqeG/yrjkG93nyMPzGbfpKofeutvzBOksy1OhMNLROUSnIcHPtDR+BIjGJ3OmvaSh3TXH
abP+PJKsRMuxRYurpqOtXdk0krP+sS/9Hys3sWrfmSIxf6+quBb5qCPLSBoxWD9PZbIx78ZROpPg
tjUYhR0eG2Hp0o430hm1kp5DkAWR3f3mZTkw1z56imOVVFAFpzOLW+u9X+EfbXw2odzegAMxRq5L
R57WLKJ+Ct4MIlA1GB5T2wE15t4c5tffxb8bXWFqVm5UVhsLOkGAw0oQy4FtwJwXuC8RSnsA6OTF
DxOAIOxCkFs25LBR9S29ADWealMCgZrY4iobyUjt/ngagjHDnWQO+Nm/WrHexILguhubkeOkqH5E
TBzh1ROuV9dQe3k14r88fv11gBuFt88Sbs+70gHnZqQDx5Iqs7paBKsdijXysfiFezXnS4jWK4Ck
PITaLK5IqopuFIH+50D8ZgKHmS+x7UmI74tnYXSf6QCbF59KiU2HBaKY2+7T/4Eh+JCnK1bCOod0
m/x7hLi58Gg/yEteItff5/Cok8mA54g8YBUAbDhv+hp/XqfXOZXJqjPkEgF1902r0FegBKB1jfuu
g/1+vlkasLYilO4sqQcDPcU/Kt73mkKXp/yVKnIU/xD6/CtDh/1raj3nsl73s0T888i5IzfmMJ5f
NaUZnndWyVu16QhmoXLd3K+ykej0GW0Q6FVMUXixn4kjO1qwB923OmLSiuDTKVVuBpZcOGd3j7GM
2bmqk6vbLKpMYe0etQRQpXih8jFLzDCVMDxZf5RDh4sE3+yNBXG5poXFfPocbQ94qlyW8AEiodIp
yz1cFOAWFrSXeiJbfgHYOR1d6d765ZioOQ6kmHB0gYkq2Gz+ec8F7v38Ix8CIHzzj8txy5sRx6w6
CksfFwbaIX4IzHPfCFw9k3eVWiNG3VN42cwQy9MpVZaPaSPGOBDoFDyOp1r9bp1LaicMZfCtZiLd
e8rj4ViL2aac81vBQTrIrQ+zmEzfSOEWaGWV8rn8XF+HNskGFW3EmLLvHK5I1BxnN7lypihsEo4b
BGP7dID9RoqkEgukFEDdzf9xE8TreOEdoXnJDdO+JnhCTd0/Ged08pya+ixoaihzuS9P7RaEOcdN
HyrsSi83h3iGTatwCK//iGzLoy2fZhhYrfIcniB7z2x0g9MT8jQMc7Kk6HnvwHKLOXwScqNiVxUb
ptduCQqA2uZweXCaxwTXkokzqE5RbvDnrw9VQoIn/meAHlALioq6x/NwUiE5AA63dSA4Tac4arAz
m8PVQa/3i9o+Kso/CFl93C93miUZkf3eR/ByvGSA/+/gh3NPToXH0CG+xFCajsHGOodDC9BRPlDr
ap+T21dvfB6yh8rsVz9Oe5swGL2LlaP0txXyRiFC8LDiO5KMMG6XVN4FSEq/l7Fxo93zS16uNITD
HcUjfdBDTR6UMQY29yta1+VVXGSX8p0joZWT49pw3OfUR2cfgYvva3mzYmTVNJzVazEqjoD4uPh+
kHQejMoO4kJcJjqXMMldYkIvmUVukP4j1r10BmXQ+m9GhDPdC1c0Ilta7TlhYI7WtJ0fUMBQEYXh
NZdNNEoaQqovdn7Dd5mW6snW9rKeigPDQi+p4MqkYuzINMTKWn+KxO5kSBKfiaKc2KpNhAUbI+lW
Jlyewp4Z7CDaLvt21tZrAQAqzHyzbjpRjBy+Ujgis60U2+BJqnO6XQwtiHlymEgPTP5aDf8fRaMG
J0xxw1z69JoVtXtYxXl+LVsqHe8W5QJkgR8gjucmAqk+BMKERva96KyRQRymAI9EekbsIuXXYsnV
ihmkmpIJQZQGIkhBd86IJH6ahJqksT7qtOWm8H9TDYmjeWFJ4TSVJqFqBkBrRKCPQ89qZlHAcdcr
FTGf0BuS1ilUJYTecn6HPTtHDSTHkyJJllBqx/AiVa/IDqk7s4v/7rGS8IhZ6yW1Wxx+tsVOTuCJ
+bv8/NSQUsG2ddtYVjhHdkwB5g7blOhE4sfMEpwVFrZ86nOWwndkUqMHi6fb0WLdjSG3dQbMj2Ku
X4e52Db0qy9uz2nr0HesRMtxB2L+ONgltMlkSZOsIvSq1JP5DV1sG0ATW4AMsd8xDzVuN/8A4B7Z
M2VZhH++ztiv1sQfokbQ1podaWiAZNb09QLML2zGZcdBg/8l1OypgJnkpzBOpil/GxQLa/IhLTCL
baBmMaFkEvXWZ/mq2ebTH+DAu4HeJ21qV8MyLelJjMtLiABIQIAm9zgPb0HzECa/RXqwiS8nJXDu
kWN3BW/lAxvLZCI6uge48fxD1yj/pSGySAF5OOXNDxQUPuHbm0uhB+ghCc5FcqvlhkGwdBWRNkd6
RSWJMZWrcDEMpUd6zPIyNbETh4gBVRgsknSz93L9axbD+HCN+S/imh/cOcBuk0qsVQ0mgn1/Isdx
zWXOKsCXDAzzTj02TWvnelKB4cWTuRTpLT3SR3lTN2Mpg15KSNsSLVHzzUJ2NtL7cAetkdrA97ga
lTpwpbrYDSSe0/UVYHYpIt2/9Ln9xZu8am8uGvnGA4wtn1AiNWYExJBOS2C8g+C894gBqrWne08W
ToAU4aopglfSwrvVfGmMUVzu3FkDuu2ljnMSVDdWWMBn/5UlylRlC69MLjoA6M/WSmN3zIcKXBml
vAvnL74CbG0DKSh08NbN/f5d7GbD6D+ooXylDOeEP8sWE+dLW8ZLCzQAUr1Q7HAGJe+G2xzY2IfZ
6FIum54/aV/omyjWebdY0xZdrpYCiTdfqz+CQOEWu0JB5gkPgvp6ZeYxWzaOKskP2q4jrur71wbn
IMIgfQhHoSvi9Ir/b8e5xm1KD2zrVKS4uqi6uEHD8kXs4HEEKAhdKcTI0r2/j7a+P1EUzKwdTXMt
O8HjbiNHTfDw1l02wD9/T2HlNF1zgGMDbVykCpIQzkPYfnSXFUx7u8ZPHPZyf350EutMMVpgO2sT
+sLUMn+BCrMibbe3MuN4PwX5kMwfz3O7MS0ar75O0jCOWolUX8SnvknZ4RVmIXqthRXpJOJVb3ub
52AW+4a6tP8T2RP2yXGR1vTA7QM1NtR4YR9TFI3tPCzIKSF1aNEDSNx0vIimcu1EitdhNfmgTe/m
bG3KFrCSollLuYJrCorO4nyV5/CLvLww74SFbtLgoxSp1vLLW0rJd0RIB0fJfXdhtb/VOxOQEz9I
zUhTccVWoxEBQ+F1pIJj1xbkf9lXYJlNeh4yjectTS828my18WjYMbFzLxD6FvgvlW367KcuOjFb
RkbcSLJCT57Z/h1wQuoEWULHfwjTRNR3bskttIFjTWYJAyddm+67oJCPyZEC8rCw/Knra6GtctYW
q8cCyS20j9jdWVa/+Bu6H0U3rZvOcuyESnG9j8MPcPEK9alxC60J6elZBirfJB71mSVa0O8NkOT9
mzTShwgjEFF2opMbENzGksB0FY5lUMsT0teFS3Q7PgtUgjXpfpfX3DkyBa9WI7E4VE0/B9RlFY7G
p+RmKj+ffOPBC3Zp04BeABDs+y/BC/IyATjUfm3jEhdDvfDYYN8xgtNDIIiIY7XCy3zIkji0eoQR
H5GLAG5km4qv8lJFxSF+En+Fy8iunTTNIhWgLhsbQfVunPUp0W8UYQRSdQ0KEHT7QOxOFGcwhOkv
l2wk8oiskMD52cE5c761382js+FJH5JMVSNuboeRGZviyoCxIUPOYiqJA0XuxgPYHzTRqXoyPOAW
kVaB4Wy+yg3qzFiYOS9PUFgHYwLdRqsRglZoVOEcDwb0BehcZ878QxAaawhM7RC3LHWwNS0y0L8t
rcgKK7HtGEQI7yphTJkX8gDkGyyiskZE8N47iOamztGyRGC+dk/S1a51cwruliZspwIga+9LdGRr
QjSZPYGd0wGuuJ9qnNGFFzHfa/eWtQBuR+XOK3fmcBZd7pbUuE7ZIUmIWrpWvYRuHgl0wi4q7pAj
qodq3ycc9vnmYNWJbRTBxVSFFA9ynxYCID147c9NhC8LyCiCToN+cZM2XXDr5lWAt3PwnCKobfhd
3N14WUwN7khV9HWfD6+4qq4gn0lqmWHgbC4UeobI2o5nTqw3QbU4rOuXLzRRLzntrf2Osdr4Uqyd
Dq7I2R4AYtn6obPNzi8D9QJC6peF6jCZQSvc+Asd3B6keAD0ic7kht4erTwkdE+rxRxcB507uKNU
S4NDPnAeWQatSkLDrfMQTbLqO35vVeGxH4WVZqld2VBs5CDCE91GaR3Z6OWmuAaGwAwddH4kJ1BI
pvarBowM74VIKQhYRt8TM8q2ULh0qtgxHTvNrDdsyVObC6nsaCT3R6ANfeilu5ENbwnO4h7z7Jfb
mFMCbLstmC4NBpJDkapd9lt7rOOAZi1ROjDfEPzy7DXLimobQaEoNtm+44F8BQIIfpiT4/VuNJBA
CZqQfoBWGBBrc9X9BppS0NuM593/BS/xeeP/mHADcSNuYPiJ6nMKkXpP5FIoc+lgBKypAIzQjsbg
gtzzgbXgP3ri78KZAaYIDQE2DmqsB6JWcD+QFlUqpFn+7ukcpdOmz6/H4JEyYVtbFtaxGpOkOAC9
agywszuAGmaf16iMKQ62YKjKEXHU+xDY348Z6DYRq1FbMbJTj1yhMyFNOwY4ydLfey/INlUaeyiw
mVKL+VxGdSFQKSCWIU+CuCiKVH7K6TZ0IcyqYiDut2TBnPqTLRQzUiF/tcXNzDK3yqtu09LrRYGX
8iq5pp7zZBMzU77OsZ1ZIC21BxTwGja4Y9awF+kTWBgdpAYEEAzYmCx0GO41rToDk2s5hbGybQU5
CZBsVkBTuwqHwWSmb214A+3FXTnzRBG0/Og6dAYY90BsZ565eQam3C/6ke4rgSXJ1R6yi75Zwpkx
qW+avPrdtyHLaf/boZlnvjBogxseeDrL6M0He1PCdHYCTv3BtGym7ocv6mvJfSSsclbQ+dOLoWjp
hsFlxbtAIXbhyGHOih/DAthGjlV/rc6wGOF2DTLaQhsgGZg5i/P509g8qP7Odshpt9Gs71X3r9Gz
Z4T/YqXCqy6gQgMOJ7XhwJTPJU4xUndV1QcU2fny34XXbYkQXZ+ycMkGhjMtpS/dVwqMhQfJU/4G
LOsmUVGUXzSBL14cOXFDYJ9dhf86X6fcaj7SreHhxCdpnYg2QyEam4uAook9bvSpCb1I6h2jfCyk
PIMDqAtjD4Xs7Sf+6zc0aWGJBhkHDep7dWsIMTsfgfyrn/YqMKU2/6OL7Ll52c8aSRZaU8Gomr6n
PWKhA3gtxCFX4bRuxOEXCsdrB5FpgioZ9G7TCUM5okR8o+DM1sCYgAwkVl16UAqkjt5D/RzzpEp0
mu3D5JMr1/Y2sFCenq2Hd8EBI0qNeOZRLw0zShAVHS8nXv8nUpWh3zRmvSdmGXwwUg0SylxsMzVr
ygIs/5WbvVR04vJbPlPcu5Wjg5HTvPbh1sia7sPZ1EOLQqzaOvz9vB7N9Oe52UyZbZDqcBgbeKvF
sXfvHVifScAyc9a6pugVPu/mdoLkG3rEEx0XAKy2NqpiWK7Fz/JB169OyQsWePpsvDSGEdgE2/rE
mdK7h7broHbmgcG/avr/bX7soCRAuIbyA+nrWiasbxYDu5qNoTYIO4+m3MHFDlS6UgFMaNZ01IM0
G/bSTWmcFkCIhIdTpkcbU7zRhp+T2U4YLz+NTESoDA6ThFSgLO5ZZvSaCtpOJwt9aoqcwZvTwJjR
uxBSeeFj0CL5ZC1z3UrGuh+K1a7jm4fR1PFxak0oHBcCi0vrnFCbvEOcK8zLjtROiJ6y//35bTNv
5LFxpFF1/ZOBYAzebIjysDDAWOhKcwA2p6gV7T44Tj+dFEV3RB9uUFd6EisbDfCfLt9jPt4za2GH
MmQOwOLwmJBsF1+MVthxUApgOifHqeU4F8dhiFRGd0TbObMRY7OkZWATs6444B1++SjSAP/306FP
P564vpV0D8FfI1mtTW+ve8WYP8hj7/Bb0zQ+tDJ19VYUc3bi/VBy/t8/L1lQQNu6W1T6hyzA2vOg
7Zzabf4gOkG1atj16px1bxOhPnPlzWZr4aZNoWnVHqJlijRAX7tpkfm4tMO7bWF8UOiPFC9z0RGR
ejDcy8O79z+hnY0nbLy53HP0pJfFSXECJONmN12qjWLrKsyrjkfYLCTwNdK7TpZjk/kDStpCT87E
ZfmF04S4MyOfn9/0aH4NI//suHM6bKhD0g/J6OhfsHJTuJsdx8UrT8LbJbaPhs9t8f4BEAkQcq6r
Ep5+PRL8+FuTabHmurskdhQ42+AEhR3qYr++gZ0goK++t37+yr11lcHkLnh7qfSXFfAB1JvEKCGr
3yWcCeZe7nhuo7bFz6yIhuDOU3gPL3mTQ/935YhmXSXWyZ8uyT0iGdlRWw2giQRq11aRxO5lRDB2
lGLaMoVZWtmyQqzHu5/mYfd+2NczOgnmCGtU3cYmjP29gtMSEeBOHFESyw/fC0lkxoRS8av3uejZ
AjsGhGCRZ+zW7PR9aNG+GpiD5MAdCibZbsWCZnuoZnCfU8NOmnhI9obKt4Uu0t9AVns73pOLNJmZ
Gak7cHCO88DOTQJlVs0s1PslylUmQjNmBW3QUvGP0LEfHMPfl8NamBs95NmzYOphXBp/Hhe4fpuU
fshcgHcO+mx3Pj9ttUjysU5UiaRymqmPNHrfujhT5ifhurPvwU4wU+Mk5ABqr1az+saC4VCu041K
KYJHvjNIZ6AxusvMV2S7bGw+PiJo/9Hr9Lpqi8AYtyzLnrl3ixcJC7yI8DHfdo0waglYYrGVGUWo
/slJyLSRpC5gFveeaPIs/GRQ1fiaakVxQ3+qTX/O1GYiDrLzq7DR63lIqp2ZZS2VVtD/RlhSo7dY
9ttjBVg7gIg1ZvKhVnSGTds+8ktOcDaoE1OwdF9qh0eGk2w8o1N8Nhvgz5ZX+iIIaPeSlezXCaOd
1wn3E4AFYHa3mmwncig46hkrmedWER3AuDi3HSipxvjICc01vtwfViJJrCwLAGz8Z29Xc8OYwmmf
yRd0R+yt/ulf++G5XvtCOKJrHUmU90xZ+qHGD1TTtKgNKLtmXynatMOuRhc8LuKNQfmAhkqd6YE8
c5o5BeX3W63MN0nBhVBMBWVzA6iJsgd+BtdWFeNyklLySRQkPvDdzyxBNN45n6nZQQLbAJALnrTZ
owvyuGIkXQzwT/Cjd4/pqBhM6KQWgRZcbsfrnleeltUeTCUiFndfoqWCk07DrbJLohatyLbsnDA3
dw4oGpHPK8jgEi4kKA7fhdgqyfesVyp6iu7q5embIusFQhnESl7DDYFueIK9IF2KZgaNjeh7ir1V
VQ+C0eqLnWAA6sm3JOQYJsGyTzNkTYNKmrao1rERhuN7ftwTgBG5HawtDyfAvzX98N89cMZbIbMF
ko6tJOSYkx0Z9LNdGXTBnuZ32FFsUoPvHyrcxKcbm7CBxTPhuH8l7oNtEL1wqmq1btcm5O/SR356
Jf8GJsjWQxELlFLm0o1tpGzPSnOTDFnmEM0i7q7ekdLuetUhbDQztsfckGDtMVZSsJRkAimctwOG
4MaeDrSLN8YowKFFEUOsUUcyxV0+hMyw/dUi0P8Cx3JJvTNZZXjJeo692raHtaYnc+PkFkjzd09/
xU0ldQu+BpMiXvduw0H4wLyvbYFNX9+BMUyQBCsXamdHnsjSKadSANUasQt2f0mOvzH9eDLpRaa4
Fr4OsYnIMe0RXY5iOFHvL+i34atA/j+4wawQU9YuaDBbY5Nmx9qCim/BsmLlhFnSCAxyyqq14PcI
4vjVp+O4JNEGS/RccJ0GOkxPa+6w9RZQdaKaAnUM32K9+Xsvwkm+Jd8/c7ZXu7EdAv0cR37Q70bp
O/9dqV6igbDWgdOT7uQE6souGVuhtAze9J/c3Pghr2hQvTlsKZ8f8jdvgLf6ndtkNlUi7zE4/qkW
PtaM8krXRMBTMMX+dtyc/3HNgvszTkl4a7IBlUxwZW+eMp0Gz7C1AIByT4mBxRXqRf9BKERC0chb
nfBneSBH53FRloBYnsYdNZvlTG4yxDndrUypVqkd0W+RmT2p8TX2nOJQkrxke/ovbyCGvDO1aITF
ueuHR8VWWfJaVS3PPUmAPc6R9Ua8qJfbxQkZbH8hnulj3YMV8wlfeT8TxPfKstaCk7yWEc9M7F5G
RD/D9YmItN+PVCJ8/Upu9yttS8PN5FMrgktkLo0aHlIttzAm9ZmIcVJvrIoKiwqEW+H8458RNqLG
kbzAMy0NgZf9HStWj2xOZIXZro80BiZsoNhUx5AwHWsUNxP88oD5kli3SNntZB4vi/T1KB71NZ38
2ds7uU8ZfhTyk3HhX46Jw/WTvTKP4mgF/NEezO8JKVhD8/6rC621Lbeu0aYhKXSgG8bovk1bNNoY
5GANI6RBXYDK3EGy5NeGHAym70ynbSkKKNrneUCkWW2ycG3ksY2Aon8nExzyN2jLZ/CzNSzzcIfJ
68/a0IrCJ7sT4gMzd4OJ5XB0tFS39dBF/mEfd5iMNoPoUwIW3KazGrZMpzcsG0d1UPSU9i+lKIUx
vF3vLMoC8i92atSLK5eFdyS74NHLJzAhqrXAHiBwqTDQOzsry7a+pas2Kp2ZKDM+5yAFc4REd9XC
3/hVsSevaVsaY/ZU/mImJZXd25zpZbXPkTRvLM7cR0UAJlcCZu29q4Uc0zGf24vCit5ys9Pw05/f
JNsZC6js+9+wnEA/6eyfs8vUfm+DMrIeQ/3umSHW2nv3K8YniBRuWzBKNGaZJdxbv+g9TyLbF1EM
lPi9XWTJPRbLGh3IxY+LjYoGbHYNxVuPdIig8RXka0mgh2Snv/ZUsYXkuv7LVUPLN0ljxxxCQ9YP
rqL71+gcfU+/hcLZ/1RoXgTChZLP573mLlsL4rCN4fwdlN5IR1OJP6Mrt1ijva7tJHbg6kMKpjQL
mLuTN8dbXVEg00rwlM5YMH0RLhvBPIGCR/U8jDUTtNpDwzijaqdR3SqSNpeygfAcI+uKrbWa/zLz
0SsA60Zv/kUxE/KO4C1xJ/cSkHW5dCo2aQC9boIli/AwtfdTWOC+6ZetLujX8CzfaqwzzJhzgsDa
Bpn91lhu66qB5AmFOE6ME6oaC72l0gV3UKiSOllcb7pD9wui8idUUpB+zbZAW8MDyKJA7uhhJYEJ
anr2Exuop5CmOj9SvSe1Ue5pFgLM+n17/0efD3w8miOr3YDF4lIfT/ebmPtO9O+ikBBSkl4IXlEn
c9qKQBbD02lLg/cJFm+qVjbcskTVzxN0dgqbxCbJ8NhoeAE93iCDoYsQf5t9YdcfY1iyzRN34AZY
pLDzvWPSYRJL8PGjFjyzlL4jkxeeWzXzTcnr2dn/XPlR4jmVzW7+dGJyxe24SmfWH+A1AHJYY21z
rKwgw+L1X1NWqGY7dTVUb32r7iTROmXxB3K7B7p7J54djaqUbf+TYlH6Wz1jYZRH5SIxa9TJKEmT
AS/6SmRWWPaWYpxDtM6tr9CMxzKoACIFdjHK6B/nA+o+t8i5rIfZ3JiDG10+vQOmvOy+wCZym3mc
UMemtxitI1pdIhVFFf3qjLXlFLIG6gOVo31iy4AW8sIE7czBIO5teSi1TTiPbQeJ0K1TWIix93Lt
j3rPyHcM5496e1kNnhw3UWNG3J+xsP0E7GgBLrEv5rIBRJV5IS0D2FwhCqInqbosy3pGBZ7eaULy
ZSNIyEOF9OEAgA701rqUnfOTSYosBVCRcHgnaEUOdYXXvficgaSd/63zUCg2pGMZ+ExRi7l6oJcx
9fiFC6TAubkts5Q1cLHAzSbVVN/jX6aY5nOApyfKkIvIl7m8t1WoITQkYyFMUs7yn8g7Hs5MIjZc
Ae8kZM++m0fEY5NWLLR2Healec328brKPQ304t54v9YVQqwVrvXsx5lniX2lIHZt2L48VVK+tkOZ
4fFR6L6WBsCDDqtZ78fHq/3L56sUIO1XWCwrapEVk8tAF0GltX0Er9TqK+lh/saxZ2J1aX/Mna/M
PLmjcSNS4VKDYsFBwsKZb53w9ecF81/8gCNvV12FGz2tYjZxe6Pr8FedQqamBSozNiobPE0SDTeQ
vJir/ldqAOknmeHC0LpSpaHb9iaYfVIAns0pXyPe3q9qqI6tON+xmq4vso5pmQVFCyohxbIWtqUf
Ues6jKn6FhzoS291+xPtRVb+rtegjr9YS3HP+a9b6FdQryhr2CuXsWzanLSQKnv/x9F/WA0AmiGt
/mf9S2dn4bMbgK0a3tXZ6iS8a1cEgzpIz8LvuQnggR2ermBFolHpcyu678z112xlJ9QvjOMdtWzm
23VxYy5Z28eD4GgaJTJM5R6+sJ4ysGMiuCNEEPHySZHyrgXonVpwZ7iJwBE3/D9omYuWPL0zeIQc
FQ2bpe4l/YMPWImNGpGjOwCH2SEAjSyoLosBIWSDVyZt3Cs0/U+jNhZiSLoKJJpwxQS+jyu+5ka9
jUpzEja2dN0+myUwUv661fPPoQXYpZP4e2ThRFcM61dmynhmwCn/7JuIL6olIL0rQK2q0TMesgHZ
OHixD5n92W21gqZ4DWwuFU/+1ZNwLAL8swaNJ/qqKact5O4FF2lP1SybIw+0aba7lexRO0WhQLqP
dCvhJd9/tsAdo8lJLFJjl6z5aHZFGcjDvvs5FGvwWAYKqkYDjXq40zfuMQY45XSoKjcRSSM4dWtj
Cmu926E+t9yYIT9uBCc8lnn1WinuNw84ktXn7RAjwFM9RiHsMRflTuKc/RcZHbyIiRcGt+DazUEA
GPrOnx5Be2JZ/8USpVniyu4jk54+wJeis0YQWOhpl/LxA8QBoqAaofoECgvpfTGn5t2JU092SCDS
/VRPDKPb/enbV24nk7zD2vebr2du4T9nxb/YNZKTuUrGI2/2ASaiC3RKporg/2eIB4e5DuKb1V0D
segwwZmbjjHTd4cuIIs00U6UYictZm2ex+BrUcoLPEiBf4oRygfv4Fbi5ODnz+9RkEXDbP0MiIuq
07383HyO16SQIsbpX07sQV8mXEmJJNaUcTNa2kmVvd19nsIJkQ77SAJGfpGFYDmMTiN03UZaaD7b
6wUv/HTrKuIVZLzXJmW6Iq61Nh+uNGfr783BLQhaM2tpsijn0cpz6CWYxlWZq1Q0rhObNPvlZnUc
12xAMlOGcyXYSXMhRpej22Nz7CoZxWnvhAtb53xii3PbqP7TVm3p3axMhmk2KzKCgvAcIEKoFwt6
Aj0+EPyyPF2tnrAvloEpF9avfIA/8urKAP7tSqdHn8juKboTpkzJ2ISb9LCNqtr08fZKEuG5avR+
zT7chHZmkeIi3yoNIc71f3Yw2A/Bdni41EYOyUkkFdnafC0s2BTHPOvDS4E68nwqrux6lBT3H7U3
dqwrwZJmxlqbTMinAwLmAwHbTe6n4RP+kq4Y62wvAX0RigGWEw98xMRYkzRRPKFxr03ImtAApWW9
uqRrykrCw87ltwmtlZBq5k7EP2TawCFERqq3AtB3xOgZz54qZFRRIwNBfBe/IhusrG8HaQTbkFkA
j1CxTyfKLTSjG0TAyZPs/h9+AW54Zq3ZK2oRUYz35rpRANDNT4tidekjW9D2kxDWtDxI6t7083Hw
cyhSePk6hSHMKWXR9gfDCz7L6qRlnjYUAz6Gx3Ao2Iazvb6dvG/BtHafDRXJbhFzo55bJT590DbH
w0M2BFSGhXT8/79wIyQhu1SRzheI05db70fN+dLo9vN4rgiu5UH+YMSuDTTJiev5d1lMU5ZDLgpJ
Mhe6yHKKOJAbjk715VA4Jon1tBocaX1cnzVjQxA0dNjecHWzA8WMs7+IRumGnEPSBocs4lchlx4m
o9CdEc4AUV/4sbTUt9giIGoUeXr6+e8szntXGB+XtzwFp7qNQer8rnMaTH811CCgAqJWO/xxGVMH
chZ5hjxfoypdHw/7nn4eBeJXziLIAa8cQjKPgzD/CmndZUjqbPzxX6y9qQAu8f7zTPnKF/5i2S3f
OYCrcdqfK/zadiv46vWaHbZS1Mfmvr/F3v2Hrt2TfFTBr5WlP4sf1Ep/n89Bqq5ZU1FJBYly1ZLO
OdLs4ATtfvYHwJnk5hyXAufRXbMLfO0r2UaAtj6pvYY8iFq5n5/Q8lEdHm6It2IgYpbR9B5yF07g
UM7yb2+pYVlNS8aMEx+WMU7yaiD3wW0CYU8QSMIK67FO8aDbbir5EaAk1k4ui8HhICC0j03mbw+g
1DhahjPH+uon4sQtbmqGAJmDFunHugPxilwGwxD+NC8G9dWIwDVCGeUlGsYtxdUwO8NumBLmYDAV
jMWNuKSj3pUHJJpJZJHNnUzW7k/n3I2KjeIYdOaqETt3sYWUCtLIz7lqih7AVOcgzyH+8cjzJTpK
ZTIZRE9jjZ1iI/lgSGtCCygvblJH8WBhoJf80KhzRwk2KGX2eDENef3ZLmt9I9+dcYmPuyDSm4y3
1hfkbiGHUQevQILwB6PnYXbvg//6oRxU7zTHgDKyZ7dp4wGJ0fiekKJo4exbeoeIx+POrRI7ql6z
+cNwtJ3fuyChSEgAKU1fdcabz6NiiarrItPcd/u35nItLRmdXz+2qryBJuoIFO47dqKxJctwM+VT
C6GxeHwkpRdY+VaW2/QI/i5KrK5p4xmha+nEMzmghIDeEe7GkWMjiQeMjnsM29OO6JX1IcISt8NK
JQ3a3cxOyHcShIdF4ltbVdfhhBJ9dgFMYa/liTLd/ZvFM5LQS7mkaYiYN7WWS5wRjbGMNWnvH/Eq
hQcd9hXBuZXTm6/y3L04EZzC28phUZQguA3dq6np55DKE+S37FxAG8rN10M+dLOaTq1VMrn0HY3J
LMF/NtTf2vqarpca3YZhnecPD5ZQqcPZpuV/0spmL02tankQ2dZo8R6tJd2sWQHj3/By4fzpiaxq
cTzeCUVpFN8ZZo+QBwZV/cDTX3ycjb2Ek3XDtNBtAdUULbOT3HwXMPqz2QGh4kWn5SNecLqN7gjd
EQl2TyIgbMK3DH1mdrJRxEdzbs7ioSRtFczuqfw2sxOghpt23YnNUM3M7CmIMmsJh3X8v9tPrFl2
KyH9Txz9O9ozU840SwAO/Jl7IYHshVBuaEWvtv5yOzhc139lDHN/oIAVQNECCzLK9MRi58+JStwD
swh2s5mAGdlFzUhgWc0ru2T4IGghC6Vqa3kVx1a2oMv9XrxSdzRwwOnAr6OhaDKe4+aCDKhTwLN/
ife2l91oSymkOgHXEAsOnFdGI+2Az0l4dUHziOeuR2rBxqi+pBhhyjfocttM/sF+7GDi3nrNu+G8
YrEzydcICUGvn2EQAWxQDIbTaGLhizNuV5U93o3nHxBWmBsVHAVA+LmuI4IGkz+iSInX+L098QiI
Hxwl1UsdHFPAd1KgplBJrKnAcYZcnhiM17DgGSKtqi/XFYZv+EyaIo/jmuaok6KOy18KnfargZBo
vb4zTpXXXp3mMvDHQZnpyqKeS/scWBIqP+UvCoXdDNyyuvHiFSxRSPiLOQ1Lbk0kw3vhpqD1LmyS
G9Arqj5qjAXbMyt7frWjerthtSjDY65ZSH9zlI5uZpXAOkXA6MOTEALrUe8L8sNs+NWSpt1VPGk5
tPuixBMkgab3ci8OGXO/k/iiLxSkrfAXBN52FadHIKbR7HcJbGqOtGGkJOHvy848co/5RB2mDaHL
W3c6YKf6U1lVnXV780CPAzZmdPLk8w4OaQPG123uTC7yEDoE2aPUpsquAPTnssJUMQqWJdScrANr
FFxKyZYfFIFUw1DW1NmlSwzANv2z9yAGOr/wfmm8RWBjze7lFsgitmOsQRCKNYqLhfYIxErPFEVI
AKkaJM1ji+AAFyRBv3BNUFZd2Dpe8MGbjbdP8j+xkACD4H0GeqgT69k2s0Mc9sJHwehTu0arOh7b
z6vQvv8G34Ngpg6JNBSBnnVhKN4fTVTIBpTWU2TmOgtzONoS/SZzmM0Ccaw2MkuyF+KMD7piwWni
cUSXlIWK8XrMQq3GEJohKdxITfKsY9CaaadQmS/cCJYMyNE3eu88EwWlZICkX0vOKmlKaVTV15iB
SaR4yEIiN4h4lYQY/VPOLQ83EPMQSJced67nf+FoMnB+/rwaBfc2Ecdjc4bEEMKygBTKZ0lJO5iR
Ww2vDWECoLoIjhL+RY48rnCXHBn3AxBTR9OD4zA7qvA/jqiCzD3Q2wRB1Tz4ZTPU0flmPY3SN+ol
b2di8nZaeB3OI6Uuuyhe+bWmWX8BSDYiM7yV5T6AuKY/SRGNkInujVKNsdq7MFe5jgMB618aBoGI
jnJJjNSE03PEOqz21NFZuVRdP62pHkpCrmfj5DyHCUSKemudmRoqdHDNX+TnZodnAas0jWoxOOjV
WFmccn7xzPYb1yqvcKWAxkkTDExYQdyHbOg0j+A83yZh+CaTTNo+Yy6Ok3OMjzFdPoCK+UGFePoO
pUyOWSJGAueJXeKPNVhdiMVnwx6VxPvaN2LwJ9jelOjx+6m3Vzl/pO8qSF+kMPu1PQQeOoOaediY
XDFLeV3hwnupIGfXnq8VtefoC5CU7UvDNRA12JsmelvO0zeoeKI/faJr0OtTXs6wyzBEwNPqQPE+
lMoE/8ur6Y0g6Dsv6hQY8/rnItmBo4u/6TKgjqJ6WJ8gO1xK/a+aWG7jS3PvT3Zh6AN+TI5WnrTB
AjLUTv1poiqf5PlNjUFO7TaGUe+86+WH9XBOLGtc6EySYjpGSGr22Ea2H96pwA6z2nQY95sxNgo1
als17HkoikJfxWLRY0rkQZoL264nYY1I2A7tDum2qbCAW8V8v+TmlagrbGvf7pS+Mb9fvm6IzBBW
NzckSqg6ErGwSJps51LUjvJ5KrSITDBzQffbMbZNJkB0C/5smRPAG4a4mO4b6whNeomxD+zAryBa
WkAEHL4Llempf5BPDuHtm3ChGyi4Fvje2XDir+pD1DWr5f8qdjOFFL1DgNltoBGqOA1dX+kl0fQM
zK/tOcN8Ueweue9it1vTJMB4cPDD7LAq7lq2dP6bz9US8vPU1r/KUld66fQcmcxnzhIMKSXhXVXH
5CLrdt0Wx5g+tI9ooQPcxfgUQLM9RI6Qx7dhEQbFCv1xOiRMCMJPbKkvbxl5BOQxxp//VmgI8Rbw
n5Xt4pie4id7OHHJajD+3yvmo8UF/zB/X/Vy6+R06GOlZSFy8hjvVRCX1xevnKIKrTrMXOfu+D3W
EKntDzRlUgwtD+su+CHffb3VtJtVEdg1WB3eZUzfqTJ2qYz6/dd1f1+4GH2k0Q/ETufwN5i8sDR+
Ye3lPSHZABxTneSS4lLcm1TUMXaOu+6PqVndZt54uFWpPebjqTfX4sIWTODRcrZD6wWLLpfhiham
dzMBHW6e1S/Gp+QDRsvVn8d87QOpOXf8B36oDaZl92RnyAeumZLOykgrczvb35XKIGGtHD9lf9mu
bP76zNMTFDdjxXt4kgi0w+CG6RhH5Qq0uX/Rt0Qx9H4D+Pu7UPq9qIbVAU7mOSln/mQGr4pZPA9q
LGxNt/SmSswSpNioR5zv9ALvZ9WLTNi8p7mz0/EH78iEpgayrqAyH30AYzc0OVLqG3FdVe8CFsrB
tlyx+C7eMT+PxwmTa7xC7CdkCHQmcadvG5j7D0HjfM3FyktIGd1zFwA0ZXtxh1+qWDoaPQnUGNua
xmTq367dHleNJ0SpjaZ1l2r0GSlwmin1LIM/cZXOVBuPgePmz72sJlyBUWpSm9xUCE2pVbsmz5a3
VKDYzE5f9rCThphkvD8stoFNYACRXak6H6tvxyNWV6KyTohINJXV3sVgxrnyzLRH7cryb8JHK2Jl
uqDcsgje9O69s3qWrvT5IsbaBqdE1E1PNEiy5FQ/KdMPe/x7w/8Y5WudYuUyw6gxSVYNoufwf0NF
0JTl9zwoAj6UHdjXXlAmo/zDKkVWEjKxoitNShSMxmykp60fom6duGkMhz2SfCqfG2HEFfvNsDD7
ELK13U9B+OzKD3cRpNpjpMRb9/DWNJkIV9QH9Or4Svk/7XMOK9w855+8d1YBssbhqOCL0TfZI64T
Y62aWs18TAWyUVotlCxNoulr13EEzOMwqBMdXdJgmoKkymI4fzZuyungDPaIqQNLgR7fyTWj1pfI
v6Q8FCYbTE3MWNcfkiDECq+QpOmwBE4j2OJzJEh3Cf7DdD9ykPKJzwq7Iald2hqmjemOBEhQGMTp
6l5TNXF/J80c+jyugdiizb8jCLvLhEgDzeztCF989Bj+bSLmpksbaa61IDw8fzxhvZV/N6OzvvdW
Rg9PTvPedT7DIzSm4ciIAJjxxrabX8gq1nLaupAgm8MHV9yqpFehp3geF6Rq9qWUacxvEofQOF/W
6GR6qs6BDNKtGxLg6UW3sSb7hh4pEbRXTgBM1MnmJPX3andZ3b1rcT3WxP+p/w6AlKoNOKJJYhcD
KzRMZMNwOqb3K9Q+oK9MCRv7wVjn1CUyGgKDOwinpMMPgGoL7nMTIAt/FkFtzAUYeLzHeGuTNVT0
nHYyZzw0w9sVwXEOT2AE0NQGmCMlw53v8cZoHvOPXCTwcOlt27RmfFkZYoixsb47sZD0oTxkMXIK
IPSqkWt9HmsAP0lTHMya64BMKCdud4b/a9cEcuBQ0YInqrB8a2WUpG9zisqCc354wjnvz34nRgdm
qHFCmHmKCSmSoVTKCEj67qII6VoUK2HfdNElnwJ6oxfyOz1yWHmMjf7l4wci/lfEEiAukdF5JQnD
BRFgehh0b1yX8e18AWrCv0UKBNhsrWGIFTLfW2+OZ9m6qSv3J4gjtETLBD3RuEChvLA8D6JxNsUM
f55hFhTbNiOneVjZ55YAE8Qyogs8SOZrvl0e4xALoyDthh3kF7f0y9uQKRf5kG6AJy4jIL+srLpS
V4BLg/sDGpt5a63N/BViXO4DGeew7Ml11bYB8JEfVj7Ndl2ri5J8ZTdzkSgpLvcqfYFNP4Z1SwLf
z6m8N7wpfc5uEAS86YEpC4pOzE7nDUMxaLp7AJZn97zAzzjQrIFvDfIjYfZ7kXbQIngmPKVBXF9+
SnMrH3aIEyqkgrQexTRbmC6WBsQ8db2qJNlA2U+vnuP+WMrZeX9MWczru0csuFRhFNbryzlutSQR
Qpy+7xhJEezulK37H5W29YRxwjv/xIBHkY48zZ8Y24UlQn91DmFYASSJr28JrcVOyspxC4beCpG5
OQdZ0cJHlSGPxk750+WkiRZs3tUtbLdPWNNtfmpRBasRwe+llUNecMwkOa97D38tAQRxhKExvzAC
e1Nhf/uhyACtdKcz/nWY6gh6mo3fWVbkrsGy7fK8/T0OipTFiLv8wxbkFqLLyF9whqwQLzcKEmFD
dcjIopm9dxf4MpPSxcceFsk6aOTDNsw3BdGRTNQ+aqzRPFxXPHRGH2nt0lBx8TSw+p+gSFPD6Z+y
CehrpIDbfnhsLhpNfzTFOtakWW3lU0wZ9Lofb1pZY0ZNcTRRwc5ETe0lmnZsENJJMOpStxVESS2r
leMuDmjoFEZVxQ0KjTMiIC4LQjfaIIuzKnN6qvxzKPt9cEAWdcv6pBqZ4D+CejOSRhxeucwA3Wqq
16Ty06joxH0TEx+UNWxy5vAhGVrkkesunBi7/fnEYXsPLGxUZvLqU23IiWx/oyL8ybG1wMNnkxXY
eB7yWRpxAg/ILtUAPKA4442jieBE0eju3RtR3JR3DQ3w017YEkbiHQKjkS/+T++l6+PgviSfPnXU
Jk2/hASAJEv9qjvJoiKFwd/Yfmd/Mxr3HZ93kQX135Hgjo1I7fgUmymslEOpPZH/zQe9svw5tRCO
j6OwoL5bp+609dTOCzPqD2v1BZCtoaUi/Kj3E3/p7krsFCymSRozeSfORXItflrobrE6f4sYzP4p
7Vw8SSOqMgC3EM9G20JuN7+MRPQl6hnfkgLKWK6gjh5/xJCxqR055koJQCQf4F4usbeWTUoHC1a/
NjYcUIs5P9jtT/hyAOw2objY72vsNsUMPaDSL3JgY8aN4iCDyaX1DeuNstMluG/zxlF9j/WJ7gKL
+bugzqiLuv+m4upucERKRadSkdSd4sm00xr6c6lnxzaj41B0kRt2zlFjAg4cKdcvtkL9ZfFWEyHs
Q+l7HMnT9mcCP/uUSbDwvfXWvMhq07ahw5wMMjPlzxZRC+6WQBzk9LdzNTL+IbTOs2eD1gb6GXyE
8PubL5aLewg8nCPr8BHI6tJeuigMTRYBAFDs1hMv7BgrQSpMKVN7NO9LRb3jeY0t12NrKMjY1PN5
NHJA9zq39OxmouYcOBtVZTGjBY1qXSlTmqhb6Gxr0+0+FaWu10RCw0TfDSAMr/Uu/0K5TfqK6C4R
m3Q5rHev2BF0wRcC7vLmy+4HSKcKBRqleDb2F/6xQpgs/Beh35AOLULDVEVZAXIIK6Nn+gS/JQTO
JaSO/eF8oy7lXg7Z8yUvwyCFaLkgeUVqISFDYa2Ptsys2gC/CNZm+5dZMxFoHxB8sp1CZ+9gIeGq
HQwvZ2lIrArqLoV/J5HwAt5CbE3+4zaiKp5V71nsLUzLFIYjMnnNCNtj0YhgcrTHuu6YchYzWmkf
zmHqjTKTDrTlI9Jl7wSCszppUZb1j2US8eUwa0ON8A68yY/xGR+Ar7JAChc/hdz0mVZH2Jpo7D+Z
q1vg4X3nhThpGh9W1SFg/FhgZ0ueIwesft4/VebWjOtsMTz6aPMpktglZrCawVq8Jzo6SCbJ8lvO
QMEjmUJ2QrFtuOOGwewmSHGWywmkVe3BaV8lxsAHL/fk39vx7dckFTVyzE5rfHyWE/6SyGT+kT5v
i7ALCTEIGPT8A4NI8Zlap6nFnL/jPjVJ82+rQ+1eS0Tph3mgi8EdN41kwk0HRnOi5zw2DBEA2lz9
Nx0ab64ZXaPa5LOPri36d1wPszeO37/zuIS8yfWOVnbLUtLhsXqd3v+QbBUnsag9g+s8ECPusVAt
LfjFWloUkxXuu9FTL+wVw0SpVmoFk2rHh4nlRhF5F3OLAQHOOjVmrf4UxFBtXR7UhfI0uSH0xcf8
RkCyEilcsFdvh8xxp4haS5GGlj7ANpH04mF29Rr24fgbNcfndwPLY5BISBiNX5kFaSUP1MBtmej2
qmcdTmneAIEF97DlwwmnLRZ9GNyR7xcPtTv/HclaQ3C9IRTzzob/kMIIdmkUKOzWZ6OJ+0zFbi01
v0Z22yNj9lDGyKl7im2e6Afs7yqiL2PsCWTse7XsAZlzFSz9kqFWzSgwoOjVxPE2o8M5YWqnug9n
IAYlj6n8gcp/SXPriWO0zkXW6Dp15rATLKIwHcyYDHeTlwPMwXceR6DAhhdUraRolgooAXhHMFUg
DHfVwJEULMHA20KMBUn9ABvQhBfUCMBwySI3RF6RiugvaHAVYqM7QFO8YmiZZY5ywugGpd36kenv
yq9b5YATaADRWQeMNjZc6mN5Nr6DTPy1+8i1rVFTw6i9wEBW0EsLWoaN0mz6lSSsrzOvL7g+umtG
ftaNGVkMArqdlpi6vPsm13yWw8XTogzflE1on9JdWqnrT9aKwbGzecN21BQAzvzfBdnhwQoWfka+
PXuqIS3aVb+tYKhkT4qM2aW8PTnc5nhUNJU+O6/1Hke8LfEVd3zby7yrPh16NG3YTkLdE5QdBCww
9j6tGsQtg7T601DVUe/QFYpmXy+s2MBX0ULhem0MJNLBjZhnwJUgSv5o1/PWqWHP6lhCy58tY2sJ
3WX8OVLTt55rn7oWqbVxD03ObeLlTdtIo6YbtlvwLbOa66Rs2tckVirzWp0dbqXjY7NwPq1CLpzR
9qoqtoe+8/e1sn0yGZiDEmLlSaDQWYglPLe2N4JJh9oZh4yiAMoTxWGPxxZaXKyK86luRuHsXGh6
B5Wy73MOyXsCuaDmEris6kt5Sm967mOywV4htei8ps5JJXFLcPWG1h6a9v99eMuMJ8axnWbWCJHn
dYsyiqWKM17bLOBVbxeDVTWGL8fndhyQOCfJy0+oXHmdXLdEbuQOmXvlDKOC2tWYmCCCStIBQE75
ZUMC/lRvywlQn5Zz9wX+ieEGLRfQXGHD17hzoUT6czr1uSn3uP9foGLbfCP7OurZd/l4gkzmCsaf
iPZSL/4GBNJA45Mdq16F+RVDGfJlKFmECvaxlc3EXoevxJB1WMgB/oAZURcxhruwZlyDADxiMhfD
LaTDuzcxJ/UIPFexkb3uNghP5WlliEEbVXsgH+ifSyAaOgv/EVa/APToLhAZ4yqwDVS6VZAUW2I6
E4Jf1usqCWAQSMU4icr4V/GZULh0pOnlX3g6gHiZB5rZArMqNuNLX7o4MUgNG3ZuFVPC6qBc1pYe
IlBhXDfsw1Dh85U93o5QGIlTYM9saLgQYX0QG+M910hRIyXd3K5KMPvO7dOF3IZ/bFFSqpRIsP/8
oFE3oF1hOs3TWYgFy2jB+Zd+QtKw4205ExmgigIpP4fbRUHUjjmgFSwi41WR17abwRhwqm1LpN+M
aeOrM+NRaYYaPOQbzblK0gG0NBO+gzziHvYViVRZ0/q9Hdonr+LxMMY866pQj24PCNUGMq3FK0w/
0brwgQrHSgRP7xTH8ERYzzDgGVpSPyGeLbELX44NBCBkdw/zNacQLaXvt1VgiyBWnDmevDLhWsRn
bR8LK+mEoyKAEJIdNuRBoQ5vDmzxYEZyBxqI+eLMXiZihmdJFX9+U+yDBVh1Tghl9NZ9QLpJf1++
o0WpgxaaPmdYBy0fzyXHMJgOtyMcqChnv8IPTVlgv5yOUk3vJxzZ5/SCRGvppv5+qOynQhBkCUfm
c09lPJUkoDVDQxVUzNQSKxNG6pCgGTKl907ivCZku0RPmYO7a5AauQu+DewgCD05nSb+w1uPFm07
edL3nfwDNg57FJNkhtnRkGfUAOEnIL62AMe0P6LBDjT3CoeXHvKkixAo7KaADiii33kHauIAkyxw
vlCVe/xM83yBYBTgQCMLGP3I7pOwmBaMeqILXiQ2cIDjjGiMMn0WYa/R/St5blaBtLMyImgRb3+D
zjptXK6tpboq/OZs51njvKuBnjOUyAZHnYenVvrzLos+N5RcCo0r+F6Qmo7cnpLThgm/l5gzfenX
LG9kPvGoO3rLSHWHeMADrLRviN2wwjuN0hwFkrB0Gk1lAFuvoWgIDOYYP5EK2aPV03sDpgB4s/RB
hl56SK1IDEJDqQeuX/2uIcZyZAT9NcBt4V8bGSN/ITRONnqsEQCgnH2p6dZZa6gBw99Z0i8Y8dVC
GBuUGhZWswK4sQLIuY3caBN/KAtXOg9hM3UbKMcapKcxDntl5BT3DZnEo8n16Sl63vcCuV7iCGDA
9wJbaby4lY0yjDegehOp/Vl1ocE57pgYKqWQGiY8Ra7nWW7p+cNkbsP+pUXe9ezCmNHxsejHYZ7I
5dnjNHqExd86RajRY9h8DHnNLtw/8uchtM8rCbq2JFwLYr07o4WpHn+Bnw/9p6PKEiMJrFTryeBd
2LwC3FZVuppYAg0GKEtV3sq+kkr5pe08kONazMLpRBVj0Ds2lNtPBlgY9UW0ZvkJaqBNG7NZdBRU
Zg1LjqenSgT0jvZ50jdL23GySsGhqEwVVrUmFfbxzAwC4eoPlai0JwX3BxTm2P+FvxH0lmfbRBU8
JPfePBl9KEc1XZgPOK16OnwYtmmf2Z3yhG2BEDgd1cUQFTATIiz/KjyAu9LEzPGjEr4c8AgbhqTO
cZ3vZ7dlgvewD+PN2vpAp5hb3/OUpaCCaYVw1ZP+aB1eDaYKygai+bAnNjeWWNZLxYHB8oBvYLMS
Lgl74rkOdPsQsVbsxyYEzohqPigFqYlwacCujAzG4gYgoxuom030CYb5MjwEQdSaqPVLiyzsiTJg
qqFgE2jzGYei6YYXvcg+5frDdTdley5WVPputCEsHWK01RWj3eOIdXuUinsVeXCg6pzFQqNvAHLJ
DmAY3T8Ybyixdpp/bts06dmB2bhsn9Ucja8oe+555H3OLLxW8ZtL60qg84UAWTIHmXykz790xZrx
7tBvr6E7yMn9EjFms1QL/c2JvS8qSGduY+rMhxEdFj/kRmaYM99de47mJit/+RFjySC4+X90RABY
ex1SZyrWIFL2J/eoXVctH5Ijq+E5KCTt/SogSJb83qgrrlzT/kPuCNrRSRYaOtr7C/uC8iuGecu6
ne5HGnWNztYVdr/JIHRrMNZmLxTyovmJYrBeqb4/OgTHyQZl5E8v0ab1rCfaQzqKEVjJmDWIWjx5
E8VxrQBCRcsPWeyELrFqG0IJ4IxP/t7fzDUloRkVMR542GULznc7fOi2s6IPaAzqzFI2BsMuf+ns
yhcjhbBDU3AoICpWkGojnLNWFtSRFtjRdN/r846P9XHTEHMxdt2XmYkRgZROV+/YtCwBZ+Et5kLB
3oLNDn3GvUUfdclW/Zs1WqEtGJytyVuRRs63KPMRzvQl5BElXSqNZg5nAld0EAzYv+Y1Vk16kM6p
3XJHIQ58TkHB2jbObUcDSQHNUfUUrQWZMnffvyEQGhAGuRGXes3Eb5pxsZ0091H3LbWZzgf3z1U5
6zxge4cj19q8L5YjDqfGPq4DvVDVUZwV7h1axdrBRa3K2IJ1I838MriPC42z8MenBJe+jlfwyH+W
kAZ9eiZPW2Bow5WvlwWCpaAqKlXDhOzklFrtbXFqzVVqoxKFGcS6VDzZ/gozfa8TItDUclOBZTTc
35X4oJjnH9dDbHuUNGtEUYrqiJ6shKvhu+09Se17ZRXjmCTjM82qTdVwvkI0t5zNpRSvY1TP5CaE
RKYxEMnrb/qw/UAWxLows7JU4IAXqde72vk1BAglVNOAdCcx5rXKxUJ/y/DmUPBv7//ER9U3I5m/
7M0zjeFoWS2idFgF+0LtcwKDVYloaY3qHDKMmn2sl4eealkicZS/y/X5cpvT8cs1aXBVGnutX05k
rscovCP7DjklGJQ8GyRwv5w4J0bp0VtYm8AAArNGYUIOofPj+Mfm6xuOLVdi4OBvWpZMu7xS9Fvr
2wp0ho0+bpPvcUxzInaUX0USfbLYnaqipIyxo8t/ksw7i8P+pSgK0w17hg2yKc4DyHf+VY+9udqM
c5lf68rss9U+9z+AfY0x89wpUWyI7LBnOYL/lmcsEmL69EDU71uwb2v9vAA960ahGu4prx6OWyyY
YhYKndWSxUdrM4RyrXCLzZf1kZnwYu5tWyORejjsi30UKthADvljDtpPkJ51Qo+gmcb3tq0+mQJJ
WIYarz0qLMEY+m+arVzckLfSXX3hnWcYjzl9uBdHNbmBGngBW0TXq0GBVsSjthxzput9V91Il/ab
9VgUz36+JduRizjOH0SgsjCjod1yZRnwUvf7JHO/bWyAK6LnlyezywDnm7sfZ/owyEBObVjvvIRm
HfEIiRIsJcJyIZpzXHj9v5KWOx1xZ8NpXnnzCBvumgP13LWiuMGjZkcW5nyLj2Z7JtMWgV/sVh2/
e7WvsKVfXoZ4SlpIqR1TOCiEL8nGTjvntJpFplkupmjJdrqXsVoDr8XRgv4A/I7nDSkDDZjIrIFt
5rkJwqNiYhGff4IV+k7mCLisDy3GMzZ06J8jyQ3JU2NFd29QYIUL9uci2ZKBpvivrJTYVDwHQG+O
KPV9813r816fkvatA13UiJnXhroUehfJCF4JobLcHU9rZzYDGdWrNMLuZt3LblFpJrmRMR4e6Q6c
CVgSJg1MVPR/L1aEGPnMUdNPqbEhK31oAQPpJRrp4nLrw0SpvYg9t89b0EFCdGZm467v8nq8LHbx
FxAQUvfxyNoXeGijqcJbWqwD3Q0J97Wj1Vpes00Z9iG8bf+WISGxY2p9CZqBKQ0z33Ij0NH0UDS+
mmp5JqYu98/AplRWIThwzxYdnmFRK5cwxspxs0vIyyzwvrRrE+51X/wxWEv1gFr8oElyg7+mw6aS
G7+VG3r4OT55WKRicwbMG5jbfJGxfQ3LWX0FDiRmV92gh5gXUcKUM/rMj3cuSpIyAA55Rf45xWDC
9frtahkUw+4IrCs9mQQZMp+gbsQ3Iuy0SAJuuUUEcrHR77uhK6Y5ggoU16WUHi5VDTdvgPim+0gK
WN0V9A/07KdkKydnp0vVxaTYR7gk4BxJ3bHnok7OPlFJr9jwX4a9o6itgFd+ufLyT2WaNzaw0ncP
VQW3vx/PkUuYrBTq5s8tvZGWUuVWwYYoy/cNo8RPWeWBRn8cq8HXlmwmK8oTI8n3WuSx4VIocGqO
Z5zm1a4SJLXY9FblYXoJl8biY3lJAwPWkZW+RDTqeNbRqC/s2hYk1/0+ThT2tkhFcRBW6PTAyJ3q
55/EGq7w+/JUWTfOsTJIVSX7IxUFhL9DvcloXCyVnGK5yhcJr9d5/JM54IP8R8K9Y+wzTSj/XmHB
JbBddmyD65MUc3SQwi+DN6xWwlsx4NrkjopEnH6VXXAMN+uPxXE2+TGQgdk89sP5xiP0NxXcT7D2
FdTk7UFvBRkArV4kw0GXFMe93Jwqf6uDv/Efo0a+nqQenZGILdc14T4KCa/7Ga36IWpaHewNHuLw
OqU7I6ROnCyfm0/mLIxCDRMiUwgtIK59R/sdSoefW8pbZllJHc8JJvPujHIZ6wFOZ12EPmosx46q
Xtxzmddlbfw7eXOde5oH4mqcoOs6AHzkJCuBvauT9SrXqBr/Uj95vmPSQE3B4XBqh54QnuzcAiiN
/7z5dDNxY8/gmTzois2Ovv4i4qlhEzNjKtk8Kd5+EiVjwuRC7pOsn2zvsQrGVGdYqu8XJcYmdIdy
c9KA6z2Ke/yXvE3p0/YwRvx6oHuNnBKsCVo9uusB8bpUIyJkmsMG5aXEdcosaiwiaN0WbmN9sHk4
apNXg3OLxox5VD60agU6QFqx7e9Vt1oBQVT/3W8CUUrP4JHgq+RjvRk89jizYNMTLvsYlUnPoQkf
sQKQZ+vyQxVnyC30HxBshBb2wysrXWJXFIj8olRjRFZQIIAIGJfpyf/XflfWumjNrakqxRGug0Pi
9KxcpmeQNf6p5GVS+JEjZOUfUvOn/GaEQtgbpKU+OQivQXQlUY8g8NvGm1ZhqwPsKrgXe76tF2qc
KnP+DjOPelgkdhP7auUndotm+DgbEYkDg6uSFwJo3hd6AMMS5rcQanof04FCI00wNyDC5tBAjAEg
R9+vsjasTd0URpKVc9fO7m8Yxiu5tFbuOK9g6Jr+BxW2z3h59+ysYMGf6B+w//5RQurRc5DrFkn6
mFA5O/CGbIiFr13XITJyMGiyvJll0rjzI0p2ONZFn8GSUGpW0qE9GDGWmcX9f5592lGq1YI6AyBB
cVVxvd5PYkPNGqlH9CVXXWHLwfRqysZQeY5Pqx1cNXzsJzoI6Pndt65vWJ3sOJgvTccslJRRYZ43
AGg0M8MsNxjccKzTdf5vmQJi7MrTF1yhfycXXh8TssWIACa3FH8MjwpLLPdDla6xuqSi08nTQStL
W3qMsXQUkWYapwnNMND1sZUcVJypwprfIjOWtU3eoYChltlVaD4W0UgO/oBkCx+rjd7+vtSpegT/
oMaV1ZPJoGf+iJVvDKJvR/kzZKDZkAX1o4UaZyPqswpjTOe0cgigz36A6DpzWy8tF0IUUpgzXJ07
aCbreCG6VPxEhGYolWYYAyCzrWninVvVso+1y1QDykqj8qbhvfnDzVXnsgkGxv/2RTkm8eww6EXR
zElydBp2WNzCZ1nFHUwnSqGRC00gpLKWgypKyj5ktCNKpZRdzxac4+h4eWPxGfcML1Rv4EBHilQH
RMD6kOJu75hpJtANlqeLpSV3CDOVpo4MnDdhggDpTYsJ9hxGH/vXTEhEEZIKZTk9e6cQTRle/Ncq
NRQ8kvLO2mkuUj5RRjercpRcFMfagniF8H3ynyN+wCp50od4DygR/1lOROmrjFHgLL8uhjt0d580
2XaGMMx0nFz/IxF1PQ58iCcmG9TXlSqZH5ZxKwflMfJOIN2i7eHTdFyB7FNP61MrvtjkSUg+Y0eZ
ro0uzXHarP/+lSr/rZ/pHsJSZ2flGOVbRjq2ZqUpEuhijvXWsBz4xuksHWPH3Of9o327N09GWeU6
Lc1tvRDbS28gUdkniub+hAmROUVlItd/Zc+YP7RgcGPP6q5JdDBu4ZHiix2RedIFGdlTTMNgdrf1
RjtZJ2fEUm/z0jxtprKrzg97qhBFEfpgogBGwOD26H2HC9+rd73Uo1QhKhEQAiMOqJC4asSdLhMF
A6InkpoglVzRNEMzGx2paxxsPM7ETdZ3fCFeSIPHhaZqYswAvGhBHZdyzmVG68QpDWK1mZtIquRa
92r13y4YZ2qNthdTzf7JC6XO2v0Ym3l31OS5TFHelayCZiLFWGWWR7YPdt5/WHZH/+rPn+lcddDW
4UtBxkNUbmKOsCS7H9cbROgTAsMNhAB28kouT59YClTrjrLhpGtXUvEmQX3NyGfCUDiIH2aEJhqC
5qYb6Nls79YaVqyy4W5wv5heuMMJKfSUtKhHwaE/Z4NZlAy2SyjX07Srn7acCcbNH9/iWpIpjoEL
kWMxxBrrXHCHzW7JWRvv8KjbMcM51ACQBSZ0pgYxba7zWMKUPc9/lMJtEiuLKHHJ+Bzi53yaS9/V
t8AA/EpvxEn+kd18+AhUNWgITjRrRRtdglPHB2zb4xpC8zP+uwrC1KdBN7YyfrgRoHKtl3QC8FE/
V08gO9n//y9CLM3KBs/GDiu+yiOe7GFAGP9RTX6hyzh9lgg58ZSvgkXSwDbbNo/dUJo9z2WovAV2
p+0l6awb33/c6vkUdHzijUWtdyl4MT8aMA4UgG7d239H/jAQEMl6yPsIpPBPY+DGE0iJR1RFqWA2
D8+FJJuNXcW7lqFGhYUpf9GEQYHIZelQIdAI3uYjkZ97AqaaFqoFZ/pnh3lnjbYzxr0vZijxMeRU
SKbQnCbki3TJm9+o3fOpNFLANabRsudRc6Vg4AcGT1DCB5o+rgTh1r6NETo7+tYMc139QYlypcGk
1VUe9ndzH7+lfI80TeGTKGB7pbSFaoHluRSSGPanm8DW+RJn5dvGG1sWRPCv2/aGvduJJlZ2QZPd
YI+YdSJEZlOOCVyipxAPOmaBffngJYDLjRHwIA4/fTSLFu9Fa9ET2nRbDERa006KgGaKdlRVoJTe
wSMxiTmpVqlnw6RjhQPKGzyJ6rQ62iRFzh7T7e6nPAGTPzDQFyGCFwbocq9VaGGawedTd34ZBhLE
ZUSpQhNwoidw89GNx0AFpynrkiW1jn8me9raW3n42RtcrNd47YEda3BCEsislR3uJ9+qLov+JCY/
TGeQCucm9V7u6sk9WtBJpiUxMBHWriCeFEg+BiG36R9/8zL4/iDsdjQjRNRfEZgGSMQO6YBYfnH/
NGD1grt0XYLJnTbyCiJd/FsAQmiq8urwOQHBHnpZkJXvMZQwzuYIBMxKGAMsWDVGjHIsH9S2arQ1
w27FFGMKQSGZWcjIoTzwltCjB/L1eMDBd8eGuDzfvWE3jqh3ZTJ77AABKCTW6gUMNDdnJBcqSdS2
971S7+uNn7H6EPvHlnJuNAIs3UtV5c7dF6nd2IKQTun7hlhTvbXt3FcwxrP04sJ2Ppd9SO5QlnEG
Zt/x8wlPDYXcwgL/bfi57GbXAQEAgkIG1RHDbNNSWZOH9m+5w/cfFzKn5xURvt8oyujFZ110C4u6
EMAGkb9QDLVls9k04F0iqU54SaeXM7Z/N+n8GxO7mhphKOMtuE10xmdcgdPfw4EH+fPuAE6opF1w
zvuK0rg3ued/Q/h3od3L1O8hb6U5H631raY17IcQwlnu+El1sWM0207flS362T+McBrDwsn+VpOp
+RxM0VDhaC1JzwClcEr6VS7ShagMxrM4owmbrOWqiUX5ZGuyyKQ7QxMoq/IPkcku1q8xP9Entjxq
QEPQ8l7c5zjVUgYQgd9IIMX4LN732OHSd2VXkuF1u2+vdlzAvx/KEYvsRdfxIPAobAeP0HbJWXpz
It2xiEXay3yv8Qnk4ojSYKJgRdqSp7+OKSCHzL7T2wq4jqsC6WqserGWXfm/pzTjAGpyrMfxyUbe
09l4+ojRb95WcFlewFXHYs32JPCyMU6AoB+LXfiMpmp36NQSwHcWqUPbbO2PlSLFIrljteeM2Bms
1Ida/6HQjYQ+48j+DIP+T9yqP3/0G8LATbtlimjUTBTBYLI39RnOojP112zcE6dJ7xCmNiManNzk
eW/wlJLdXkO+lhtG5pfkiEpwjg3qxKMlED+SIm2MykfFLs7AC972DjrV0xoBIUeTyRzRMJKojV0B
+D3sM3UW5XNA+FiLOpuDkaZGsp01WtdCtFK5uX8Tspiw9cgYN7DGfpH8odu1eiINpmdvyxYXFekg
XxZYwKZEoKuNVjtv6DuN70T16IJD7ea8tkrJHBkDw/Rv62hM4kkMbYuqisRC/x0mPufs5+gLv9yY
QjhglrYmjP7C7YgUcyGK4+efIIf1I31LKNnhOT+x/4Gt6xYZnYMememcBwN7TZ29CKJ2/0sa7dRe
XcXJqAKVDMcbZYdjGI0KsvOxfgkw3tX7CpJDUBM/P/fLEkmatKmOc/AZ9sDDdcBiUWw8BhD9Qf3s
x0dml9sPxnmyhuC7Xhtouvy0lFNAojsTQ14zwwSCGI5m/jqeGN9o05kai8xhTefD86eDzBghkUON
dPN5hDtzIKNzV+hNFsq9J6Zirlvr5+NSTlF9RWJHBM8INtwglp20PN5E+NM1Gk1UfMB4K0PNF7gz
ujhtccmaJBc+ZDlQrX3YOalOxwnqWPgG58ExrcfmElBJIKcTuVRIiurpb3mIjFT8wjCiVUyzTXOf
C5PEx1kTBhnTuwTQttL3D0Ax8+yS4SR3PvB0uQrx4lep44IB2SUfSjgd8FtFgPW3UUrO0ezQN5Xz
zIWSBC0YI1VBhzDKyvi0ScGpZ2CrP9Uk1pXfeECqrKxr9O4HWPr3KWhh7tiSbikTeR86/NsKPjTL
17ibhRCwWLqWz2ysnU3MWZcIcnS8qGXxwVrk6Ke/iBW/TLHeaJbblF6s6X0YxNFlMFwjTwg1zLir
cgQuYMtzodAb2AZeAfpV4HlDK62dXvIe6QvPRZWxYM5MbKFpPKzC43vFrcEnO5awTFgxR5Fpg6pP
SrjC+kIo953bbDJQceLUMjXnSUJ8KUez0+woafC1Q0u+HOfCFh5m/ELXrX7ORJqk8Jc2mEmDFQhJ
AMKZra2768kgUDpQM3JKy9pLHNOP2X/gzvbqCR9kEDFdFUmNChUPUePxWqPryxgT2EI8TJZ2HXn9
jRwJRsYLEJduOJYcwgV/VcHaDhgV7pKPi4KnKPD0m7ODk4rzFP7PzP/hlkeo23fHliLtLeElJkNQ
B+O581/evAArujF0pwrDagMbdnLc28PYeVwhbzTtzzIUKStidNO9F/xaes1rhuYIBcH43pPl746P
D0rnRxgytUqIyQ4gkKL9fbWbIPyzB9LJgZajWzNs1rS7Ty9jq1pCiQYC7LLIfNdnG25xow2EmebD
kbey/G+asHD9mw71OwkgGKj5oIGCZ4EXyU9N3hQOE2iYcnD/yVwsEeuuCNvBhIB1SNN8sWPQThVb
lr0q0L8xhWdYHfQefp/fcwNCZmoIphC1KNsMSY4PoRJNuR/oivflbPnwTZsSCnLo7jP6SWf6Nf+u
mPX3NsQNnZJ/ix3E1pWBv7BYZVeZpuAT8t5M5haYAxZ6gf2Uo0kHbK5IgYSsxcuihF+zEobWf23e
OOPo2ZWi/eBKPZxejRBqrqujQiBoor2E+BIq82JgTWjx8TXSRQGnvgvLx3JIGptE4E8VScEKrmou
ra5dxENtFniBhfVS2CleZMV2ZhWSCRKHQWIwJ7JRncWthGiD8MGnjY+Mk0oV8ikdbxb89DjNQZby
bs3e7KQP6QC3GgcgxAtn6LhYrfHM63tKO0nCTuv8NJXDj+tDBSdRMk+GEJGhmXnXxJepvQS+gJlv
9CoJfvm1YGid4WQycSJhT+dz9l6O2zxkiFZsLvAWg0pIiiTDxDUC24ylj9BQWvPItDLaQVcxRGV5
F/qDNkAC8y9SjXGUjx2jPATyvN0t0EXmpHtadnRJp2ZtTHVamFTuGtJFUDszLtOG3TL0pUQiQE0s
3XruvcyL7lgqWk3CUCwPwaxpmStMG5m1rObooffprnUUdboMTBarYoKp3FI4XktbI2+MSjLMD7Ck
kmNpISBuSCzaLa5FNOTHhzdJwkzj2itB/zLiGcpLfpI57xmXGQ8oihIXyYPvKxoR38+WdmRg1WM5
atHxS7DuPDGpdUzqjcrm46PRtec6BY6RbPTB5iQSGA9Kgo75fq5iJfTVTwcnltV+U9yySjOCHW1t
CH+JsHQs6EEdzNSKEsWZeEfNQWJ0Lm386G1L+9fdF3fWcR6Vxx+aWw9+TyKOOj8GE8JJnnbE+XKY
wq6sMFIuHAIraSl3aHk2bvDIC+OD4fJg6nFGMct9Fhz1LQJibYB8B5KZhwqSSGtUXNp76RGmoa81
jhdgTKiUQ9IITSYlwjyTZXKjt4a9ySiCF+TFAMzMxRl3ae9du8iYqUBulAlCPMvmwz/5LAlgBUCO
sz8waZ3JXZBBmWBY5msc5YitZhUMXV4kiegVuyE/UseJmF0NX7LsXizyfZryPR/229C4btF75DJm
5lIcJ9acSTPegD76MtMGZ9gcc9iwH2j6wSl/vfAwI9G2SfBArvcBA1PnGr8hlPDhgZXYt0x75i1l
6OL3XXA5k4bVWVN5jJn0iKa+eRB/yIxI/kAJCP0hQc2uzXGVNP+4MBeBtVzSIjasg4dViz/8LLj9
Upd2zJfIv3AeJ4BDLkh3UfNvz7CQ3Bv2441uHeCc2IiEYDn658LCbhO2IFcViWg0NRFRrizhVuUi
9eoUSWU0MmkLWj0u2CtJSiqipZr+wlDBBEyLKXi4g8e5yG5hH8KeW0Uh2Ga2PE47EFMcue2Db6QB
GINen+x6MbGi4mwPAFY0fc+rjJgW5A86Xhp5nMKI6GDqQEEupMZYkV89qOPNSPh9Rv++L8wFUBN/
OZaStaO9j99Ri+6I3IhErZk4zl++HEMCnrVIBfKUFeeQN99vnMneVhg1BwhctwyVjHovjsmJla/w
F1zlriiLH6OU0e82Yk1ooTzFnL9YSMr3H9J7tXU+Zkv5cmpF3z4MF8p/Un3LdhQyWly0QE2PH84o
rEfB0OAPQTTfdP1pW5jAoKrDnAJbU0nzlKl2Fys2StCSUNYLj/38/jH/VbDOn9Jf4/Z0SpTeRBCi
kYsxJVHhcjc7cUjRXLOibeCBLKt3CnWy9rPc2P0aT+9rdQYBJAcIU/mqu5jf2L/obyLoBWPjFBGZ
s5Y755hwjWFeyHADMHDFaaueQWHHmBvqJMSczQP43jN06zNN25mgGio81bZlotsqI2WU1tseu47Z
kbTIqLWkfU+MNh1Vc8pARgYr/5LaCoWgcv5/g6u4dZac/oGE39/qvz5yI9z/ttLYZ+7V2QphP5tj
WNN/mIZ9Tdfu08KVLLhWGK4FlURUY2ceflIWSxo5jwUAncrtSsmg400FKXUUNIHlJtICP4fTVpHn
7oHFQOHIUn8cN8b7qEL/kG3OebDz3gXq8GMMHtw1AdFZB/f5KfFTsaPfLiD47Ln7jn7lTEYlpeZG
HqQwzJ9zX60ZAH1+FWpT1xsozG/moS1eeIeVQWDII4UVTwagVU3P6e39Uuz072iVy3F66XADW0XA
w5gC2QHKEexr9HXsnP5PGYf0C4WzMmw7UFNQa7C44W+D7Z81cfebrovD6qKnor/ZIYKIP7Z3Daea
M+KJVpdFGxk2dYjvHJnQs6stNefaSQzzr7bKtdN0j6YebS1zgKD/jY8oqMWjZO18aWzSD4/BqNN9
kSqaGu9oiy0Jwa65Rdk60hqpTKMjmHpKWayKhuqw41sACKdxcIdfqf1/IczaxzDUW6/qLKhe/vVw
kSfqldafwYVrS2hD/oQnxsTdNahDH58dU9t6qPIHl51Yq4Fw+DFGmzULWUB+BEjWvzg94BFq+1Hs
N61RXs8WIMFOHRhtXDHVUbl3Numib0VRjCWed0Rlbtrs7WPvWlg2Jx3NM6TnIxPPciOhiSHa9vPb
1VfIo32XSEl10QtaJOl91In12Q3Y9uwtbkX88xpfweSzDs5qiP3Cvtt2bODXs6t9sl5J3mj07L6u
1nUafZRyk8Q5dDEuNkYTpYwcAyNdGze08eZxAAnUUCgGVLBv1MNpHXudOcIzgz7KMozTyZ9jKyvG
DgIJjRwOnf2UNmeYkpRvL9zo33o+awOQ2vn3GMANy1vrHYvOnNVF+yz/rC4EogTqxrmjc6x3qP/N
umrmKYB6nQrcxzY935bCRUcg/EjYLQ9hp66WOGuA9VMIcMhcIc2F63YOMftB8up+AbbIItq5kmM4
vQ6aGsz8L9UM4f6hFMu9ZX0EA2ekAWUZlN5ZRRfilyVZ3NtgYFG453zaodJvAcwAsbsR3cSvA6sX
CUDRNPkjbsHvIrevnz8frjrFa7Va5VGV+rqNSDtE7AXo3uF2Nf44zlKaanywd0QG/1LfiPKOtn4e
57Oe4jL5W0MS6vX5rVjfA5AFipriYjlUPetehRI6necED9iHRNz2CdVwdLtffaRcbddJVIGauyzF
q3P69C2onBnFbluKsBPniDSoN9jzwUxGn0UesIsFhn2GQ0+mjarUZMecf/+nQrnmOpMz/+4KTvp5
+HvAa8KbJnC4eEyf283dyTxqmhulzd8UTud32KNoI+Eduevpb9Og9j7knQ+ycV4fK4iyUndRlk7S
mRMcyGsjmOeI92iKlD5gVxFRVcTiOpX4/OJqsr28hwNJPWrBRYWUYdCXNdwl8zQsdJ2XHSaqUgpq
HJ1BniaMm775Spgs1OmkIkqS79eh2tV3qfOABZCfmjRazm9KCYkZaWTQn7kbiVf5jee4dh7Ghn9T
vxU/u4bg14Pv+DI7QzyjjlogKkQdg9eI4VKUggjRY9KhhQd7FtZI1ZRXv9DFc0qdJa19qwYb4mno
97Mczr9dd7KLRvZ3pZg3rTq9mR+8gb0UJaMR0O/ATy8yZlgWlD16Wl85qP762H55mjnajn/O2WFP
PQ/CsKxEWc8zXWUDzFeIPqL9F9Ca+ZxR4SZcU3N5hahJFHu+M4l3RKni99npaPe0CBBQPt+/OfED
3tIPfbzqE+kmx5FoxwAlJvbejTgJxYV8brvAq/WmaIVVXqQSZlYsLEPp7JIcFfYJinyuCgDkgRxZ
dYKI//Z+4UpZJ56T/Gp1CczjT1s67gPr8jF2GGhrD/6+jEOuNQr5FPvxRoLApl8STCcL2HZiq8Je
y6k92y9gCmMGxxtN0kfany3DycabJT/4xAZKNevk6/hj47vjLFgRlWT8qU27MP0SugZP9ts3hPQC
bj5EowUDrdFHzligz47gvXMTy3C/V6mlUQ9VyABJIS6pU7abl+KaZKTrJD02mt0GjEXr4Se8ECfI
VloeLelHylGGct9AJmDIwpn9cwM9TaO03L0e1P8IFGHoxmVFy7efq5fR1iJ034m0PrlIaCpsXTEO
wpflFcw9ai7ND+/kEQonGqXhXHvz2AwmpuMzWmoFLExTE8hWILZGCy0zJ8M9a2rICnUqm+YV+JI3
Y89VSvtvR2uIQYE+4ayKH/P9A7cT9YuSN7RcLD2ORuann3tw7F+dtcL7g5JfhvHkFpKNp6zhCj6y
3/qch8lJsJ7JhAO4M3wcGP91U0ZJUttPfTmiiA9+a6sXLCVqd1lsZn0x56kicMB6Mzk1iQiBr3ph
3vg2G/SzRcQgMRTcc0NjSy6bLxsKBsGKsfDm+bHExWK5vJg60BZxRIdEuxMhWGuRiJjaXdinyqsa
8+hfSyF6BatIlNT6LsIAp1OJiryPyFjwhEbRhSx4uV06CBHPWgc75jMP5KqLIynOWy+N01rjUQJq
gJBNxl6Gw4q9HO9Lx2bX55PWmmTR6CX0qts9j3HvP3fDAy0LALYzE204gEsjSJ4S6GWss8xuc712
M2gGz3zPTkuKm8C02pXL9AsV9ktqCgh4F9xN/qz++gzYLVNZjV4GfAn35ekJ3Cp2+GZo12ufgF0Q
Cn+a2BEVBK9wJHBpIwkMJ6EawZLPOarAFoSdeRu1BlukWGBHcwDKnnTwKmR7ltgiKRK3DYmTV1L7
LcLzVCFhfaaH/6Cz6zAzwMqyGQ+NSpA7I7OwSaQHs/6yeq8KZTlbhtmMJm2gEtLPrYpmZ+++ySSu
eO6WUQqd5BV24STuX33c9sHGaOpOwnijWx732y7amLiVviJp+QPgUSH5MYkASBus2QinTOUl/4Nx
IeaV6/h10k36Kt4wR0LNnx4mZnzkiJB+DZJLKGv/juORKKDzbc6kxrPZyECZuW3fA/VBfWUcICei
RZE+niZHnAhlzsMiumHNv0ss1u8tWnxri+ohsmO197QHIDe8j2kMKDi3Z0IJwxSoFbUmtqhXrFNr
ZtqRdOuvHRZ4bXxPd/kbnOId6vj9pc8teCVSV2Jo5rketL6FrjPxi/4RrWTGP4xNoKJIuH4RNCD3
odgjH5N0XAmPA3AsU/K5Sc6RfROxKL/6+3bEV6tHECDg/Ouwn4DvRkeI2Rwt7czCWCWHLK5D4WrQ
sIb5VNR56dbc/Z9cVIlGxH0+IITBCtSRmBXD88bIZgmFPRtWq3kn/0KJRsvng6PnpCMx/70uR8Ev
8WvaKxN0qUJS9yIKfccFpncoiga01FIAt994LGkgHfCEIdJCFUX1VpYrKUj/AdEKYYRSz8Uo30n3
5P7QVFv+muQUny/NTlqr7cL2sleILsGoHZ5CH43WQDo75xWurK1VQv09EpsflIbuqG3Fvl5kFGHA
BaAJJrWVLvqYWoTWEy1QotK1CTTluCGrPoGaAynBct8Gv8A0tamYSQzQEOedUTBiTLLft8c3/4IG
/HC8Lp9UOmODYf6z/AG7wlRUHjiiAUObKDGFG1p85QqDQPW+vvyqtWut26h1LUhgX1GJYiVzhfqp
Pz6/8iZRtVShkmEVKdrBnN93/44J7ZNRo6Az2eIK4NI5VaKWsDza0kbKCmCa2xvnFga6edx6rZSr
NEo4xDU6cQ/D2pQK2nB0OybvYsYfxc+iV2YrfOArDtn0eup4jJquFri0y4LJ8UWb4+JzsTGxYYew
tRJkxX1n+svDhSXiMyrSSXQmjnJfNLXJsZHY5kX621Ed/iFWzSEuTCcadO+hxSDFbko9tzjDgZZE
EcCcP/KL16t2e2wu2+h2om02pMQR8ikMayoAo2ooVT1+n1rnCEfgj+nwFxmXu5SLnqSj+psHaOM1
GWAJGdJHNVZGmba2DiA0KGRZbKOygsFmrkkZI7aA3GE+g9MplLPUnbaKrrfLPnaZ5cwWFjXWbcVj
qytFX5tbBFivUnKq+LoNlYMw8U3lJ2LpxVTl0T2cvUXK7pV90JUDWpKVz9fo6f29YmxWG4oMlMPb
fAzRH3bouMNwjZ+odV5Hk2YKOc8hCZCbCLulav85pVf6/qrxNw2Src5V6wcfIBKGGz0V9OjZV9Rc
imGcKPtWa369ldGF9mlrKkskaVVaxiTUafCUW2cSQcvOv+6DLERvwnR6vtnapKBBdpCePoL+ISwn
OX7gTueqdf1L2KusT+tIEYr7bfb0glF5S8r1wSU4ytEqDq47QJbpQmvi0AGwMDyMOUOb92yefefZ
2ZcrnYW5RxUTFp4T0/4i9hxQfd/GlHIKOPE+04KIIcwPTRYO6uSxfr1Qk5dnkeug/4RIwR0WuxRy
oVQb16wJNgooEUG+CY5J6j8PemgI8fqVZyqPczs0almG2vokN/q3tLDS437ShjIwJIv+XFq88s1s
aCyckXa6WG2D4HgR+rlSMdBRCkCpzXqDMjTrjwWvBMKerdiZ6GUoXtZYfKdxPpwa5wnGl6Ee7dB8
lSyjy3laxut+sQF6G3BlkgPgcGUCn+4x0cLrt/NnZE56tNONzSjkVvhvmKc4RXxX5YQL/+PlskAk
Ci5Spzayt1/z2MFiLZ+zhMknxmITzFlfMU4xbQ0o+P/g9jMDFIOKVgRnUu1HtGZhihKtgX9+8F9r
hFZBBtxsn1bGcPJXc0TNXePJw5gmWkYZfWfTUsikIzX02YWW5geEyH8UJVZxHtyHwfg8lB0+MWOc
Y3kHOQ3LoCzhCWoj8QO8uV5uCvdwwEiAWmX7ClpMiDU/oA4bRXYi2hE/Q73T39B31WeeyXJqmDS5
kZnqQIebAldCsH7aQzchDoe5m01+SFGuPa4cQQ9ToQ1MQF3BsXYK553q4PKOdLsWMi6lJN4+GOdR
ktm1b/1ENobuYN/Mk1WtLCVXiKV/BErn/02QGeuGvDe7IsriucO+BTkYofVf/hyaJAfk4H8EplC+
4w4Ytl/87v4euiR+Nfv88DGtYpI3/5wYbt2nkXcK9UzoPRGcsX3YujTnzbmDfxFfJn2J+A8GfHPx
ukZuAdTfG9zINND5RxOWz7AlCtbSUjRyYXFFhoR0eTDb09MmwT2UXV9+33+zF3oCRS1dkv7o1V4L
0leojR6WHmd6uMjEYLVYth0TosvXyrx7+FyZri/A7zxucOjOXGZp1OQucGd+/P6dp86VxzhpbggS
xp0aApWFDcCvGSBAwrMcNPaMVXv1SVDvkd/dN94/UOOcWW+C8glFQmkeqfw6B9G3QC9MGO7rItYj
MSnC2WnX23YJdyynTAOWILN5qWwxWYFHZ7GkEtbAJorewz/8EqOZBEcpBN8+ozWU3XkcOmih8v8o
duqAutYeUIgHdGgv2aOlC+HhZ6DUIbfy/YDdRYANprTAKhpqn6GccPcgAVs1/Ff/O5wXtLMowYZ7
iX/TONzKUD8H3KuvtLzxRwZax1lkiZ8+C9mnwPtbUypDQNeCeteYJ6UqGwMnLcfO+MBW59N3oC87
k5lGrHv7EkCyILIrnWiFdqJ+WZ1JkIWajb+KbTuRshYdt+UBpRq00qmhyKOYapjq0VgbJNkiKYSR
5gG9O8ISASymHQc4auLkwMfXsu0A1VMBF/TXtP0ODf8MFhOD+fhIsQgxi9W3SPC1vAUZ6O6JMueJ
pbNYNbcu2UtPdXnlGJhUPTihzK1FId1oj/jzUoXlXbj2WBYG+nPGcJpsWV0kNhVPkpbwMx8eWwU1
4IBN9MPgseeBqt4+WRMVcbYTyPzoLa/YEBbsSMMC+YWGqNJzAsz9HFg088VmAuiKtJgO6A57aT+S
YduNE8vt78K416QDhizHjV4OL0pOuiEFcBMfKTBVvJgpAs1iXrctxYmsPUygIxZRwEx7uC4g0LsL
hKM4Nk9tyBaY2QmHvrp+aBUMSn0cAELu7CiKVHOI1p3+F46f8V9aau8vGO20RPKuA+PtfS2kKu8a
t1q3cILwufVe3+3P50VqoOzGEM42RDyY2TZWaX7/Zb5kTACK0Z2I9oJZSSxSYDEtAZO3rSbkxobk
MwkVCPHCSH3l8E6h1QXDf2Q7MZtlj70wJv/9yub6+qfcrH4eXmblEG98BIjEg+pKI/MYU3w8n8bz
oRGhkwxdKc/Sj77G16b28y2tcZhPpGOZ4Teb4KVQ9Nka2osknz5ANNAwn6UA1ujbHyTKQxE4elrt
au5A027g77VkzrNSxYHwjrErSg8cjG0Bx2lrSjr6yN7h2tjVFOjwyI5AOyKeZ2fByx6OyTe0PchX
2ypgkT8c/GqgRpUkJWvzA/3I0KOoXkc3yq8oaWdUnAUIp7Z8v/OpZNxlq7hkFTYOGvT9vHgbycQC
HiYPXKezVq62ChL5TXkwt88ABcoPkXgEB2zVajgyxq5ooZc9/Ivlb7rxJzDuw/4ZeOkcOo7oMObm
+J8D6YhdJ93rAYKmf0T04Pfwd9renVOFXlFUwp0Ow7TATN0EwPi5e2DfoZwcJtCL0GeBgN2nWh6M
303rQJfm1kmRWagl/I/3gFOzVIYccVAvkS4eyXVrFuiVYyYyI3uIHC3Ku7s3CrwlyoshyPkS+Cbh
ToNfqzidHj421DsFN8twd68uwkkI2iYzimSrHES9uLIz/DDx0ExDl4AvIjpx7KggAzcwXzA96V9x
rtezDpm4Q284xB0lxsE/SqDOUoPWooi1kjLRl6OmydOabwKzLUdin1O3H93ArKipbibUquqa8e8z
gdlnFSMqxTKfzXIT2xLQvQ7mCAGfr5ey5ZzX60k8TaCakMOtgxZlAHN/b/lt5Cd9RtRmEFFwvd0p
uhrmEDwxo5ZirevCuuaVWhFek8LM3eNSVJ4FKMlLVJfMrI4HOLo7NhwTpFKWdh8XlCLx+E9lFLd8
Ua9np+qPa+VfkJ7ecCqtRiIf5iTnRftG4aqBRwZd0AHwa9oLb3pkp/HSskhKhgBULzlgOS7mAcbp
hcvP3YwDj8d2xQiVJO27dxkqJ64+YPO2czwot62Or3U6+AtN9qBy/txf8MATFl2vXv09mVEa7W0v
9B+fA/1qMCaSvx3Kc/gBDLgrdeK+GZU8JQN/RMkUI4pyoBf+c/mb0UXlvfKWgbb0m97C+Q52Uwln
h9kKVvB8Jt0eUXi6anUOoBj+TRm/fwj/r48HCrCdW/9p/++ep3ddmSHkhajnN3RuOiZhgJFvXflj
6P6vmVc31/9oCSePEVupFNxpMr5BJfouKtcdjHtNRl1O3gXIVIjfG6+7OeNQHUyAeWqbmbAoSri/
b/ZTwyM4DuYM+UkGmHOJMMYK8kzwlbsfobNJ9xvK9sY7NNVm4v7zW7Lu37zuLtyBYx21Qa777WgX
QGlpl2PnWix9gPhE89JCHhIaA8mrJuNm+02q3MZ4HRbMmRRj8wunC9gGyVplYPsFAQ8JzlsnkOVA
GgS+hxuXLi4jUlJV23ncEz3ObG1g1LXWLjv2lx2h1KrSYFW5gi3J98UFL95SAORDaNsO/P1YWanv
L0fOYuTJejIwQ3fh6yaqq3LpLfpoOxIhh8mINHubKpcQVwFjVot5Gwmec7XkNdXxoM2cMnXZ6/TY
yslGA03ppUTPibB7GtHX7xHH96O5XyGXlnAzURkBtsvsjf76aDJlv4h1x00pE6bI7R4/BzrdAr9X
XCzAM+9nWWU4f3NDKdY9asHCOmIYSLMql6QhhTuAX+EEUGdzwp3wdMBOW6vjwI0y2r05ui/d5M2P
+m+9rd4SE1j1T2wswjLNDXFHP/XmMPqaeXEcH9R5V7mJPo/06y8dj4lCbfG3S+1UdawjwRwx1KyJ
4DibHEJpi2FjwLUqWhQo/L50DqjhFwxbphYAUkX6xntaWRmJQAHf2Je8lefQ83d4fofPUnTrdc5R
/WNpnFb65TLDCj/Xo42jQvcu81LXxIg9R6NeLx4+7LNREwZ7w/ko6/c+oSipbkZLTOuvkSk34eJz
loEENeZpZxyFagF4EfxYR5K1uoXw2H0zRWbRltLJvpitHG70oAUDSxEfYK1QLAW+4nvUsjVqIpQl
m5TWODNY9+HRzcOe780TEQcakoWuB5uVekswJsoGrDUdLpn8m/0nzwI5bFrJuUc56SFOypcHGe8u
jIjFIHX33f9ylewvje+DAF3/hqEK0Dffa2a4gGz4Sy3KpJw3nVmOY7JHrYzX0zAZdLrrqDcQXfMg
UTGL4dYGahT+F24T2E8bHORTfWYVFXv4ZMX3KDD5JPfLHl5V7I0xufDwffdKlGbkcMIpuUahTDLo
JZSnjEzc0OdLlXNnbdv4wdoSwCkyTzUGDQ9fDDmmL5bZqTYrCJLdNfOZyEj3+fc7cCt5ehoU5hSY
t9GOzLIcxTzggWmlTiz8NLp5QBlXlZIRipFzvVtSJ8g7Yvm34OGHzte9VxYfhO0pleng5Y8FeTPU
77obXa/13Tm8SSLZT46nCGTgUaBPq0o5/8WMw3Lg9T1eQ8gAJShcpdNIiwm/HsPlPSGIMCG/bnOw
cQKSGe0lg1aWFcX0NXd9RRmvLdFn7ef3u8yCbNMOKj1ZxVnJAyAqi1OoCtV4/NNbKNWsuowv6Zyl
FRUu2lfH+e3PfuPBPXXCLSZUm/p3voq85BQZdZpa9b9+uYkLt1dgnv4T9t3DcOcdTLM6gNfJlKZa
6Y39I5ToF8fKCgRLn7z5s8EFeVlgzoajim7RVoAmAA6MASjdGKb+aKXMPgxRsatjqFmavKMs500s
KzyAY/Q9OQUqWjmRzjksKXBrSLAMlMv3vy1Ky3Q1BLSm/k8Qb/nKu3H9rRb3DIsgNt3R7LHbedYb
DWXx3V7c9mDK1QPJkklE9Z7VWXaT6ora4ePyRHi2iyQu3moPO4t3yP3x7gJMA2M+mBD15ET1Y/yT
khdwcdoampwtd+Sl7m7XzJZZKA90k6tojCaAdTWmR/UAiXl5PKUxbVWTpHgAvtY6E5FeKCx6kT1V
OSa/eTXLeP1dWWIFx7rE0TZszZroiTJEYSU1HQ3gFDu0CX0Q3QoJ4FG76NEFIi5gdvyH8iPLEFH8
aIjtWK4DBsPMjbSu1X7x0IYZScENXW2JX0MW4NIE23SDOmRhT/hM36FCy4yIoZMV5CosvT9PcGH7
t4Hy51HjJKlha+yJdnn0y/cwIu9bdDWQAF5tNVL5iQcA7LZ88V5U2Mf/5SWl+kjAYDO5b+/MGhAw
/LXMT/HdGNolSDnD5leXcmmNScz1DCB8A/aJT78lHa1fQsoWhcuZWp97D9OVU0abNmJNKm0rYUIa
ZX79cIHUv4r1A5v/QhhgtPjlGjvfwQaptC0iWlhjutQF8IoIuoyBQW/KfJwnTwDWojzNBtnF915h
sEJNnsyc5hHh2rdOm2totxVyWCq+5zg3lEcH97eNfKcrln6dIDMLrqtGPej0u/Z4RLAcanJse8cw
ZGPOYteyhSSm3LCFAadxuoI8xi9EJel1xn0Zd0TlbaasHEa4GDbBHM+mXpJaW3DC+xIMlhueAZdo
lFg9LvVpxKkMWa2yW+wdFDImLMSogfHzowqjsg4SQ9GOw0fRzckLDzGR5/G2Ae/85co50QTsP5vG
JZliSTdpM7RfddCFSuF0aZz3+/+3Ygp9GQ1L91ULBId1h394I68L/MsfZqZPWwQXJy+UI+hufPpE
S54Mc9Z1MHpLQQU0sdIwhvSwnZo6AOggpGFcDflIw0Z2M7BYvVyILZt3qeFY/7yUpvc2fifXVr/I
4jtTg87wFywcuL3o4vJBspZsTq6AaEOTlZAIXlAnyjTFBYmooT0T+GehV7VkAWUx/9NQI2QMdoSx
C7Pdy3Q1MlfopHcP89jCw2owKWdH9543P8hIjsy0k4qLQIPwRHFMPrZPRYyTN5J32xSK1aotXJZO
609i3beFu5x1un+e1PjDuwQh5CzZB0WoQPOLcg8Kuh4qM9ZTWD0WNRzIwjhSmvlN8F3Y/lwKWn3q
KrKE+dHIo3cI0+eVZ6JYjWcLMiwpjRUpsuJW650b1Hlt5rzpeZ3DkOp5BTzDOJO70knOfzzYSkZY
VI9wpe+m/iFPePBsxO6dOzVQh5bvLUzC6aIp+uCxKYM3ZHj7ExM2QdcHqz8Z3kf9fR7mN4zBNnit
m0VumUXtTYhel2AFjUmBLo4gI4AH+9x4ao3f7xMeWiFtBvrudcsLYe450loj+5Q/k7+7Sl7AYDaP
aF6/XQpXeZJNNXJGFD+cyB9yAvhl8A/KePHYW5v4n5w+5ZC+2axRfEmwK6ztJEo56pHun9KqKrix
4s0txC3NVL+K/kSd0SuF/fpFlOxa40x8CkgcDlHjReTd+P5YFTkwXb+0Q1/Ka8JJfs/B5HE6METC
R6D7IcIH0r9raal0Uw1IMpxnjTYEZT8iU50iBWXd20w42TGYe3tsHjJHNCOdvKssMRilszEy1Q34
hkk8gWUzyGjerux3RXy5z4ZuRyPZcP+R1LAglftvBN5smkHUTZaq3zXcDg4x1S7ClKDLltvavVjA
GmcpXJVFk1s+9hSstYGj3KtIENUJXivJnr65AqA2DA919X3gAZD5AWgt6q51r5AgtvZ8QOSXhdDB
6KfdGFNa5SgsdPfPCwTCuIX3raf4i2NCZp71cmPwZ8/5cVEVW3hsBzbLzhhYEx2iYURrstqIsvzI
sVzXUro3HckF9eU6G648a9gfaAOHUfbQQrQiIZOdFto8nsJa/liLToMnDyca6Mu8zKp5hscIAxDh
0xAaVGoQ1Nk7WObDEg8foSUwKeVU+uuMPwLmvAodye8Ykj5ND0VAK/Ug0ux+o3XiEaIhH1rW4M3o
2NEwkPEt3taarQFvZcon+RBhiaDBVXnG8jx2TLBgmJ6wr+WQxkoD872Myw3lPcCGTtIId7C+ocqw
CZmzIlitRFsXCQmmRKEXiQaHnl+vizBuL3NKvxi2U9PBnwXx4ocl8Wf5/ZmEvTd7w+Mu1uhv2UV+
pLqIG+KRh8j+1/YaqI93dKFbOSW7A/E+b6KeRrE+YUcFouXGAzgN+7JfJo5x+wuPKo7erCX0bfTA
OTxKlscHHz1ZB8Zx4palWrjMvvl1kqiVwcLVwe8VlihxsRDCb/mb7v1U/T6wh8kQyF0/BIvfrTfm
/qIW8nBdCueZOIIMiFmAmB2pZ41C+kCuaJfnVFaJiXMxtqnrHspBSWHqubzYYG0AAxTzz0gGc1xR
6La7G2Sbfu6nfqLJpVJxoU+HLFmIUPgKKcl/xnnv3Im/dVMKINS1nI9AbDMBphW5S6vvMDYdvRU5
k3896R4y8jTRGjIBHipNKvaI3HLfH/eiSxv6yajeU5wIFSLdR0bhpJlTJ6lPYxF3CnAtWv9mAiUX
4JmzyvD/Aa8bUCfvxDNXWwrDcewJqX6fvyzSF6KgYEzD9E+RYywgcWKcqEhJ0BxLV6c61jbY0L95
xgyYZ/HWW3BSBE3Cj03wBduSLSA/ioiyn16tC8ePbN+DEdQMoM3CnBsWFPYUIJn5SNfKwubyu6u0
fIr1v+Ub1SI4iVgyjvVI5c+j90w1+ycX5fH3tEW1AU0SHccWhw/M9rvEwdSgxWNxh6dq+Jwuw/6b
UVP++NVfx/m9otCK/EERTpxUBQ9RMohdy9C01EkVgBlD4e54NtTVeTbaJwKWliYoEniWSmwyKEkJ
4r/nqJTwbYpzKo2qsVZKIPtCF/XXBoJjuHwuK7UT0xT3PTVjEpY/xtKJkUmgqm3Vt7UhS3CkOCxV
VwkvLN2nWFl17QfmADhP/+ZQ5gI7eX4ttk9qIpZQ6mgZZu2cmwwugOIQg/AumT7fu8ufncew/wch
SRNIUo8QseRY0oxPOdIobNXD7YoDgPsfdu0TFBaq6jun5wE5hTX6fczl/s3WRsKYOb8PZYI08oNF
/ws1se/wi/TtsWFeHm1135pZ0y/HLi4rzIeZVm/15q6Fawc0JZBjYW/1L2nrX6ALgLCmJHZx7Pdw
wAIhm+SuE9EbTZkFP+dNyGI81CXFtpaYwMTZNQR7t3FT0geKyrlFEg8n2HPuiZiUQfIXTHocemrk
Qho1F9wh2/j8U8GJijFsFLVwlLr3a7ZJTqKh0zubVNuQaPILXrShYZZikp6h3O5rfkjuvz/Fz+hy
6HRP9Bf2ZlLP2OeVJTp2Pi8SDX9NwdQwotOPqa8NL5GT9iE2VfM+fIDBAUvlZ+i4D1Yb3/HJuJsm
N+nRLfoRSAOzAgqXMuVxeC4F9IwH8Cw6DMIFyz1vh5j+TXCEfU60NxqZooa2+qCkD4CRXeIIH1U9
8mfJSv8vpCy8HQ4+QyTU3HGREL0pe8taUdaM56SEHV1Ei5jvHtZVcmzEb923qe15ZraqS7E8VUiQ
qoD6cdOaV4JfszzKew6FZLsv72Rlq3hAO8FDXVsDmzCawe44F2p/qOBExEXiNPUnLE0IAWnXZvvq
zVafakSAqGjJJU0Jb5VQF6LZ9zTEyCHQr/mYuNNeiikSnfeAl7hle5oQJAKfsTcPTDwUgtfEM/yc
NQlOSJOk6F9U38Dhx7ehGF9ZnErjqm11BgjlKXLyIywROwGm8mUpFgmypJv3EdGxXAHO2qV9MPqJ
lMTU2udtVnvniScvndguOJWqlAtOXFpfEqhv4Cg12SDn+YCFJLkO/WAfWWFlEVOzD/k/tDikci4R
lybHmRWSEpSmdMTs2eOeRy40E81ZKvPeOu0aY0zOhymi6GpWo/hGafJvk3hhlk1Y3pwbh8e1hVH9
PiWqy+CBfiQCWicCwvIUlt+uB9M0zmqfHYKRPOgp2Pt0YU+ijze2PZPSm1Fg5e9sxnmYg4GeZNTM
XJfXh55YjTBg1islrWXgGBZ5+B7nxx4EpdGduwVlQsFH9qyjjyHIng/EG2yBLrqEO4W8eU/E5SLI
sVvhhn78Oh0XlunxRL8UNSF1bVBOUtOouLLNGeADdo/jJcOqB4iUyobiUgRWpdXiZ2yy+BRQRsAR
TcF+oP8Y/bJFI8NCUmTTGDJNumC/JFc4Hd8me1JNrzk7l2cw21yjzUpq41NrrawmG9WSD7ZGrSGS
3H81G47INhQbkHypnhHFDRZ2muIJpIE5r6hZPTm7CdatvcuQZKOs/vLnbvtz1IpDIIEWLFtRMPbn
lnRHKOC4IGigsw0rqmx9LR4i5FaMsfGrudS4kQl8xwKJ7HOvfqf68yIOEvgvHmt8Mr7PJWJz5tSX
tl6OCpfdzdtYgpo7aBJ+m2z5bsIZVALZTO3QytPEX02AnMWrONQE7SS7+3UBKSuCG7fc1lu16tU8
fJUfSi4sg+gVysB9wsW3OMVJ1fxQwoRMFL5q/vkD8IU6h5omyKwYlnTCSYgHlNjsVq71eA4NKkf9
t6HX+TGDmkCTQqcoyAWO97zaSe3lKULTD/3Lq0Z1/sLUe2nWtjmqzHpwViQhZCLrkERwW6gWojQk
0ev3QvuB00ibfCXdwhGUeYlTuD5JUHF1i+ogjAaHlR/zYnWyviSzISAaEhpl48ReQrC5F2doGlSU
zKR4yeex/8GqZMvUX8E7GKUmMZfoZD33KU9/O56M/KrLagBmDnjA+Nc47t/euXmTrtHkuUvmkZ8X
kARRVdF+17tTBy7qQp3qgRuIyF8SCA5EVUNuDCq22cK5CRZNbpZUSvxkUUTiqwaY6jCGgN6IDKBg
IQM2oplc4Nuckx7SSgYJPGD3EdqzZNrapbifllFPPn5KHZJcvTOIHM+omuaAftfhZ/DlcUw8Uwv7
Fq7WAM00WR4Qahgs52P/eF9npNg4lUyl7JV7tfN7fsyrzAtG0EBOZu/4ZzdbAbOx3RGRwXvpD3o4
53/55PLxjCakNncZRL9xBglne5nvCKPUeBlWm+Juvn6v1s/4Yb1rfFaataz52q5WJeIGb0SSv2pb
DSp2rB1c/08mRxWEIk4RqHxSUygMQxfUCmgJjzQ9BOsDgu6ZY6ZUydIiQcaLNzFBtPJNSeFBvize
7ND1+pS6xQy+bFU2YsrhIkSPGYi0qvaCmLZx1GlYghnaOEyw5aSpr+F4rZeB5H7vkslNW+dSq1td
J4EJitPavtBbNjCip5vOAaYfP/HsEsCmym3O7PpNW3YpGqItXnvI31YtsAwF1ckaDBB2k9Mjo3FH
l8s0mHzbRmYTR3hOlc3UMAorjRjdj8doShkTAccfGr+3VsHIS9GqlSjwvMSr/dVuMSyS1WDC4Zw1
Rq8lqZ/XUVFaVfR10+O1XrGGeZXYX/sUdtFH+gVMc9qoxLK0pF2nNr0qvyBPPsVfrNk5Y7aBIwNk
qO5dZnXR1THQeTCgFpe7xpKkhkrWiI3tgfmYcL+eROUywSE6zpXj4ESr8JHciaAOMzsRO3EelnbH
lUZpPOf8hH0Pj7TYHG3fEvzosa/zBOHcHuv7unwazq+QS21UF7XME3JhqHKCbKnwPptv7gpFmaBk
NJUm9sjyAd+NyFS+H7cxmdXZnS4puykHNLZmXc19z+YFuHuOUARswurgI9ZTryh/lZ5sdpoCeGE/
I/uuGHwukWGx7+kHQWZlEeC3/K39rE75rZf0wvEtUJiFDD5TOhb+i6gD2SxQYVhmWj1zgHvIE9UI
Lt4L/rTK6qmFKivfH3S6cHmjTggUF/zOnKaOlNy0ikpAF0CL6J4G33W8i0m03MBMDeC4ycuLGzDF
qhhJCncSjmAKn4fN6Gvib1fG7rTxSUx707D33Ys8ltp/B+OFQEfxTSl5NPV3KkREbw5zk6YpKaH+
65+BuIJUABqwK4/fOjdhh3J5I/xtfAIkDp4axSgo8GyCiUbIya9lE/KWr9GpGirB+kgesXg6E/dr
7FZCtgcBYXZvs/pqkrdxHBf9/I6fmzlIStGdgJQLjIO48Vs7W1EdjFXlCDDnbIrbk/tFhF+eHkUs
7foTw7GaTK7vmvTn3QQZHqgVDZkNbsuZ1K4cqDIpNEkr24iwci5bIPC8kxgQbv3VOSL8/Kl9hqCm
HZWVtKK0IbmxyCzLhR+iv2S3FhquDK80mxGnDH70UhbwGPInWgB3Pxbt4UuDcpzATC/T92HVGkX/
rj9Ftl2uWmTHb4itiXCiMPuqUL8SRcc+60QA1Yu1Y/B//V1hfszkMowwUDaYzesQK3/Q2FF4+XWB
+Bxqm1tCDnpLBP+zEN9MslqH7zitxbA9mer1rFkBQWk/OSwO9mXDh5CCmizxLn9QUtzjtBJbv8Ut
Hr9TWfuYO6DFWSnLkTGuP1WR1KQrJcgEHwaaXtUvvnQO5bDVRn3nufVcvKGs/7uGWJJpTegmBs2V
ZL/UKTBS/hMgtobeNGDDyBm+xaVaXMa+HeYHw9lG0heVkYYCNydIJWPounp5a+7wOxeOlgUhicGS
o8U1cvRrkusXOM0uGTmvYIpThYGN/0KY4KcIZhCPQ77oczW3XQcuYXqJzdVnCwMlPVwoPfPdBi3H
GWNvLgdq1PWAYY31RsDKHNYftOvihuUsbn8WotU3UBr4wd2eVjcgSubgVAoaq54JMFyzi2ZxLYBQ
tTI+05vG/tnQqL7e0TxcP0la0uMg20cZd6uGbc4vCA7NZqOH8vU0hHNZ9cHk8M6H8awkSlIxnMCK
gbAPQTyMe1CMt37JV0pYoUoqyn6In7FqYjdapyttmTm4JzWzR13WsF1sRLOCfAJ2f/ayjBkMk/eZ
pfxui2FDeQ4AY6pDkRrgPmTeK1WagXQqMrmsGMqbGeiOm5BkguQvqyPix7ap+cWoZRHBvEP4X7Iv
iZlqH/c03f2RCZClRVJFlrmKA49BAdMDWRu+Y+U11b/caMjjM5MIhj9O1gHte5h18IalCU7lFAL4
18ZhndK22QrkL9gbHhOsomDb30gBxqJBL2hzfmNjCdVZQBqi1OzOLSkBlvQaLh8uex2hukwh8/k0
2Jv6ir+1TMPkzelPf9iLgKXye+v0ZYudbq3IbzBQ/nTfQFGNOKEXZhLSkFIeGpWmebrHQGQGlBA3
msuGwCjGzAajDd2fZsx4/EJK4Tneu1G7mIyxvJnTCG06uVHcfn4smOTU0Pudt6u81hRc+eQYn3/z
2zBM+GMqg7A3xnc5h757509FJr1BBmXF7dPSYNW6CcQlsr7SgDeL9wLEDNJ+uuaJw3UZ52LUWYby
Wa8hNjwRBZwmsjNc8HyY+/5hxyRFW+TruPfVLg9+nvGqmTrRiYYVV6g/JYbMVfkg4TFo6J7rOp5Z
6guitQr4q3dsvsHvUtL1sfYDiYE1+/akSO/v+hn0l0DbsTd4fPK0GzPzqYonNby3/wmrAGM5KL/J
RV0S4Qsv4+BXyAJVpuhCjtnqBsLUZ0cL/DHcqPIEJ1MjmOwzOZuqa9iSfBcHRXLadNCgsJ9CO8ke
gRskzeVzgQh16uYVneqeBc97mb9yghNSMtzODGd4I6PxcvJosEdKYh8JXiiYGvAeCQFv3EPb6Bkk
akOmSDAQENbo4NTDDIIhZeBIzWNaXsH1RyvBSGzXYKTt+fqzDzhzN2xQW/74k+73xoJsmZLDkFn1
FiiVsl3GU5u3/1Tg+arhmB1VY408wSg678yZKTARZSKSCCkh/h/qwMcXquywp28gZc6nb1eqOnEh
DxstqO8+DvovTzScDr+i/103Y5owxKz7sq1ymbn5Wp6Tla4+S0yR6v0A5kaSBlEXFb7Z9XOrTsJP
j1T2tK9Od7FO8mYIHh1bkNddPVgFZGyoRixrgBJVaBbBv1V6rglAZdzKeO+AW9D9UyvIVmR54kQl
yvSLpp+afyWgqHi7EuceXU7yIA5FVrwq0WGkyYAeSaKOZivx0tj4adTV18HbtKHut5JkVDd8MdL5
KU6xNyhfLRQc6DTd33r9wskAkI1TDF+AN4niCkqyga6eV3c1Chul9/CVllucKoTVsT42yeQsqCFu
Y3hOibcDfsiSeeD+jKLKPAEuIwfjNBcAUC1NRz2XatW4RbBoUJDtHpji1NoumFobVU4jZN10jIiW
7drHGy23m2MP8NL5nU/kQCRQ/L4xWMVAGT/ERf56gU5KzsnFlPZrLfnCRMFNVMfVaGActZjv7/+S
F3cqcBhQ9KoE0jVOa84nq83rEs2mGZolqTXcxwHCrl2v9aQJ/eSQtqBiMFLHsHdK20VNQEVux6Da
4+a8Eyi7XWJv45eJC95SmKPeFqJpqsW8GGDVpluGjytGyfSouy40ALewPCPpGRLcsmSrFOPEiofa
HWU3TRmOgH+/JPY44+4cF/OyJ6ABZj5KpD9+3rTo1aE49WT0LDrwVCK56ZtzU6/FASH/aCDdQPZD
GORHolIqlM3+my4XSBnFJBTaeg5EdvpMJqDMufaL/UJoA7MeHnFb5SBKvW63LuN3xQF1qFONeSkH
HsbV9mveF2zCnPfwJ/ckD3+qIoIzQPpiR95x5JrQHRi7tmPV+R7FRp32L4q4eMdNPS5TUECfO7qg
tops6tOtB6OBr+3LyUuLxMBkfouRBKAEPRcwXiqXtTa/9+cEEePUiv4rbsG7WmzubnyN1J39CaMh
arsEQl1GWzwqEP4Y8GJq1EhHDIOnXDys10HeifahouM9LKtYbtecuZkNpc7PdRz4HNMmeLWVa8UY
Xs7SbElW24s3nIlUfMM9zKuD58x3/YH4i2IiK0+tMlAaYaQ+o7o9CwrSYstPS2/P8KMdBErdsDtd
F9FZT93KgbqbZLDfCFplFurOFB5gEtduur1rnhSJIzkpFLygOTstODjvDEPRV/ePI6q7XPnhxV3B
qkCSKSMgrxSRSrT+yxa4X2xy4dJMYjv30GTLZCYpOblOQe/H8WdQU7vzNkTwW9lxJxMSzrtK11ue
0MwXLpNJyJMcyHfI8yrVZ0qsh4uOjr1xnX5vZiMSOrlqSIEkzW7wltsndeBWr+0RPunAeibnznRw
XyCQ0T7nsvSAXcNQIQ3oZnurVum8z0bcUDvCiz7crxSub3qa1KiMajn8rkHVGXZvrDEjPlQFrqYX
honJot1WzQpxvbOvcj8/8FEjcJolYDE15nonUKMC15+NBvAzH+991Zn3u/0Auo/mHEZhAA0lM3fp
zPehHUbIYtkCcG0Ivy4jYb4e8//7L7iNzZqw9fx61RJrXAQt9IA969eL3Py7QVcYRCAqNKnwaChS
G7eKnrpGIOIpE75GcY/anAV2Hl6V4iAzFL6s73VXDgK4pXt4ldL66gs57lFTlb+XJxycFikKtBaW
sf9PdR/qteOjAKd+RNudwI7+TOrXWJkkpjsafjlp8IfOMTFUTXDxdPFRXu2lM86AV6SvhXWOE9+Q
XLIGAsihwfblmpnZnH/3WjnSha6WZ00k3bQyZgiwljP4chPZZhtXGk0XhCHbDYJBF8lmvQmwY8yJ
bE+csZ5EgZFh+WbNga4SzW1h/+Ye9IJWtTg4xQWdjKuBAZh6CQm8XGVIluiOwwYBSt+Xnw/Bzype
zWcJ93aOlQheepJFHaY9SKVGmFjuCxUoDpUsbi7YQySRNTZWO9hYI4TUCp9GPGzW6f3TsruLveao
hMnVhWIGtDXBH5dqi3PfWxdq3VfZ2RIedysvqQccVUWXUrfB9fsjWlBpIck74Y22LgUon84BZRvh
7TaH0YFq7UiUCGtTxAlHCNt4xQ3x8LodfvFPqev/b1VyHCpb4CxRgB4wJKCHh44CaJfjBtA4ovc6
Oc5t/u9mb9rZPaOclXQhQWLGVcZ+ZDaMwJMgYXKS7vqU01rtxQWizAv8gVLbWW8bNfcbn3SILTKy
sR+dulTMbQ/zkcNbtUSNgp7NStfz7sDSEJeTMsg7QUbhRJPa+fMgVw9IYnoRFCv05Sx7PTFNrx2p
H8kKwM7ygHtu4sOWb+q8Q190CC2Y+E2nY409O0zo649l8E1qSFRniPhvvaYm7fGCFy/1ZWH1LMZG
Isfl3G+f7D3rB9zOQFvbnd5GOfTqrrexMRl2Asefg+2I2fhf8uiQdRjAJ1tZEUoFBHDKExFL/fYU
jgGcs6UjYIPY20CoxDafWPyT5D2gcWW+ZmZHgyBUwfyBQQGQAvxpayRoCvz7dyDs2ruZeMesYJ5E
WzbgpZgJHM2eSgxbilLjhseMaZEOrByVEnidJftASDZUcG6Qro8GQq1A20TLRBnwkjqH+m6/EDpG
KdgBBdbmFxWFjpswQzeUfQGogBTss6ujTSh7ckwhixiZhjxYpIjA7rmJUQdsOK9JBGQxmd1SCcUj
C2hOadcb4vZnIX0930NZRLNdT6QFUpf20p1AZBLMAdpQ5J4XjtoyetCIOtUxpnirK+XBYCt2jgpy
1d8Sf0OUcHgB82HhIOtF/JEfQas89XdD9NHMZo//7Grljps8eDo9qQEHlBtnW7f6r7kzDqxXr6FN
c5M9ZD4L5JQmiMB8FMePekD9UznchLH85Ryrn07R/GNVb8APfX5u5zKmvB0kGwZXesUmMn+O3e3R
uWyPAY+p89xA4gmSTWnd1GmV9FVtWyXHyFA6/wcbUL5+oIjn8Mb2Z8dea4IRo2g/3FS7bzkBgcoq
RPJi0v7XdT27wPGqM9IZGEMM5bXujvXe9KFlMY7vw3vyJ8YNaqPfRooiRv5nparkDCIM6ISBPwgd
QP/5ZrJDO2vYoTUegjufYpL3QiCX3dA/h4wXbSha2se/KrF3B7Iyq3IMrIi8QB1YWPvwMUIqYYGs
Wxk2VvKonzs0YxTWYz75ny2Hx2NnC6zKKmpxs4dYtN+Ovsf5Re8OuMbm3BRpKBM5/Hv3V9DzP85K
RtQ8Cj5gKfgXWuY7OWUBo+MHN+3ObDrYk4wsU+wrWYksrbUC5yIC2d4B31VtCBOmK+jtnFZ8i7et
Ea+2kZLx4PYq6AT1BbFH+F1BUEEWtjK5meKdhB/R4uw52Br4m5XzlM16kVmPIHnJLlzN2DpOaKWa
99mL15CkPhrT9R2HyNAferFdbWQxgH7t+QPSlyPk2PsgEnN8sWqGnfEWM0UDohmcUo5v6B/zml53
pwbBRBkm+vASVkQXrT+pS5y38aklN5iLBT0J+tWRrrZ8jqBRpecfxns9PeeKMnz+U3S52KeRDo3g
4XkpT98sOH4M0dOKbiT5FY8vaXlFn3yAc1ffo6wJsUtz+MjeqaANFM7S9zUL4mMgIqcdKZnC17so
M1/v2T+NRlyMqtFr70aDuF+TeGnGdQlSexXsuWYEMstJlelbNFlPZYf+hoSvK5sTQ4XCvKkagqUf
ZRW4BYFSWpdPK1vsiNASRivW5m6TFLs96UB1Ql+e0NlIRyxfehut1nRQi11sW7j7uSCOmjBL858R
OWYVGjIJ6g5d6TlwOpyzRdU5ELB8bs/wUloya4h4N+UPGROkHRbGsZmCKt616ASfgZofNcDD7yQO
nIv54H/u3jQvkI0rytfxkGVmPTcND6UzrRhPVGLIfyqf0D5eoPp1wswff+UxezapIWR9MLihdvPI
r/jCbA81l0RMSHqKzp3bpLDBWNZPTdue2hQyuzsILEFBHEAWWSHLTKRj2ZhCbMv821J6hlaZh0ps
DBNUZda/cxlrDb53BlT0T0m9SrBw+eQsdzH1vLfcB4mcmW2pg04yZKs3naaZ3lH1wU7qmh8DMRmt
IITiJN/tB6ZwBd+F873HDb0LKP23ymItKWoDNAdbtUuG4yIqfTRG+DtKQtoUelOHGwOL2vwSvA53
NOIicVaIMvNy0jbmNmr31StmZbSx9KCojY55yUAKZbdM/uEbAgk/qMju6D+AxpyxfsVY3L8MJLJx
NGkNv1eJY1lVkoRBx7xKFr3sHdSB/shIeSivSOAhrBudmQOzaaY+RSSr5z0djEfyifPzJ6AGfwln
gre2mIkZDHKOckereMab7+r3Klk8Dq7jO2sH3JN/56/E5oVS15NAjVLjQsAhvyBAb0Buy5XT8nDZ
cut9e5MWViMjlLBv0QnJdbg81rjwHdWPTCqo6moek0A20q9DA76Hpiber6CfhCIqMgSOCA0RZc6u
0VEDwrO+5vFkEO8F0MKfw0TQHk3eGJrbAAwt1oO474XtXj6xrZ+Nx2SE4rb4WH8Xc2Z/Lvg8DefW
m+DssXtYs88xV76J1lMbbU06qncler7TWJIV+LXI7t6wbtf6XK7r3n6LSR/jX8HyOMdUbyQUq6Sd
O9PhL/6Ap7xXKYoocuJX5VrktmyrN7HcH5YR+d7SxDwphlGdKnXU5BQ+0sbIK73dRn4qwnuN72aP
hpZ5n1l4rI8RPTiK8zVJd+EGHoQwdUkDVRmXMhxj0GFkHTID1IhyhJXsYTF95YcLcp+aGTiuuc5U
QoDJNXoSpkJiR5rIQv6EcNncc04/Ekjpa7fl4091kTfCxAOF0YArDGbTKUzITXHKD6ld68xUKWVV
f84qqonLUNIOJxblt6YpsNRWUXrV13gDbjY0IuJuissWBQ3UeyFf7a3RtV+SMYojfNijshzfi7Z0
ZYrdC/LO6e1YisRanbYpQqto86yQGrdvvs+h1HJViosTEAXks9BbjejvtQbVlBBUpCTEnYMNdaAw
n5YbS/QtLFJJfdawIg6Z6YAxayJfV7tCrZbMCL8W/QtSEuiNrSRqDxk401qXIqf6xWY7i7cY9h/1
PkRFML3i/TDMiPEdOL1nTZB7GJl489yanP3Zg0oLHqkOaaqWnvG3cNk+tbrygju7m/JPKdubvSAT
20QIWDHgW2Dys6m2F3F1HQC2ffzpuq4Tj16yiFwtaRn5FPoZTvfS0CfvOXpMU/HVEwvr7fB4zEV0
B6OUEixG1RVV5U6dRCO0EHdFaI8jC40/WDoyo3gdWFjoyFpUK9I5zItCPbaHaLsliYMDtfnvnFQJ
mVUiDz7DNbpUbYj6kv9RKD7lModQSc4wA7shXpxlGUFAMYBPeeLK68LJ3jsGkUM8BuYyx66IyjM2
DCQ8GofSuoDGUqDeITIWgCYe/c6/N1u4B48GB+WNx2GHJoayLm5y7cf4nAFDdN8R/e6q2ozXB+rD
0N6/b1s67YP2Zxp2wg9cvJT1S4YAqEZ56gP7tAoPnVZ1/JBpYaSaDUIFcs4CvIqiN6QEPs6/0woy
85uwwzR+I7LXdOyKhipvVqyxQ3yKb1UX2RN5xeL/zmOQb8ZjLdrNW7RX8lVqxUwva2DvjV0DFvTQ
QkYKSlCktFMvjfOfCK3t6wxFOkH/aviD7ar6Ow/cfPUPsphm5aMyAZJ8q1wHu+c/SFb4vcxNKrZX
4O9r5bvrw8wrE85QSQAI3sRE8ewmD9FSojfz+QIRqTxVHz3ZfVsTrAsTUvmp2Kjn57G3XOpgU1x1
0qTVYdILGeCO6uqdQNK8PdD+49nuVxhi+rYy1P8bZLxlcLqLiGtXjkEnJtiAX8SlMW8CfX1jrvIr
7asAB72dyRPuwGhqXKtkbheWmcNYE/POK3UE7Rmz+LZDvtxcpQOWfjXkr0hsAKzkMRZqZJBRUkXn
xR+NO/5AMlesVGfo6jVW2mEys38Yz1cbPjK8q/TELB6qa1q/mVumBI2pP/bGnWv0v2qPJnlO2bLF
mJC7tAe4jHjI9MkinRDHxq+/jICpL1zArXj1goII/T5s309gEMgUXycVDnr8P9hX/3E/Imb4wmuF
h8oKo4k3aZ7FOw+MOC4vu8VirFhfHnr7tT4RkTKnrLG3npkqAgul3UbCJYNcGJ/cbFFkpl+CtxLV
SYER7x2jJ/4cvDugyU+eqQXHQ2M/Fi1K/JDSoTz8/trf6ywYdBS6MkQMHNqjM+Izn/rdzSgne4JJ
baIT5MsHZIqSBGJjHkGUk2QPj00+x9xuRFQbB4i0J+J2ibSALaHI2gN5RbI1Oov4JwmUXN+PjMQ9
rda3yDE5iNYBj4+khmTFjVA2ePEVfcAlQlb1rSjfPBXpofIj2+RUkDiYWBT93hMgNn28Vz3yd7nF
OSAttu1fzRFv6xrblRN08em5KWisZPJwwA7lX2gEHAX08vAZDJ4iCjSFRYvGcHsE4busgYOotS8i
lT+xmaB3RgZpIRnrqP2yY0qT886v56qXUbWHKYv+bKWSI2cWTmPPN7qsV1X458jNvMylPxjmWj7L
w80TKjNyR/IKufQ1Vc0KCTkvKit6WqTIfWb0fml9CVG3FQEL8U13TRwB6VbvAvZP3i0iFjX2Elwn
AnbohBYOuaKwwdraDuXAXOOivzoKGpGotMsBnXyWThb2XgRHczqhEr0wdPXCxumnaHeBm3rzelrl
olYtEJU4VmNXArbeVE9/mVZ1nS0ady4n0WSVa4NA0T+H3Z0dZwepNBq24NK0lL2VlwwBhh0PPIGT
xvXSRElAFxLpXlUnLfFELw7wz5jKLq9/H15fuAwbym+f56kEhSV9Ynhyv7d/ermSI+eKPhcQ1nCL
LFrtUfvRRgDCX/93EloXugvdRZjud5Pb+Qg+FOUqA4DpFIc2f0lC6XM9J2OFJHX420ul+AANhLzq
9iKYgHKAO4TEJk8ByUlPyqn1qqPyo2syTdr2mzBtSjXuf8CHvjooLuKGfLsVcJQrf6wUgfIlISer
2ssmjK3mznIUNyzFw+2gThStsitiJq7NoH/BBArOeo3bwXSdOkpDtF0wRdllYnWCyM49CoysQ4ea
36VZGdLKNXp+gm/gRoqv4rK7isxtJ0Dqbbi0Q4ppX3YfdV5uhHXD+7H/3UWnmZD2sxu9DvWlGVp0
rlhIl+ZrIRvqjNTK7j/wITimyJbBZjdJHdy7+/J1lauu0iNIwy36RrpEbyrRyPiewzx8KO0RbYxo
ClneI818MolrqxUqKnEzKoklUo/+lrFJQkd6soe/rg5n7CrucLJainQFKZUpqnDeCujIFpipbQyD
iuLbLA1Gr3m5Zc7SPWjbusw0rrQQDmhPjzdOl+v7yJcraOYoa1i4jpR6J1bDUPeY23GLa82xZQhl
LBqzsCRFxzcliSMM0qdAm46pEQ8bITXPsvzJkyu1KyzHElS+0RaAWWPbD8atdj9nYmv42nrjMw9t
fBolE7uRrbdKvhX19CHlZJEaPIiyYgC9gd/VZn3z25B5RkX19bB25zvWYCKFzxbeWY4yujg+Ha/t
wo1z47MJ1CITltVui89AQeHyefTeG3oim2Ynl3oKxf15TUGWH0SazDQ3iBEWr3gxk45/opSyMQB1
SK2kh+LQwmIRW8rd+VR90LB0WdGIw02Znx5GCRWZz7PppYsojJN66aDerkN3RLPg1mApXWg05xGX
BGlaECp6+esTPC5fHUL3XXSo1skRiWq1rX+EHOd6wgczP9wYmVFlkM+aJOzTT35hnBRkzhuMtaA7
TcMBGVVpa2i8MzzfCIbigKbNPzK5T5uDfJKDeCk4Zbnho5xRLg5fvbKMh7ppN9nUWRPjF/PAZMGT
fwmO2E4SdvZQer2Rhgx10+T0WvMabZd0tVg+2kBs18KnVIE9UD1kprebrkVx4oUjIwh+TxIP+rPn
2BEzKv7qOgOxNb7+xUouzFMnXf5X2CA1rYQWZ1GqQAkLcVmpdZpTHA/28NoN7Cxbs4znI7gApf8e
CgW8st4cU1oyjYydEmmwyZdI5XiXWTkikrPaRzT4NRJ6vbE1RknPXvjIMAyBEfTK5iisflrahStj
U7w1Ym5U8O4u6SwwgZc+ILIzlRgCSOAZDs96bckpklW2XzyOF+Uxak0GWcEfiehxPTo1d6a8PfUa
GCgOi7l7VLSBa9oIxVX9EpzY/UhHMpVPafDrGWhtxy6W1HAtd9bkiffm2EptmK7eGD7jjrQUyShN
CdU0eCs6htBgI7ey9cUQjtQbgNgUeF1o9Iue5LSwdn5bDNtwNHAZn3wo8MmXBNweXN15GW9sZCQs
cAk3WjgM6uCyGYDbxMB7oAq/0WQEVPh52+cPSK9jPfTSdIe5hqfj0ZmOvRLMTNr5nfK8hiMhKFB4
2y3w24u662N3jUtykHjFTolb595g/3t9gtWdtr6hwBR3KA0Tp3o30o5TiiQc2Ipa61EJdiPLIIzw
RNhVepmtiA5Q825ow80UoflMgy1SJVYGbynlItlqb7UHb099P5A3nTXlyXvSJbuKe2dPrUs/wemN
Wj4V6Bh0QTEu1gbfUSZwwJPgtAtkrwmZwkdFSRPXbXFPgoK6mEEN6iB/HcLWqGUuzNPH/Zt4r0K+
vJKpZWZ9fBzcaGRccXZV213CWp8nxSRL2vrFvjJOpyJHplM2pHsaClnZI5S+byZRiwLlwVLmcjZY
c31HNrCXJvtoDUij+mv+p0llVdNDxJoja7kEsq/VXgWnSEZkfQ/zrTwdgZhRXhWEmFu+zW5D9fHe
cujBYPdMobKuG0eXOXnAe/se5Aes9Qq3DqR+vdfL9psei//ZTgTRXXHcMTLSvVAhAVwqmRfsW/VG
pdswwpxSfvQdBV/rGEUmfsnfzLqdKtwcRlonw68CmDKV1Gu2/Wsf8N641VFRY5owwFp5B3W/866r
/Y0NBfSdzOM/067KGm31Y228mtGr28UN1zMBOfAU/zwDPPOzPEuYsJPMxQH+oYh/2UMjPZbk9enF
nw6PRufwf/y03y6oJJwuzB/Tke6hebmlB8rQvijxLFGV3zP7/4X9lnCX4hqpgk4Za39L0kEBwjUJ
tG4voUMrpFroCMJ1UIZk0gh6Cpoij3ndcgM4fV9uY313JyHyVwNmo4gMC9dCWRF2xZ1jdXUEXw44
SAYX1wUsq44IQPvtQ1ssYID7ZoazgJ/RHECADUDu+BEONnO2rchWV75uReYcfiiR2EP0VmH6Kt+g
o5n9oYgFTIS7N5c3X0iAzuIzm73coSuSD5hs5AkL89rcjXOODwJIYfJD/p3lagrs5mbB6/6mKIQr
cJV/zMt44IOttWCkb4WoOBHKVkFsJBNkHT5csv4cmPAo3HLPGx3ZMrq0vOdeiQTy1aZMzN18RFpc
rFXdnUUk4lpMOWfzD4IU/5yVlLX5AlFa2l+gkf8HhKcJaoY/kAAKFbMr7cNlv9T+ibc749qUy15i
vHI912/3yVOCpNqbjFNXywbsasLOLmpm44oHVedi/Cyv2RtXb4NN7+BJaXw7RuaVYfzooV2iD15H
Wfumw3da/40YLm0M/hSbSFp8lWw6r3Nhe8cmfkEWgwXWlpuU6lTgYctb5a/JN1hiRCOoc+O6z8Mt
CUb0yfqxjw7ciXzlCGjog42li9yGrS/jtcAQ4UZODPr+LHhSDQbVfErP4D75DuJhNVBFs4m2mUOe
Sh8OstczuHF6bTpRIgPRU8I5wWZCezFl1gJbJONwFqaQXW879DTVYpxUVQuYTTrXZkxU6cxYjLx0
3nP9JoJNA6e/xSy+XTksmkQaV9m9E3u2p6u2yzQVMqxNKCDpjjR3Y5KlE5MazwZnU3lw3TRE+mtd
zvaVXZKLGJilA/8fXVAh8iUbn8DDD4TYaGLMLosDKP+NV6aOnNwUsFHxrkdH8RnWAcqHGBvVCltM
Uq+x5aUbSZGO+jOUoqIhj/EH24hmmcj0K1fE7IRAO6Az3Le81CLR1Ea+MrlE5y74iXCl/VTFr43J
eWgnIvrrolDf5n13+YGu6+w64aWg9qz0PBWpJCPzYWcwQUMTw5e0G0jUo2ZMlWvLw0ptycsSF1eP
940Dcj7NExm94ur1Oy74aCsnhRYZj6HNGCR4DYxdPqOFfCdzrAKV84A9dCVl/oNX9ceSbCPKZ/IX
XT1vYAOfRCjcFJb2srmWoB4G+QrHlwd0jO7uv38OI5fA5gNJiYNe51QRXYtbbT3rt3E4yLaH276m
HqNFb/t7a/pvOpd+8LgQrIcpc7GLLi/6IKtQNHA9tgHjxYI5YQQDF21Qbuwj35YeJoy4fPthbYpJ
59DXm1gtZtscce05usFwTdH9riVpBrGcVxzIr/ewrR28kVNUwmU/dgORxcYTFcduEs/QJSkGFNIr
bkht4krQz/2012SEA3ruGsDxuEECxg+KQP4JIe1RdZQGgjrPfg1s0sqxFsIZ3VQ7rtpDYUXB4emc
oh+wj+NvnSbdwD649acwTiIjlTfdG8ffa1fr3qn8xRDwPmIR2NcalVdsX/450pYKymTmfBZRtEJ8
CFmXFOWlgJ/hfxQOHlltAWEBUqnZhqRLpz5PhFcjzxTHDRJoxW9PNkeDhOmJj17Km6hQCODEIzjK
9weyIYW73Me8X0lBUkDZbWDoyERs6Z4UdOS0+PUvVbP5YE2sRqqlpkuCKvWWCGsebnpX/09gTVpC
jOG0dIMY4uXiA0+S+6pPDUzKJtU6T3XpO1gRgbkKIjXWjfPmwYmqOQ6fpCMrykEcCf/CyPOm+/yz
qgdDDJZgfNQYH3my4NSLlOZJnZ91PK/b/7luO40N2KrmoRXfG5NdUDRy1d3dPdPQHZXKpDW0rceo
2rqTtrUY5dkvMg4OKaE55OR0CRWuNDVce635si49UMgMX4g+gwDRfQ59Q6XbY4nDS+TcOkJXA0DN
hUFFXqyC/0RIcNXjHu1B3dUnfnuvYsL63Io4Sd0vfGyRh8Is2hMOvXXSuocq797TiOeyUufKi+TL
ErL8XOJEDzHD0k3+ac0shRDOFWO9RtUQVQXpSQURzstM6YM+saIoO10wFQMW/cD8KKqWFDRs7Rvg
G13jW9IutQz5IAQFvo0UgbjaziKbM1kzJ+qUB8MNkwbw+MzXm0Bh9rK43RhKNdF43zujgL09cFiI
/9LuhyTQ6SxySpGCp0JDjUdW+201K5Ymv4zf5ngg7eUz1N5f11KrG8jO+4m2mD2IdEX7jbj4wRyY
58NiryQ0jwBmTWPQ69Xq2G55dKTyC40Vn+1OJcVy0DAbsSI9g99RE1jIgE3hFVl6tNmiQ2XTAW3r
rBcWpaJDiAxRmoa2W84Z/jXbxpeEImB7Pr32cMgVuM474lfdf4+6n9n7XQwDRpCQM7d3zpHIajKp
N7UNVWEJ10xeYCaFVctsiYzM1ZuwxvpDzSfljaqaBiek7Y3kSbcp1tq65L2hHbDlx5pQO5w6BqdU
GpJcMefM5fLLMFjFLvf6p/WGzDgsm0zTxjqRuXd+neooe6AkpwHlyg6VCziq7bKrjWwmTzVndnPd
i/FK5p5UCkvOnuKrxC/EUv6elvGmEbi1kC9kMmGRtg2b5yBs/WQmw0lo41QWrs7sNortIBMgb4+A
jrlM8vxpp8N7f2hxAAcz8mc3nAAsRHanXIorEQBVQLdSimuiXaI+/AOXga2jU631CODoUfsck816
zaey27R0QMfJ1vXnFt6N3ePLfexvcqBZqbbFr/M7m3f0GDqEWIIQ4prAr9W6WG1/p/fCYJgGLQmd
MQTG8kU53sMehU9vBewU/yNc0bySUqLf3mjNQh1rPymqBom4ODYj4SOsEt4WwFLolCFbzolUkAHO
rAnISGIvl8GzhoW1WOMyqI3nFR4sqbcp36IzJ7lrRVVM79329M9l2OgfTaRQN4EoShilexpzHHrS
ylp1zkAUY59e+KWBljW0JAVYGpUUMXGcW1Pug/CGFexQzmJQRFeUf5m8nwu8JMnNArojZFAf5sZ5
kN9zhoVVx67yBho2rp8zIZahUny6ZcaUp2s0O8yXvcSzYmjQKwVCjJ132iIVi/oO6bUjygyPh/Qy
S9toJbdAF9CnnZz05H6fWtIEu3VY583HmGeOP+Oc2lEcNa9XzJ5C/UzrUk0jxTuVAinFaB372c0c
427d8aQ4ADJ6dQxt2ZYW9cL8DIy/VLWHGbWNBg0/e5Gs6jEWRnryDf3svORj/C6fZOq/Slw344On
yD85sn3cwKRfH0E2VgnlnT+gJvpF1jUN02HB0CNBKjngaIVsrTEaU3kj5eSRIx+/9qLIMtr8d+wv
bKa8YEnii2ZKQUbXX8o7khrIur5XRyEihw8TPl8Ksi+a5DUo6lsC7xjyJls58mNXIbowvrnym/IX
0hgYH7r9sjTeUNPyr3BVzy2zT6cCIGmUMsMDnT+nSb4biAzuDDj9zGj8F8EPKa+2A061L2jR+RbN
T1M4tGku/YrdTEMZKSQv81tTO6nSx/wWxsAEP/HU21d7+AyhcO/O5HLenQ21Fdp9rajb0nxARQWU
a2ij7ItqmsYlpnjg8OP8TQbDXMLD7vaxOtQMjqhp9oOeNFy95fjFVTswkaiNoAQa+z5cEfq1+ZzA
ugY0DN8MDEwFaj7E92lq+k3ImyQzsbLdSJiibb2PZ2lpNwBXC72Eabkmh1ATw2nyuVY1XuAnngiw
Qk624xkQ0cNSbS92RrDqPpVVLnw426uBrvL9q9H+INH8NH2faBrTkqsktdtWZb5BkmBxjB8oM30P
g/SItGPkkmlftCRhOizXzEJAGTtVCZU//FQ4V1pNhogWnnMh5iukNjINJuPgYt59XOWFCG7KPjyb
bhgfuaDDDWpu37zflnTmFdTUDVN36DtvAy/z5c5T+10xxS8g8d4uD+9FnbrlGprZw/zDgoSbD+Bm
JBP4hKKWbQkeoqJwtcVeFBAHoD4OPAoJO8/FzuZeW960/P+zL7oVt0TFnenaWvMTQqrOjyM6AqQh
su6w7MrBqpxdEIuwOQwfSN8Nfi03OQeR+HZKxuQ5smjnF7suEXnSr7LGrqlKZ0DH5TMM2KHV24EK
aUQIN4MiA9OxfjxUNfQi23S/S/WGtlpZHLv8On9ysGK0oP9Z20whRt0chpeYQ0lXB7lIeC3IOuc3
DBsoEb/uXtegKFXTbMFUwlGLW8r52oWHDaHFSVeHdLzZzJqJwU8nBNpDXZzEmedZY6V1KEzBib8v
ol0Bm+6a9ratMdiErUjO68i9O/9JQk5Nn0vqH55yfDNlEBV2xCUZttdJd1MQ72TdHFD+dGSviSgh
gkQCHkir7n3vpAWiEKrYwg8d8mvocMSPw6ONxR2fHqxGuQ6vns5nsFLRD4/14o0lJq7murgw82BZ
dtf4OeUi4x661eAcd1kVSgkmkMGoX33W3yTZH3c0e3Ojuan2wqV51J7ACvWLc2GZDH0alWgDRaLq
87oMbeoN5Q71OtDlxgwF3Kqr4yjYBS8SqU84hGjGjlKrqTnsUU0s9sqhtMw0Fw39o47Qo5Vtq/Yp
WJ4AbNp49uJ4ND3sn/jgryXAfkAloMrp5QEVQzIYyRYQq+DLIZp1VRXNF34ZDhZkbOj/UCJnYyFC
4hPzPsdTnGjWCb4mZ3bxvkycEeappWsvbKkz1AcGj9SjvxRzNlTKtdAYBTT6sp4p8lGpOLNllkSP
dRLLDeFhPOUFA4XBJHhDOLPQhSiZseFQ90UqY8QXOxYqhaQmGxa0vOzyh9o/OGuZTAWf9u6mYC1d
3E6T8oyaQGfcdo8mwkdXnmW0YR85RqZCgNVx2S9ewIgsdjy6peT9NmZXpPwY4nmR0Gc7WoguZHi0
5aT9Yu0IEatt6IP714P04cwIe7HqmNx+6Syq58g+/1uQUZtnMWXLMUOzmiTejZyk4mcfTblSerl8
HMiBpWY5nuQa5N9V1yP4hNhAQ8xqc6HQPW47UwHMguXZRxYl+p5O+y+80usA94Yikhdpf93pvGxb
L3Capb1VpuKVJpHGC0jlag8Y5sTqIk2IHY8O1mvmhpvz5pm2dM3syRHTbeBNsCZE70XqgdleCl+s
wPpMfXfjCNUaPFrk9cWaslKEmG/AXk0oU1g49E4ja9jzcjeKIdboimKePMfB8BfnxgpSmUyRLGBs
i0CUidKLDtFhlG1uIO2NLRuejv4BIRNFi7x22cE3m0GJViKWexoPSMW2JlMFl5wibndwV9dwVuY1
PoaCC0aZGCoC5igmGG93iWCK1pPqWQ9n2yapMnSaV0e0/o/9m3TrQwRjHokLl9cyPpuwaEdQ/nwM
Qcb0/yPdAOIf+H7ixORYi0bJpOc1DMaP8sUz5vk9JWGBWfb1M7+qQABHZPIrTUKvM9xyrcvh8L74
60wJ/+/vA+cwC+n7PLNZMw8W4bPCitB+4muMN07d2QnWfsKZsRrw9sEYmoXh7+FqMi/6p8Es0vE8
wtK1bgxqsXBrB3HOmde/7h3mL47PsC7pTHgxeaB8N/S6RkZhU219NVqcktPYvETKEM5Eza8KkKYg
ATgAAEIPqo3aKB9vgWHxJSUIqjR46TbLeE2DkjqzjnXiEFUfnpAy1Vv64+q3ixJtDPvXjt0xxXq9
eav4VR/n4lkzpLXz69shKp/vdKsfZsuZLFbZ6fIMU9tZhFveXDumwlR5tGGLjdZUgTqXdh0Wpr6G
XFdiLu132qe3TcmbOtr4xL/Q8WlaQSFXCyTJHr/quC/GrVRAR5BndFN/EcJjhg83ctMvPghmMMGB
qZo46xZfs4vng9GJ/C9KVANdHBnEOktWtXDhytLeeofEtEDQMEZveDgwK+w3VnQviFmXTZlud42m
sIlYs125RQzqgyWXi9Y78Xa1/xxo0CfEFsZGWi7XwPC5kuxCZC+Hbu0opjEv6GoZZmmc6XjfcWg5
9M4xNnFMxysczJORgj24x5UrrOPPH6cyTTdNMDJ9lmnNzoV/9Je2NSn2CrCID9gioZ1wNQThdSe0
+144BdZGrBsqi6DiBDy6L4xy9tiJn3IX8Njo3xppWuHyHjdXpC8ovhX5MfxgQU+gR60FrMCHjeVl
eUKobr6SirUETOI8MIZovkHNPAcLVdztQM6eH08eUvV3g903xfZ2DDqJjZcTektG6g8sR9pYL50b
yEk2BnwrXV+dT4D3iEh84Dbpat311jvAoYmVndm5BdpUGAge1srAST1ie2IE1pxwVuwyyxdvDZ5z
C/84xv8XHcIqIdZ6BvnXYHfM93gOcNd/riByCu3KGfwWpxfDdiSH7lq8VTabTZNN7Ss2gQk/UgJR
H9Dt5PPPkL1KA1e8NfkcHby4Zh8J0GzsLRyFF3dQbRaERJ9YsKjP2/feA5JzwSf/xIEJXNT+3mE5
xKnNLy+0eousrlhA1C4ABoycM4EtK6AVOMCWb4FQfsaSGRO+gmZBOKYwUXtalQc8MpkWMJ2MHMWL
lZ1oABh7MxtCfmwm1ek3bfFwroJSOMTKCgfmhDnD+6iRW05Rb9djBD+WmNxRC5N/qDJrIUdqN9RS
363OHX+znYNx1DIJUD7kfKYofFc6Nw4KGFTtM/EZL1P+a6D7WMpKlky96/0pl9OMaTGIsjDATXpQ
KBSna8GM/LCGNdiDO0BSPvdTJ0WLYYNN9ebUDOHCwIUEkZ6KAJ+LjlPvpgot8UP2mhiK8KepMli6
E/cjpdgEbqYH4BnpPV9AP+HAtCe1NeZzNvgDwT84w123jf1n2kpiworSm54Kj94d3nVsSIfvstLD
LX588Yljz7vLsFpfLtjAco9W+jIFqHF8CTNh/lVNiKyDlzDHA8bMgjLSrUofN+8BsDcycHsYgzJu
/wO59NPS6P8TgbvFTNCl3GmvGCDn+XGYgLyZNUb9ED5bWnEobBDSnGCXoI4m+COj+/eodJLMf3K1
/RorKkqZxa+hzPVFrs/5/1yeLRM3j8vh6RIRFeeG5PQdSDpFdIApngQ7toE20TZwEiA22HKDGiZZ
kfTmTbRudU+hTxxwZ6eI7qetrpGA8Rs1kL76JXAtLXQQTgg3/rvsyzA9LzjCZZoCSlEu5Ev2Z5tP
sQIkMRcF0C+noftBZGBIW1qst+YXGGJ48b3EDz6rbGpwVz/bcyxycZ/KhX3bthzemCGQdUctaC0j
3xG98iTYUp1FPJ99Q0f6dL+6vtJt7wFV3hzQyfVCNRD0eCuYD4glIMILGgKLnL2v3p4a6PxQmHBU
ym52eCIV5CGeECLKqz84wOMnAVu8A7Mag3AP4XQxzd5hjQwJrNf9UDDire9kv6RUqvVAylHJr0kZ
f+4ROp9cxm563GvztXFDRjkRfLD/ckV8EfyL/EmLLiTBEu/k164o2YcrhMKPzO2yau1eOHkEefMn
V/8CekVsDoNyA1JI+F6/wO4a/2RO/tpZamH76wWtgYDJDdx23p4Ky6DRCCBXTvC9VXI1jiRRBoW+
NJtlKol+xV3y/OYN5Q7qTuaG15hogrEbfU7IHbq7zvGOIfIQP7CGe9kmZGbNApfBoeHYchLLU84j
/OizNvs8DeNQrR4mTDN3hqBYZJwMBuz9fPtm0mdv8emhOcO3wfRtfOor4cx5ort8OW3lD1wz5KL8
utnQ5sq86J4PBcXyMs7MzEzm6Ey7G1OqEPYq6la7tE4GwlOYCy8uA54m7oEmGzTIP+JrecobOdaC
4rbQxzeytYE/T1L9s0jjQmtFRo+TxG0Z9okGslceOkUST4Zgs84IGpz3ih5pna+23AL860ozxGRl
xwwYTFiZtJQtP4BXRHGvXwIDuMy/uvQHU6T+nPsxHsYLijVxOeXquPUCxJrdrIoDmmLF0uUJ7fs/
Fnm+3DCQ5pH7lgPYxff/ROfhZG8SEik1fC724SvenmonPscwY+CDomHfy0TYGMzcRD9WOeBm8BKp
UOQPe6MFzPTKLHwlS/h8+5BLepjG1bXTWi6atX8/XIxqJpBnalYifXhtcFDbuTLWF4EyFdjGiogr
hC3zH8Hu4A3Ke5CJgvzwo8uhFnGsBFZij5Ppg0nrrR2YIJAqaFLvQU8XNgWAm67U3SWk/9Ph7lKa
r+0m1GbQwmwt6QlHkzkLu6NF58IAMEx+1PMs0JjvLDQXjY55XUVLY4HSojxvsCrRsJmdVpOz0KqF
pfkOjLelAcFItN32wFcoXXYqSNS9xJIAjkUPPCGuOGP7RSelpMgHigwfqoO73kRjSxD0HlOQ9JZ+
6i1js1Cvov2mSCV2qi2wfEMqsPFvy2UrOyr7+eaqT9dAV8B0teqvawUY0c2r6tWm9rUcbk0OcrZB
Ezo5Zh0b0bVDYOBySePkQu0isG5EL2EOiI/1Joq+3TKAy4lCptymIzGM6LTMnFoXnYnxloB7NLzZ
psZrLzccUo6EbziV5EuiT43ZF3RW2zJMDpejreBkV+kKKfMYHejaGAFUeD53pLVuD9wRsflpFZnB
fb+/ZwzYqPiVStD0Mnq4G9DEGLRv5eGWZ7ov3d1yhwKK87uXFymu3UHKtMB1aUskKzJ41Z+ZUuTz
2EVYp6ayQ0rUNA2Th5I45aULnRTiFWMZNEOiB2R6B/V/YfVQ6Atg1stgSrr8RQPPZvZDZ4WQ3LYf
qBElbT2CozxJ26he6XmcOPD4y8V7HQoRpIumiLQ4RMOzWveE4ycvxvTfmhQPUlKRgwL1Ng2lPs+/
WOJcmEK6DJKusXGRRfex/VFy8iUfEarALvAdb9dgXGHeTSBy5P+lS+ptA4sLX8LX4tXZZ2DR5jH3
8DV8iGOBYiK03dLej4GYRKql5azbeI457tw9nLXeQNhK4guRZ99cdQ5LzFcxtGlj1FVLyp9pEcRo
2m9aWRMfm9yN+J+Vgzz8LvCKoHFMxSz9LoNRtfakp2iJDoaW3BTw9tDLcTqWFiQK3wPrC/NvUPDF
BWc9RMJSAoPbWXFl1dXkDonRDDK1rR3+9OXyuj04Px9oMKMxhuCRTx+jJ5xIxFa+wJdAsR37mWZ2
xnR/WyrrWwsWn1zFttyTUaVDyll91ri0VzkQQ4+BUniYVGohYbZ4z9j8AqpsTzpwS+tBg1RzfGqT
CkfYqH5zq/4Bop3Nmx3zR5zs7eMWfyonLdMKCFo37/fw36KoKwF1COhwbaybpTb/sJQQry2TXndu
JD73ni6cEzm/9LbckbdVLM4gM7oiVG7nNO8QBfbRsp74VhIA/CpxXqzzEO3m7816o5GxYERXl3ei
Q+r0XYDKjUDi28Srad/tW/CuvE806ifflF/f0H9h1N+LQUMiZUU+TrpN5vfNJQNU1LJnhM8z5Vps
WqOZxM5q1zrQT2zfdCxsHInYFnQLCPaDdC4Vq8JoldyvtrfsE3zO0GGoUZqxsp4y9XPYPDxtOa/6
AaqRuECXWbMd82zaAz7iu274hog7viagD9xw0T3sU3p80ePsL/vZ+gCBM09LrDP2GsYnvPSQdBYc
c1uK/omRPFIhkAsFGe1qayYU4UT7wqnqaeNzq1No9/vUDh8J5nLzB7YQuFE10erB2eP3IBbikOp6
pRp0rZDmbqcPCPKg9p3+nfF5++6FPZXZUDchV0g+XyUjm7ejpuclMNjjmoiBgsjAxaqlq1pV9ICr
/e/rVJsnOH88ZwPGhkip70NTPRxefMIwhdYKEiAjIAE7Ktj5ogGn8192PqzAvhHKrLiw1M14x89Y
MopGwyQHvtAmYKX4emIyMjIPvqUBU9WCELEmcdkDvRZuYLDMLB9x8MYYHRTku4MNew9jXNRJJBsB
vsAh/45Ba7+oxir/98nkzrr51DrUKNvgasEtmw2ZXHHd4YwfyE+/JRLgMdGrTBs4TMo62b/aawYg
SjBnDRi/NCoJxyZeAotFDtXxo8Qyql9Q7n1gEgr9sqb0ZuyMy7GsR2nF9woJsfXTid1cVeA3i2CE
JOMWqHL4WwJxxtqKCLC59EmD3YLqEmlafY/W4i1KBfEQbyebLVi5/nZ1GSclzloWSyXkAQ63Lo12
l3aVJ6PeByQZwKfAdFhD6QBgc8BZKnJBSAiWff7uMokSq+hLXY3nst4769VxNNY1Xcb4YvcwgpKo
HvnEvUvdoULwH2GEaXlIvJJ+TKHov/c0sQJFbog8JCfZJCplT/8RcbaFNCktJId6RkFHGenqU4U9
1Nk1qpM8WWth82dIjyatiDJbCpLmYGZXAa1Daxfc0iiuzXd1FiExhons0pQbzvkMUkAOenFkgW2z
8vbjXqdcBwL/U+AA876dRJ4qL+5KQ+P30TBb1EnMPYrdmuy+bXVS4RizrC39xdY5Sc53r6fJEQU3
WOenFNhUT7bIjcW6KPgDI1GPCBRwqAyR81LisGuS5tLj8fo/VqdJ73sSmrPyQl3WpxtVEolvtI+o
7UWHmtXkPI2s8mpIvN0Lb+po0QA0sr26UY8JjdqyIDiXj9pDWEFRnRfvETR9Z5fuxu7vpLItF/qB
6P5r0tVFUejGhlGnVksAMU09wyh/jgDPiEFbY7Ve6XFaOwl1RCOY19n7mpXgLNm7X/hObf3B2Xm1
9RWbpeuZkdnedDNltB7yyMTSA5pnwpKaonhbKyo6dPBMoc9YTzLAvAbvj0udZTOPG53s3/clhz6m
5S137sg4Aj544t5WP213IrHkkjcl5dTdrWFtIkxuqZjlzzHozBHMgAGFeJ4MRnJ2uYllvQMIDgfI
wakSyINmqCw4UyuFEJUVW1a+Rrr+Xv3L69o8w0FfDhO6e4AkVejt3uBQitpFyko2WKY/vVmfzjRK
YTzlEh05RrLSAO2kVy8P+e83f4xY/vxzmf3ogPehJeJ1nl0LQQ5bOEHZfcWYRbyRwPnD+L5fb8Jw
FJR9oUrggCb28EEl0i/IhvMAP3N5t2k0IlBKkX/4TLNAN+Bj0gN/rWpafg/UuwG+GrO8a9MyICIh
NSL3ZVGHDW1/HoXkGNcKzpS/dVyZlOOAQAGxOKw2UvjwcPaZf+LYXUboPtcWwxg2c4WKXIotA9Vb
0myG4ClzLpLYGAGOUc4tofkaEv4EyBoceJ3FklxF/2eF9Y8x6ku3hzGDNfCTtCuvsitRJqfWKlgJ
7gPq7P3bjvq9RElArl885l4qbkzmHz6oByZNVV7XHU2LrTLSvmg/TEod8dV0uwnp2qKHvkXC9nHE
EVrQNBIcEjmV3efum77awB51QuzBX+9o+aZ7ZAmvwJPtqaVPSy1/3NPfplItLKrd87yPfiDIp1FH
sdZt2+bZ+he3D/BzR/CovE7VsAYzFLYZUX79PrURqXvfSkFj8kn5H3OcBeEQ0QoUhe2sOP2WlEGd
v5gLzlMGb7/YDc3Eb1P6J5hQyFC/zQJP1uvPLHIFTD2hqNRGDfmMPQPTP44DwqMQdOtMzSL+D4V0
eWMr8t1kJnmd/mgrk2Kd3VIqDeIOHkeeXfRS02WslLLNslGDH38NJ/Ve2o7KmOQqa/nWEy9hC2of
FMKF5vWNxVMPwPAJLHBqw0AO4pAOiS/jRoOzcwuKPPSsVYEsGfmprg+uzIA+CumminxC2PDict8m
Emlsk9XCix3fVwURvWq+GyJ/2fumUJGrhb7F8eRctRBGryShuDiy1bTEb3SPw7/OT7WLbFC9pEdB
xO+6DJ/q3LJXegRkaevux46RIikvO45bEFmWRt75kLquYOCRzw2Cb18v9YzEtR9Eq3WoTDSEd7Gm
kmuXrApdaz6Ib0fQfqBKbzE21+hAWdAwgtp7X2Sfc5/wpKElPlPe39PAa1nds92nCfTbz18TP6jE
DYv3JgneiXz3wMoImiKKVihiAe3akmhyb2FIZr3W5RjhM2Q6xdWhygUwQrSkGur8YwB7idlPIyDU
Wm6aQ/Cw9QcnxkS4QkdWfmCzNe8E6s1y9STeMfDWkBX9vVTp4ReU517hHJ1qiFTosbzbe8wdeh2I
EkjSxXMnvF6eAs0JrJS6xaBZ3qwj4ajyuBCd4Yp9+zBeEzUFfBSj1aY5xFs5AZy1Y9d6UC3VdyOS
VnCt6ArDORoGauAiFce3LwtAGmTc4gbFN+BHTwkerO69Gny43zt8IghshHuUVmw51p7N1/RPTYtG
kl4QiP3tQMHKV/gPky+5ykiy4sjcOxNPAOCaZAZXWe5PqURdR6T5+cPgjokewEy38uYiwofiREqE
+X4oh2A/5CKwp9sE8utqjZHAzxmRXuJMd0oDoynn5twHNQiGOUppOkJYkDdv4cAA7uN1fXw2d6bQ
RlP/O/DSyZZKK4459FLdMChUU+gZPRrU7TEIKgbXnqAn8MKVAUEznjmLni/fSX0ZKKtnQMUCbTIA
Kjvp3RiJMp2DEPg3NxL/qvxDDkju2zTyIwfdiGukU3gECiWG/2Q5TM3bdb1Nt9bAYf2JGLWkPEVB
sbwK/pEMwzzUdWd6Koa+SC0s6tMZ23Yi/49mM3TYOeuN/CA3vVoyR8HJuIt6/1Ti4otxkpN7pzYp
4fvb0oOG/BYHpZRueMgTwrfFyBx7+48GYU5b6RXjA3jyv1dfrLJDdMKnn0yX9ag33MpXCzOL4aCT
O0VbqzJ5SuczcG8kgniqNE6wncQn5y/l6MhG9ktuN1WuXPZXFHDkgxFyKZW0DISrT9OnabbcGww6
Dvc2HdNPZ4ckU+NHjAEx+0iNpzpuyO+j8WuJ643UlxdgWv4anrJ4BxZBAGPigcrTpUzLET955cxB
x6imgChs/KA5VdTvq1uvS0o0gxlyJXlKmLE4CNCVx4CAtjn7IFwsmgi2Z7r0i4/FN9HY1eN7ay2M
T78pwMqc9azUx8Cq1l+b4WcQ4EKfziIXUyQ7OOClqsHMcXn+KY9gk5ZO2iFRGyqRyxO2xvcQl3fK
x21takVZXiWmN5hLyWA8BhJkrbqWPVWVFKj+ptFOSH5pORhKh2/TjmF72zyXjGk/Qt/TLa6oAPB1
KW82bBqrhyBg3N17lSkBYYbnVw48IeXbaVEdcHq+EK3Ax6VUcEgNp2KmhE7GsUnbt44KWUq01D6u
ZXTcgNASNuimSo2JZWdLmtXvJQiV5dVIiRVFHHvG/6zs7Ag5CueVd4wMjmvhDu/IF22/8VIPur+b
L5DSVgisirj/z+/aIrs5hygjvU0JAdnwXHCGG+421k4nk1bhTomjzvMrtkhtTK/eZ+5bliAhlEr3
2sha3qUfNXkZE+EnkqmgJXt+45l19uQ7JlRLgyRrgoHsdvZtgiRGQBpH60UwWqeUgyb7o/0wguEG
axp/9xC83YJ7x3N/RgFwVbC6gjRZ7GKOWNVEr1uB7V2KMUmwMf6UxWU6wVqKLhbHsmShHsnGJ9d4
dp1KD0FE5zFqD9aXDzgCHMSReIcPoQP/TAidv1+MN95ASR2RegeLCNIS/ZMyQfl2hEnqNTEfOd8/
KG9FhoA4p/z4kD2UAtwxuJY88W5w0d19G+2Y8FRJ1vFs4w7w2MfLjSqTE2D50FVYY0/ur2wbxUae
odUUlATOEbVkQwRYV16HqqaVojX6g5uOy7EJD5TfnMtLvHGNIILCAb4rgk6m9mC0nofA/eB1rxRH
CjVSUDquUaVk1RKOz5G03TBpP4FPfDcLEfzo3PUBM27yZs0ScFWEulIfyJfJcH3oJ3c93qVUDG0T
3Y3PAdDOzOLj/sGmB/lTz4dixMPcD9iAVMkRN+P7SMH4uqvY1y3/h2OUmC/446M0ab4AOEgbo/JE
27XYYdb+d4wKTjkWpyeLLR2oOvUfbt8lAmd7iZiB2jsWaaWJclEsEz2tcSaMEW7CcQScWrzGoG/J
QQkcyEsNR7j5um/CseKM9WXOW04mEbzkrTfUHCK74BpfGP/3qadafs4jkWk+qJS9Q4aDygXojpuZ
q5x64dgFP+Ukg19/ZQbXG4PzVwtVKmpR0s1YE+0wsoezbW3A6msovM1bxQthm/CCcUGIbphZimIH
bIJHIYJUw0WWRvLWpIhBLL3hVP8/fAvoD4Zz6ua54hmsMEw0YZI9A6qsBMW7kb0iaJ8YIAAcmfY3
Svg7MsxbgbZeDZSJDN3TlWg3n7VVJBBQDmZJbmiFoHL1wtgPFB24X3v3b9SWEE02hPWH77/ek/JJ
p7wwx13zZjIJqvFzBunpwaymO6krHwOolt+ndSQmUhjydUq9m5TAbx7EhArC69jz64Zk5bnIrBQQ
+Mch8sLb1M6P6IxjHPe8r/F6IF1PrXj5IlHHh7NjqlsftNefNCFr5kJZ6+kph6ySV2TqTfMrUPmH
XOvrmgZFZeEL8wUwP8oTmB23ZUcMLORcgimivekIq8aG4RPc24wBZvnPZosr9JLyy87e8g3HZbFd
t21gkF5i3Jm5R2KCZTn+xypk1GXWanXz0raxnHbgvZ6uDie0LoFGdDO/6/GjhFVTVxAZwOeP73uF
EapR6xf2ojGptpLfgFrvAS7EwHsr2vTlLKgrfmtgyP4WI/zl0XPObsywSAm1kFQuH5zgSY6pwhDX
VnjTLeJ8OmNm9WTLsSbro3eWDYiyCukLv4ppZ71KaZpIaDmIzkbKgHj7iV2RAY/frSg2AmboU+vc
+jBAnBlU0AhsQkohMzx59gLw9SXjAzJ9DoAzmkz1tD8T7Jj0h9YvcBDz2dE1mEAOB/K6abE6FUIn
gKf6wTzzhZHsTiFJ/E10z49QvC0a+UCmgbfy2fW8cqoTT9HBKc8e0RjFd0L1a3AwLAjOyGEc3mob
xK8qWWRlEEQOlSsiAlqgPycZsTAtysFeGGsdoLEclUOMYKYMk4XmKq66i05OzCDi2BfZC267AOCO
Z2kbNq8sgAaaYg6xXN24YCGz3/UrwaLeEB/i90UHjlpABT/I0coSkiT5L1ccPMzKAkXqoxaUbZfo
Mk9bvNGvPNe8wpwPTEkyHOU8wEfUzsnrdv9ZsPKAz7VMJ0E7MtLfehhyX+3FQaIgTOBJ097eMSez
LcJzaSatZwQMSTt4k630Y91iOkTR/T4qSfDU5MRrQRLj2jKBJQGKfiIQ6Li1Ulq5xljdIMo4JBaF
3jwx/KWONGQ7HxLjD7xacCT5fi4v+0SCuCtp/0no5NaTsriCJgH6XE1SXpXsrs9FMyaIWndmwZ4t
bRBMOC+WIiEGFdIGK4kbVm4c6HUw1XSh+J4Vc/wj/AtRYafZfHMIKi7OKsfiu33puRcOpSqM6iHP
zAJMZumRRpp7RIujQBipDfDNlmWMAzZrxZXNPhIYEPhZ5kUMBEZG+rw7utEgHlffZd5yssJD9wdy
krh+gD/741GDENRo9VQsNn3ohKJtcJ/FqcLz3tuIaNUwghcIhPcOvgs0lrFLQ+EKcUXvESVmSbCi
9MLGpxZOGk2ATrLhpXCglky1/jj7/ZL9fLhp0COwHmnzp+apwwktyuAP3mGDzkTwZ0LstqtmUVsR
QmthkkEH0v9OXcsp8f3cp4MuiI9MldBvJQy98B5zIhpk+6m0lAhki3jZemjxhFR20Fnz/ZV/cZ2Y
xmbnHIKkUzcTNZsa8nYzB/i/Njjol9cc230NRNTdIkBegJYy66uedB+inRREsh0zMh8jvkHFHnw2
cpDpG4Ofduv8U25/J9+Oz+V97EIBd7/KnwQCFLTLuYyHbgPB/+26lWREAswpXElWXAHoxjZ3QKKt
K951qSIZTVPkhqBZAsUjS+4OLoVIMjgigGnCQOweo+SHnVzztGP1aZoWmREfKw4jb1fPvCaWvawf
lkWnQwT2zCrH1MZHoww2E3DxwNowm1yDgYo8mnZl70aNu/1THv6S6RxUh6eetGRvY5x12SlSICoR
WsNggbm5AQXokautOg+GacVvrsHlUEA+lVKI2VGeITLSKTrNhGXlDmta3pvcdXEgdhFxHxEQF6B1
oRaE/+VLFpr1MxPpnGkZf7/6UcQTIHJDpQ0eoRR25Ql1MSCc1cigWgXiRioptcYlTwaiHPcLNfkl
pxg7kdLlH6CQwF8HvJdK8Bc2BMiN92NZoihaYM+t2bvMYOg3Vjyu6HIs5HrQERfJyTcI15vWvrzM
SMJUmAjJpcq6vy5Y36ZeVoelDt5D1dxIKqc1zLeIBm8U2/lcZFSbKAHe0p1IkgHoPxirVaxqqefa
2vGZRESW0UdjbUIw3+3+pnpVNsyu8KiwwRgfISP3BzDIW6X1mFuVR50m3Hkdq0xghAZG+mKLyNY5
VNh4S3OeKhKDnWfIcTUtpM1ro4keTLTA12NvTjV90aUbNxCXl0z/VjJzKMLKiis/I3o8UFehgAhl
Hpti69pQR/sMBI3R2KnogpX/XFna3NlACCjWwlAb68d6UnWThyRK4nw9OjNxsqWPSBZYc9lkkk5N
JhQik1hT1ka2Zxxajl/zo8BlRYkBluq0av9yqhM5i16dgq+zvD5BaewcMVQHcUFV6ISif898npMF
j9mgRO9t9xsj6KxzA0pEGVR9aV28xMOj4KBavwYxhLDv0UrUZIEJAxIA4ocoKWuZrNRwElUUvZs0
WBeAaM5Dkkf2SRLQnYugkmZBmzxFA+z+eRpcZ4CdRGzqSJ8EBKSng6/fWPgDmeDrbkTeqZFOOR8l
FHOzTp3S34UPJAYeG01DsY0oOwQtzAByROEBBOq4bgtWIu6o6e4Hums4zBoleuXjiVhyMvJ79Uc7
QgnApIiSqV1tir5HBq5zy1Aj09/bb/EDk8VUWCGDRFm+pa0tMvaYJUHGRV1jHtGdBPQpBA31t6Ed
eev7QBdY1fcvY47Dyxygu0BnWj6dIGwilxKuwQFllA+26X/4vIJi+Jb32wBM/U2L9qFkgu5JufnW
+UyMTKT3J5ZbJGm/pE5F6aHPb2fI2JtnTN37uwWizaaxrqu5wzrfS2zzPg6o7gqcm2/iW58y/nQ7
FfHWYUWLDP2NyG9+dXv/Bza/YmCiTS7Y5dvF65qWbc0MyvY1tLl/8TlA3ehnMJeUZHXznojCi1Vu
Jyou2ET9Jn9kHzR2C1xU4n6EBkQ+XxbYx8Cnh0pGFSQTs/xpxuRgZt51eF+OFewmrlKsOiEPBQka
5vGIaPKgp+WqUZOJFfuLr0KxP3UuvXKpX9Zq77cMgFb3oA40D8oKXxTDmmPWy3uQLlpN04eWr9tl
yDAhGYbm+JdruwMWdBPRv8RyVQJPCBqgOs5DIjm4vHwtY8eflsJe/5QMZON0EhXJPMq8EQ1w2riu
qQ6Z5H5mj+gEIgxlb4sEOh6D3qXC0HSfcpdPeVlHOTDRLjK9jz3QgW2Kwz3Pzo8wqbNvTnO+2dZg
tAdrA75tSA9i1eShcIwnPjm41uyV3Go05keApHRfpPbvTFs3cLMzb4HpGBz2x9lrtNoWPtgLEui7
ttJmaVdVfsPPCBH61i+G1YaV4WvedV852MqVdGvE4gMN7mjdA/0cHcqy2KLT5sSHpRpHFj6xsjK5
oUcOmVJDByS+Is7C8muEdSgVs4pg4lnXWvSMjlfy6BUbGmvx7TmGlMWCgwZeAs/PvDHdRh6SHf/7
7MIlwOQ8tkxWVg0vgJl8gZT4O0sPoggdtBxCQLrh4YxKoT5BNPbdhcVpvvOHVO5CX6LDHZdRoOrc
dEeiogA1WzKpotpjQSH/cbjqMPvZwt8RCh0inJpvq/r+f4csNLT6D5glHpFE7ihBP8vWlOhJWaMO
w9aXISb8yslsRYRTzUkzyrzN/7XqwRQLfUFVD00sCbnoluo7wTzFUugHwRhbe56uPcmbjxP8KuLy
cvL0AZQf9dMrj90hVTmRrasJDyW002UUVII27aK1pT1FAI5GWN1iNgFJVrZvfN8CGhN/MMMKjHf4
2CK7wct09wnMHRYzO2vQl1MOogM6E9yDtcV7f/tsnx8VH4C0MPVQv3rWRHgYKlUJgL78fngz/rbi
U+7SEZxT1U+WgbOYmZxInVV7uK0OlwIlw8Z9QGn29muhWWE4svDVPAZoYA/3PmmjnKlhpFoKuzWt
lu5a0z60U163JWzQjtjAt9pm+uU5wdSI4cujjfH0D2iVle09JAJ+Ap23viJ+FQwF5WVZfEQKcACL
1Pp9nxNlkzoemDSqW/mREL9+EPYeUafHo3x4zEryADAY8K4QSfPFvtjTnp0Ni2/GOPMVOlexoA8B
c4Tmwkts6hXcIdbWqAT5yoGyU3IfJ94G3JChqRcrrztF3UzlkOZcYuUvkvyizGRdQxl0mw28azXY
xSJqP4UqpDUhfWuQPKZ4sCeeXRj/gt8lE1fC+ul1ud3zqb4N5uBFBJTyEkoAkfvimeFgBDiEJdq1
pRr1pli8q7MslEAEcwWAqYbhAqXJx2u52pnWIGpUpTMkz07UwAgtsDu6itbAYfsT3b+WvHu1gD/c
C4mWswSgtzuyQPTuOe8TTxs6KXeb1P83aoOd4ALkVzUYa0NtWLI+oHBAFeSmNWUCWaA8r8a6znsV
2sRDTNCdAcXnmK4F/SXDn/dGSp+Z88fPE1GxFR6l/n6SW+isv/fNK+jEVJ0bYD4Obpe/mbLEJE9b
LhLCjEO3VDVtVFXzqHJb71Myn/Y0oWQ4hl/pAGHUJBbMYvKEzCTaw4guel7fz2alSZOWQiaoVFOA
9IxyuKiHUH6wKTAg3SqU2dFygVa2FDOGFP43aXevxjM6TAqsBAKr8w0Xy1tIah2SboBs9E2DpcJ1
70YBzg4ClVUiBqfna7wTlLSAMrbVMVoqE/7i3FtWIzBNK1PTcIdt5y8ONaqGBnlAKOpMhIRNoLEe
tSSkTUHhkS66DYMqrgWbrZY+rEhh5ewXAOh1jdDzKS90VaVKUK4C2K+0fDwjAYbiO5yfQlYtiJp9
4uezlOYQC3nqLklK/kjpOXollWfMDQo0BO4by9DfYjeWQHfoWX/YgfHF23h1kNuZwcmySwja5vzR
xhVYJ8K0jziMJ4JRyvDEnif1nfIbBs2tHLCJeYaFKaM0Tli4k10bwOgylTr2HkcnUTaKfIbkRALy
gq/YC7pXlkPBOg6PoG1fl4uB5wAx4AArfWgZyQhMbNOiJQSy+zn9f80osenEATDgMdpLjnS9ZtWm
ECzwy/mWdxuVrA5JdU2dxEFzBWdtJsos7xTN+W4/+UZcQJqLmJ3gyRf44aGWJpU1/L/59IPAMk8G
dD0WVkbua2HdmJeCAK6KWF6mwUlH07lBo+DA2Ps5KEaIrasQefglEdFDpcR2534+ffzKYc8cXyud
tIhCOFIuh3q0QZOczbQ8g0HGYhXPM5LkEfvgcjB1DljBsRxkr2hBDmvHpV6v37gGInXZtEmw03T+
6pr6Fu/pitQVJfCMWzKgnmcP5tI67GnyKan4kkSzon2VNzzzUaUuCKhULxmEeEE5XXC1qF0XV+iJ
qASVptRx6l2ZBn6QjEfLCi6mj2AFDDrTR6wq4A2NPeWiZLeWKxjlSn+CVrts8vPzoXT02f8dmBH6
7xmpc3ElPW3cLeypO07oFpiyMVBAI9cJZecBUdRRPTKAIYQhV4n2WaL/AGmgLpf5uemK9o8L6g33
kQYoU/jWm1a+4vb2cM+/8XFTM9z39yI/+Kz+pgimYBrxUTUh2HaQgBsjZxT35yk1nAHpJpHs4MMY
mHTfRm8gUGxjVr0oRlaNkc3u88PK3Bldc7ZebQMzvPbdARpX0NuUsFwWMTO/vJwfaEvXzc0gO+6l
jgEM9//eKyWdSJBjj5HdLXh8ZsoRQIjIq7yYf9sGTMP1kgT502XBXlMNs3CbLUx43FiPOdos/Azd
qdqEEBOp/8zYOq1ntSjrzuU2i5URWo+drry+vKtiH8C3R/ODs4e1dhpHOEh3s6Osm+oOrLB2r/OZ
tvl/L2YUJi6+ZuFuHaZlLuMD2IOp1pNAo9zmZrOmQVzL2lSBI5tCe3E1jPeme8x3FuTE/APtr8zm
3YpA4xaOEjcAgt1jjWxe4Tdn4BfzLkv4O2OJxObUbjWiu3AM4vH5AaZwlCdnonDfA9RZvO3hSpCT
IQJJmGVlKah6CcgWvC7AFck9TDbWSW1rRIE6LUXbnheRo9v0qm6lWcYz/dOhqDdJ4+TI729aUyw1
hgaVOQKUXi7YS0wwkmxjEIpbgYcUopGHVUtqgFKWvdG7Ef2QwcysmlIzHk/nPlnzU4r+3jyW++xt
0hcsqtu2/fqME4hIAo1D9N8LRhvElthlaQZp07L/Rr/7Ei6oRCuUCNAr37IBMswFT5mCFDOWTdJ3
x1Lma054GEWSewqCHlXX4AADcQ90lIUGCtlq01SgmQam0O11N9SCN+sjGTKnRSxut+eYaZe4gSQn
1TICHUA8aK5tm1UaorqFI/9DrejzvUpef6pM0lLdQMNuSsSprHg/L3L//WK5xMnBhGJgDoL79gb0
4gQXnuCzNk4LqHmFDkC7Zdya5NaByiZZUc+wlsLrk6Q62V+bHqNL/67zGH2s8A2yWF+6TWKrzTT8
q/68lmQs0s7kt6QUJZL2PynGDvMjdFUhObp8igo8QOnqlE5NdyOHXA7vGm3OcvlMIRcTeRgV+RIT
rhSS1XlHZd7JuNz0bpgRT3tEbFfkjeP17qhYyZsS4ZSPYrDk1kW/HxDUP5Xs2Fnjuol3/B2AX8sQ
n3PoQiP+2A/ZKvPVwvMxOCT8I+sJMdgN35VDmskz7xUi1lHZtCRnD5a974nbrO/9H6J3F2t41P0+
4g2RK6U90rgPjtUT5ZEI7JZ2LWPBpbCgjYTD1CNjqsxSkVhpKITDZciaiVoq+RkTvbtYOgy9sMpQ
SzCwgKji0cRGh2c0yJ9xgtjXWPUF7vgLzOERy1OaaMrHdy3Vj/NfcXnFf1fa2Yux71aP7RUow95a
C42RlYkeK3ciudyaywBx9qMf2HaSy17Mmuhiy3AcSR08hFWwLyRizqJYDkS4I2WmcyMQexl+PBMV
mTOBJGS5Bmd9gl8l4HQH94MbgqqYRIZ8YdOM/0iqiWMUfrNMf1wz1nFCC5sqFzMDHpOJjSRZFD83
1f31ShxKAvQamOGg+I0EH8YMOgEOer1wUOhu18fne6r8wfH4uW08E8jSn9hz0oNRpJFf5Pvb6Yv+
uAWX3g0Vnt5q7OW4sCXbckfSegKgg8j0QfFqktmzHnTo/LTMysP9x/sDQzUxCDp0gbQWIVsIX7v7
geatWD4y5ltXkqEgqteq8I8mxOh4ADbVeM0wdOwK4KAakPqyK0IhIAn41txT6/tFDqwzu3iD5poS
Skik1L7L6+zNhbdGMSkgDSLkmJtn5qi/SUNFpqb2zvdtFvu97y3YC6EZIoYrCQpOVY9xeCfqJ4I+
Ufm5mQ2lbFe/5dcdJs/xaWp8Pb8biA97y39Up9vHiKOT2m5czCW1Bj/31rpSfuFSLhLumELqSaf5
HbCnUIKmNCEnixwJWR/fWA5qv4T4umx+sBtivhGupMuTQ7a10QF5GHSGePx/rjW8/QMt78G/QROX
XDn8TWMep/YRaBvLoXHr1m03Ns/6uAh58Nk0NcuGEzmqT3ROcvFhCFAOIFwEq5jepSBiMZeb2GxE
hdDllRFO/U5KKqhmCRqcGqK+ODWITvdIaUzFaMza6B5kqfxsy9ADVrn9VAfPMMJah1j0aIMGRhoi
iJDf4jNfSogB8oCAmTjoB/D1z2hiWgsctrK/VYErjN6MPfi7RYQ0xgbdFqvNLjvWpDcEUOGhB7nQ
wLcyUplUZlQJKDF/Ku22YXsy3XLxUsFbb7LUU7rF0hcgBXVeZCcA1XNzGc4BY7YYwNSOzM1IOA6V
ds/a1s5HhlvdscQX2EINvqIVbG44xCEyiHGLcyapSP6KWwSGaPWBW1zabOaaZcu+oGeSV2+3N2Tl
9fhG+EOcHadOJrmvsBBJoc1Gk9e+jgKQvWnCEDkark/2RV1zy1CogfQmb9rCEmM/YThNG/ZRQk7k
bMiCx2Bq081uejiwU4ovlckuxc9TV9lqg+KEWVe0gC8GlfO6029H2c58/Ft9ZXAHh7OsNI2vazGa
JeAZ2Du1k5w8VM8a+xudMXOkb58Y6EFIPnzGuv07dwjnLXBBomTxSZTSXR6aji1UkljKEylwgaga
1IPVZULfpKGmnyEhZfboVgyv6Sr3H6XOE5sJkiuOa/2XQ7DapOTpeV8bzBkjTKPeEOL9h3O6zrmh
JSOZuCTBRrR/E5kFC6H82JEEsRBBvLE/Z2QalZjxtH8CkF73d4jvKyvNrX8WbrhJkPfWuqmfbMs0
q5RAuM6qBFsPSajqV2NSEdEfSa6G4Un9RQxL/quYvYb4t4FR4EH+Y7A4bFkOEToBqXMtn7cHPTZ7
K+tGqyYGVa0/JHdfxfEeNSDOThGq6O3bMb95VKQXvSoMqY4yVPtbvsbgbAUUDZrMiEqj6KxmgPpq
BUvt6K+vyIW29M6HAaS85SEvayN9HHbCq5NaPbgc/MoLEZF266AOnXfEsLuJaowWaJ7hzdKNgKjI
bfwyBBVeOufNosA90/CmhqyqP8o2UdyG8CRxGnw2rS4QPd+SMubkoSWjkkIj01FsxPnm9nVVMVnB
9Pq4GaOtY6SzZFoNJX6jQCholw9Ghn7kBOrvDQCygkZKWUq48HfA9CncFcmJgUPHhXohOPzQWLjZ
x2ohyoXmbfe0OUJwhI+Xi1OHI6A5pqeU0bkiwR+wgNB9Gb2QW6yC8ofC9Jk95L7yjMP51nU2Z2jw
kcF9bukTOtVjLOaDYb9DWZj7ueWmue3/Rs7N/1ZjSUHw0NEtwYu1ywsUyMj0P5m7z90jww7YcyRG
Rn3wMdc1jOuSmRQ7LUoi8QsVEojj9vwFgCelcJsIwhSJmTFWUzbCYoXRrvTVnIuxAAU0yO1u0763
qbhRcvjhsOZvfkPTHRoDLuzzgUxKDEbWh1zc9QJ06jYQa1vPJ6PMv/4VQq5gK4ZolwhiJVjbrEfZ
zb2uSqMUdQH+6TEnqxTuuTgFnyORDRmeyFRqP/QJwMhPTIm/yk0FCX0o558bnHezlYuTjW8o2GmZ
MVPILags7rz8r4YuLO/xtuzNz1Ja60x3ezeW8OyClTaGiZaxeXBJOWazoO29p0vy4wWwLUgJrqxK
Wx/PpKM+B+vTpTL5DnG4xRgpgZZTGhSSuFABvCgxXFArjvdxMg2bd4YzupYFu4qL0STFF7GGttZp
Ra5fo1JFQo2zTp+luVaAfjzAF2bOa33zVQAIDkootQCXQUY/TvHxeUdXY/dgoNFoRy5xv+6RoTpv
7hPDdtu/2CzJ2hzGIsRT3bZ/JTwquqBBGEa7Cg8Qc7HA5m8bhnCZDQgQdcSfY030hWOfndsYVj9Z
KaV4RYHb0Ap2gNjUb048g6+WDT9sm0dymKO+t2oYw2PVrctngTKYXN54nEYjyuBJWesSc2y9YU73
WoGeQ01MgEi3ArSEvT+ez6vK5uI3Rsl8hLfF5Gve1i1AKVHEIPf1AKj2dbr5GmYNdwzBdkMdWB2z
nEkS3qUUOwtRyLBipxUgcgOI2yYRzNlUnXbyzbBYQ0TrmkADcD1KPx5IHzVdSp5nJWvJMDJbuSmO
vuOA3MhQeIj0isFznij9Bc0wH3j7G4GaIlg2jMS4LGwFbpcafyuX3e86i2WTei4k+Ij6EN+4xxOJ
XCGOqAKO/gSQ1+6lD8tuOAMjiPDRhHlWrPQt1QUIq359Uhht7TSLyJhVBMkwBJAx80WsfuxP+Lgi
dm3GIbxEza/U+NZVZX2OIWo2MPOmvgfGSEXRG1cdSgS1XFgYPf1CiUofFL/QPWxs3s43tvgdqtfF
0aqbCITmfeL5ZNnU2LScCm5Ny7kgashTIYyAFyk3CvqFfo7IC3Kq1wQFyZz18PV9AYuEqSAW0TUJ
Ij2Rxu8K/babO45yAIpHBI9BRy6GjeiUIZlQc/qEg0Hnknx5JqzzIQM0FWyN5hcE6fZjF3nAa7iL
c1pE+TOAcv6WnIl4jgqkHl4Tvl2mFYOdoDvGkmW2eHa0rdhKgGZbhVK4dcDIso8tclLYiVr9KY7C
QMiNNnJmmlnIF+LZxNmJR/WF4bnNiPRtniV0fD8JOicsyiYgFdwR9sNTz+ZmRgoNkJgIqMEALGjq
uTFf56Rm9Po6zdChfJoTrXltRVxuygXpj/bpxrB7ofiIDHsapAwwsYZr4+05Z+ZzM0otJz7lyKVK
dAZWeyYOMwAxipGpLyHOEGl+HM7hVEvE8nwtL/hTlSaDtSg42R1m4694l8d5ITzubPPtS38Lbz2L
QWwt3cU4K7F3ZgYX5sy55CFTUCTvu40SgpDGG1s88F4fhw6yMIIjnuEYZZ01/B7w5P3h+we/w+vH
udtkjfzSetss6qupdKWpzShJi43soakbj6mQS6YVZZ5qjKSDP+yA0veX/LNYfw5isLBlBW+rdNsP
70iDQ0gjsawCRFESD6Gc0I5GV2BRq4myHz0wv12rACbyLqNlgOcURkaEyY0OTX5e25IyJIofC1J/
7fvKVfsqhGQvau2EsuULRfr0SxAxjdATdB6JIdu9OI35sLnrG9Ki5CuYxRBTjEn/7beb8iZzDHoF
GdsmFJYkay333YOzl+/LXy6VlHvR05Hwz64SeffVGa4CIcEHzZ1nZERvqVyFepi9trk7SD/vzqng
4mXZ7vqTrpphbqMWqQnBqUyV/pEHyocHYfAc3Yq5T/Ev1oWJfMh7aWQERmpmh8Ls2x9fAxeTJGhn
ib58kCsuclRHrEj8kMN/GxVOUYGB8vwzvALhhfsJrhu5KQSDMLLxXjwcizxULBCguijZ3U3BbK0D
hwwbIapb+xfzLF0ejkmk8OZYPjVuryAPE8bkTR8kqwuyiuwwJKbsg+QdJN5xy3xpcCr81rXmX7OS
3ghewAman+q+noeEvcZesHEbw+qN4DmK35mLImVWoW/by5iBwUPhHkRUD0VjhxTL2pw9ENbB7BFv
vWbbMDZ2nkbYjh92W3c5lRdf9s+4WdaTV7XX5ppXxQook0ubU76Lxx5bvCp0+BTirB0ixGoogKt6
z0Coa8UDAo0QTfxKtFR8NyJ/AoIegLTVvU1L2UfYQWFIPtZLlM01BXOhsqYmcvnmyy8AqH+wZxap
krCxW0++lIxxu05r3NOozVt6z/agdO4cHHe7FMzoN7HDlepqpRJSeH233oaoQho0o2Iu4aCpbuDy
0JxVozexao9Ts2KvGj1HYSvROUZQWErjpGnj52/0ZwVJ7uF7WyaD+6vA9oT/mg9q9P5UZCTCTd5i
smCoQpzWOHCJY2Tc2ahC9MverbvyeC+PQi6ZC8k7f1LAriHWwqH2dS2Tq68lngd0t+tcjgdm93JY
FuNIKjkx3A6qfFyw++PWsJeasQ+Oz5blBp+0FZYoMi2UT3zmfZQOJkZy85jFCtNDa33nSrMUP7vN
oVw2E7pBN9hWbIaWUXnP87UUd8roINLjZaUPucV8JF6p2oZcCfUMgwFeFSBTjxdnJJC+LU+oHoq2
RF4UW94p/iy7bIV3YyW8C596ODztQYDqoiiKOI6HCS828nzazA2siOR62m4XXKiBx9HuQY3x6wyS
McYqOPZmx1X3TalwHVcDZEjmE1pKHlHMgyacgefhjROnl4uU6Xfph5g/jlg7ceJ3jjrA24QBjl18
Ys+VLB+FIXFbc26RGLdsC0sv7XWc0ZmzexIvTcGL5ccA992Wyv7WWU1bawbYsYp+TFiD/VLgINde
T4LvbJYPlORVlVzoMp1UclIjTbRRZEAwmrv2m+1uyQRTmDKRC6EtM/ouDcoomVxTmC5zXHqUq/Cd
bEgcqTp4fBKhHRRPmUWeBrWHuCsXdJ9mom6jQjqGhlFmLeNoEy+g9jFmL+/MC1EwWDZO2dBxnKes
2gVX/z0c8OQBIXCrBW7bwIjvGbq3Ihj5t8q1cVLqnRaLTrnISX1F5EcEzUj7FDNNd+MOCslq8AZj
7kcNRUOO21VA3RY27XuFB+7ZzkdGRl1uAtRDN/7C3un058qiQxry4QbnWB/nOv25i6O0lq9ikuRP
1mlh51h0X0vyzyUKCufwDJyj6ZR0WHeLvdiRwENoMN0iadT+OUm/6oer2WNlyFelT+7/B7L/0VSa
Rmn2VDCWtbsnYlxM1mAq1YYXBpWuBQtC1nmKeyuKd6uaKBF49z7sZOP1wu1SMhRLUud8fZ8CG6R3
H8G9l3hFljwq0gPvEFRBYzeHp/Yf/11D74P1sdTzApLhnptGm0KWYcBdppXmxoqKyuJH2w6w/wAX
AytmRT+OyLHQnHVOXiNbohWeZQr0GvQHWFKIVGVBjoVcNXBxhlwTRmSi2ZNSOvhnqtK6GnoMJ9Wg
UIHflgdk1aXDbEhtlMJjRCUUx5WwpJejw34P9AYtWeRqXvZH7iTtFPbBZhGGnQHBAdchnkPbUapN
cLwNIPdbueey0ZctWT2LCXiDZ+qJMxuxRctfrxkDZXrw2GtATPB7O9kECjJ+xzTzyswPTaSFnAu0
eElozcTD54GlmiJvhmK5NvsxJZVe8GxsCxZszTLxGYZDoNV/o404n16kKYsQ9WW01flPzMwl8I5g
8dRq2/WpV4SoOf2dlSKJsVKG7ghI8CfIfACMYW8CCT7bh3tP2rEUfmCG/gsatwPMMJ2+lLCQtSHf
DJKrpxWG3NvMrxtdQG1hKjnxTaI6/lBPXtUaDzzyfQDOYy8x9vhHFABy9gwq07m9BGMYJiL/yyCL
lRTJhGPUHixQCMia78/9FeSkrPN93Ds8EiO96dqH0giIn9+O+cB71f65VpXZo2h/dOKs4Q1JolDZ
++UGm8JFxp8LCl2jKoc9M2An2UsC0fY5HcluZeqI0E4GWt+WdtnCDjdz3BxlxwswSbws5IGxBLOA
1aoMSr9y6BY77p6SadW5/ZqUGT7mOnCikCy5egNMaUpJRgoF6KrX1Xvpnr/BLAewuZHmawhVfjyQ
DExvO3GMORlENLhiMT+bUsy8VboT7eGDpZ79+9MFpMXTrIJjJWYCe6HF4lGwpgnygT4nuhd/JOWy
IzegGo/0UKZENA5rKvEvbFtzsbVV/817KhijDqmdURhJxh6vnqPOdwg6lKKZkkfBSCVJviZ0qqqY
KJZxX3gwsAnAU7yIp/LzZb2t3Rmu3/7f8i8bxqJajdMBgnGegs/YyCXro/j7TR7+fUEuGqX3YEea
MpfDuoY7pMxwcL6zBpLqCDiUXSE0M9OnOzSS5Lr2X0Vp4hXKNMYd5G3wjQutRrVU9uVV0Q8bAxUx
lr1wMBQEemcbnybAFkt0diAiHx31kM8pIK6in3pYXCt+qpEQxGG0vQuu6VizKyVC3+xKHyubR63R
o0IXimqbSIUt67Jpw1YAF3otBJMLHLTJo7WWF1CZ6PIOTcI/oJ/qBEGu3KWjxxKX52H+LJ5iGIQl
7cbcPq30/0snZWayHpuZwOdf+dLo9l5u6cGrpxRnkahoy9arbJzDrsi2dvH/fVbE9lsFvhbJn+fS
sJUPIqnXcobsNHeUmiCdMR+C348PKDUlQCeSy3ss8lYMD6bidKwZC1xdXyWw/qRBAeZYJsoqnWgF
hW5N+vZ0LDrTLyqQGSA3meKQ9+JLNx7VhlIioRbGcdTuzFXCoGU7KLy4lceusN5LrXv7X2kIrInB
N24NXZJyuSSOBN0X81vshjJEQyRGzpmXpruDQYrey4vQrM8Mi2MEC1O/Pjp/NaH/rn/tiVOHQieY
Gh1BOYoHFHK52Xae/plID2RLcAZZQJg8NWglT2NFWANSlDBhaRta+2oFBFp0j/dFJnQ/4NZrt3Iq
G6PDZGh0iAag/s0y3uwd6EdCv0XOdTV9W6WMpSxP62FFK+rkhA1ACL/4NJoN4feVenw0R93t+Iye
SXG5vLTJ0XMZuQMxP129rfw5JDpLmE4X7IL1grETVFPYlmL3U2UBTyPddRui5de4/LxyKnse6U2F
D28pYdwzZadjQttX2tfcG05ISXUF1oMC2vIU8a6qR6PztYPRWaBAVUwi9m6fUSv+SyTh5tR/PT6y
3Qd+E5tnblxh9qjR6Fzg8F+JQZwZQk2eBOcGeQFJ7RTFkouOCoh5MnBGTsIAi7o75H62dmtXmewY
RBOTd+Ub19Iyx6Q8cynO8W6fPWuoSPc4gqbaPc7zE+nYEmCxUvOX/55UzO2LVOHJJ7stu3U+Yki9
hJYsaomYvGu42iUhNkH9Ur28i+g3MRsveVzq8ndC5M0z0yxJOXn8VeiFrvsS5eeP1fGebyM1i3J/
89yAyZXOM35MED6juWCm0tZYhpm55o5Z4RbknHlXAAI7J2CwtI2zd9YfQFtDCGk3LirRI0kRRz34
ucnWEqhd5mKp2t+H3oEhqlQKbSihF8nzKUNHrU87iGBps/NhipFtDecAAyorytvo9HyhUbo2VoYq
weMM4InuxeR21OCJ4UkwUgDPjLASDrrYpBfg90B9nv4z9RVReH3M7zelrWvuAlc9fSCQbaIJq/Tn
1yhIOEv4iEfA/54e6z6g25yBPAKxLtsWIIkjFGci+x4lnoDqFXsz1kZP1kyZaAGmuJY1oFeTpBzn
uF0+E4a8HyGG27/4s4OENZGx/H8iSBQDxWMsWkdK0bYFNCsR8gj+qbE7gx7684vwfFaGyjadV/lA
JKL9YMBzRCj+zAtPqZEyTyo7CXmsUv3v4092C5XTsOv0KOHZ0FfeYiiPNokJqZDm0HE7Ht+7ragr
EITYZS7w38dsplmBCkRriN9JmPege7ikM/bbpvQGjSDzuBhKS3tuzHRSOpDUAd9nOrbNeTWVuHDY
Rrwa/CL5taW+mcjhhhuAE4aiaBnMU1lDOj2U+RB+7IkWkbefIb9YiNVIuUcTy5tV2fExOgUc6N8m
O0ymtx69kx/bx+nyBpF8uZ+7L2RnGBfu2NT52Tz2dB7NG8HwuFgHc5bJlhg2/hwrk4cOY4lmdlb7
N1KAPOCQB9xuLs64Cjr7B1rgP8WOz5t6pIeDZiPXFFMwauNZS06XUf6+NOopcxKOp6bKPrbj6TvS
BEyC3I9IzYAqjBjmbqzL4MEBMwyqHrlbI6jOgN9bT6TUwv29RyegwSByQg0J2xeYI3coWwMIy6aJ
ov5hOb14u31+TpdsKJxO4xP+e6LWsSNEedtLLRDwF6mYsJVnthmGYvF6aja1qPREtbZjmXGB6YC6
qQh/wVZbJqUFp1fhY9M4uGBfIW6kwNGDCdXCH5sAub9V678DxpY0Q+Iwxuu7V/EW4wXxPII+W3ey
Z6a7iTf+oD6u2zsI9NdqdB7u/3N3tsDZIsNVzrP1CYrKi/Vrt6Dvyh3L1+1OGvfc+dIEu7s2JLcy
hYYBS+1CAf/+y1Rfp7GAwcGxDIMY9eo3oAjaHksJmPMVJk82CiPFnvFZfytljga1CzI+Qfn0Safo
ztDhrXm7iO4AG/1gKglNK7x4AKSNZh1fobgXyScA0/XX77ung14XhkqSZplMneXdeIfFHaxf/rY5
7F9O9hdVtyIN/CszLq83CSqLavEYawSpiEcI0uZazwbUy3wW320XowOGXMcXRgbCapzfAr46ACO8
d2Fv4kZnAvxXycal13jOLIxPaBVakTvb9KmS0sVha3LjLcpM3BazgmrspFftRgqGpijXgeC4WKpn
KUE0RoivxuFyrihiU33g2A4A04eMprMjGlnVv29rMITnQ1urhlOc9R7+NmXKOUHleVCCa/3NEK9Q
F0SQcg6/o59IBs7yqjW2eS/8T8X326d28WxgcukO/hnMKM3ENzJgRwtl0cgWiLdI7zODVqOP281Z
bePrFQsQr4vEd4IRh7RqVTMsn6lbvLz2F2XKr/ff1RTiSzI1sSXqIm3+ekiMUoUaobhvCyyVA6P2
9nRMK0Gq8RYo3cY4yjkymC3Sm64+YjVUKkoC7fI9AlHI7T9hKTR0puS0qw4aW5cuTlzQ3oB+zTyA
IDTCvoDLg039GQ8Wa9+H4xXZS4AY+YtfAOLSRpBS3o79XQQ9RuB5bx0CsSipC4VMVmY3EFmSH8/r
BIDKTP8xf7VfBwdwPK+wUV7kjbRgp7ouH5uQUe+m9GXYXJ0maNI2X4HECHcF1MIeYuVt2QIg8Hn1
uBkGRcD4c7N7blWFAZxu2vRdrgiZox/n6MoXk1f/OrVIeO9G14TbpPXHEsDAo7w6huW14+VHt0Iy
M+C8oAxYALbJ1BBl18NwX0rQyncTqv3cT1WyT6b9t7HlcFfQ0S6Mf6QndrvvSYHityJvzw7DvkCn
hmtHrFDgX9Z1xsbuzyKo+eWM2tzqF243IG8ekxgDh0apMGgShH6+41Wjyg8W1l/PPCQ1aQRWyUp9
miegLZxY5kxrXIHkIbgAEvL2a6ofrTqAmNpgeMbYAuFoHFkhHHi3Kc7t/LNCNRW1FA8KIlqvK1Wz
nlM0jA9+90wiGDbJ+CnUNqZb9bhYzxEdQJZZ7ReGTrKuzO45p8OgCbBcXa+YShOtoUgjVkUcMYNu
5e0qzxDS3Rw3CPTRwcwDvqwgwagWsbViN4g2bqAmwoJS+LnsA7Q6hZHq56LlV1/5T8gDKD4xQ2MI
Th9Z9XoyirfqkTD+b3L7Qyuz8dNbuVzAsnG/MuG6hhSm6Sz7wtfv5Z6VE/1i0k+sAfKaRGdg4/vF
SOslgF1WTDzoAQtYuRFTRjQoZB6Vi2m+rFzw5v9tQ5ObC5yZ59ysFHZkZX9xCHcw4YjumprjiISi
zQ21Zv9WAqsuob8bDo16OYZzCOHM/MAx4+eF+6adXaxlkUJuCgAgnnfWLWwFx5lkVgiXIyHRunfF
SankpBo+rSRzpmyU1w1K9K31zn76eQSmwKzy5nMdPTp5OBwiA4YBztb9bpD52C6CpmO+w20mYMmK
hL7ktfTD9eSU+lqlV9x/ZOeTgDiJ4JQlzp0ZZ7fbWEyaVw8lb1wOwIYbeZOcmIA2SyZTr34KWzwT
XHo/13mO612BYfam3w6wlsdkM9ckOl0HZh/jFaPOSad4QY8lu4E8/odhIK65tEHyEHPaWHj4/1sT
gEIeq3KVZeVy0I3NsraGuAnUSJQTGHjGJKks71YLiDn0LLt7hMWebGaM/H2Wa+qPkdP9D7c7hrc9
uZdVs5KCr5Hl2uxcX1cMY03kq6o5DFf6rVDeEXTDJBqcxP3gROhMFE6g1pfd+TRnGt0rq4MtSWRA
5GCkAaRUUJIFMqP6P7zJ4hlxnLb5rX7FRODy8dZY/hg7jTzzYWgzy3bXlRMq88HNJfvz5tKLF3Lp
tRqCLOVnlk37cDzx/gpYFDXzTMPD5PBViBOeFGakKMS5ye2vPEGPQA5wBX6wtAHTkdBtBDs8Cc5X
Iu41tnXSgCzBS8tsyDIphK6k8jo59fuFmBmuxQR22Fjj1neTeXa1rGtiR2eEA09EqY1KQkpK2h4A
z+/zDtgW+1NW2GV0SLOQGSocdsCgvl9NK1kj8kHYfpOeW0ochhL//n+A0FACjY6eQh1fF0rEMDeJ
/Eq8/fs26Ys1CtSMcu8YdTEFWHtxq47u9n8Vx+ijSZL+MfmNn8gc0u5fIvaQCfF25nOaxjE5LRdC
pYs/RBl0ZjWFiatd2tEndPkkD6rAEPpl/GqgMpB5PtUR/M7uOUPVWHMYo2R8Ur9TKgV1B20iBZnV
SNjupsOOlQkcN6wABWJRFFviZ2dqqDdtU/MlV9je5BKcdQMjy87iGMbmVC6r1vCLkJMhBoCFbf5+
ttufJ7XeOmPg6j50gb3cR6c6895Zv4DtFU0iMBOtXIGrZfhkwRQfoCSuz5XyDF3qiPC9UcnpTesJ
FHQB8a9lWDKT8wbGK255oiM3c+U1jDyJRVZIiXZua0inRJvLkeRABcn+fhbSV3utD2F1A79Sp7qB
i01KwCDVhLy/GJh6TrkvTuvXyFzM9V0V/tMTrPVEtc6I+vJTA0tlEdZSG+Ap2a/WtISIzVefeEyT
5UZkF0T+hTEUrZboFVo5ZiAfGnMCyvB8pBbXFgh9WJdzMC49CqHOzGmeylkvKTXIgtNMeUbRZNDw
+Oy/ks7X5ITgA75gEA3J2ek+rmrYqBx3sHfrrQ8lV/7PIJYxh8wvxYuoBa+LXZi/0I4XcXXTHs/U
iF4CMaNppf3Qde9td2OPbsH8zQaNDLPiemDEGYiPGYbXW13/u2uq/jTv9VxXswawr0IwKGxwK4zy
jtunyWbB2DFJuCPRAAic2RDI0gaPSgxGRpaDDwlsmKfTuziEDN4juf8SUhMNS7QegufU+Dm68Cmn
vHDaH/S5uUDCAQHSmJfdL6MVhnOkRCIoZLsEFlVjp7mzdpOrNK89U4O4g58oDWH3+WmguxDfLfcT
0yMTXqlb2oQyRNSO7i3eZut0fLaRLt+yntNltw+29e0naRakW0fziuMQ4lOZ6yItwzTZqkkzinzH
gWawfrfXHPwwr8u3fIxvSIo2oaX4PTyOfXbXIltG1dmSjV8E5nDq19ebHtEcNSU0Nv3uKfZUPcmo
RcYsBsvjkUXfkRrorHUH9kIwUh9ngXqoJwU3Zd2jGZmsCsh4DSJBR6gUJer9lw46lC2uM90xQt8n
qbi/BRxv/VXAI7vPsFbCKIlerXTwrJle12WwQfB7Oh8mOEoXJwASEJIbD+jwUITWgFGT+V9we2w+
+rFXp+C0LDZLsnbCpt582dUVgLLrXd7ysRf5BR5aW3guRXVmy1XUTAXNXmaN1mTDpcXiNA6e3FEI
ypOLgNSoui13qZEPUisqSfLMYyEcxgCc/MxK+4LhPJIuXB+csF5gNAzFFEx+G+FoYXo4wPV5/sHW
GJdTPzk31mXSZ0XqqJg985uvfUVaiM+i4uLi6fVKtf4G00CuySSiwA+ZnrNNosV/0qRktD0qW9ox
dk+hDzS3F9VFpLus+e7OUer6/LJZyJZ7JZi+CdGba+Rn91Iozl7Q/MM24smLeUf8jLP3iuE26qHe
c+nvrWaIld9532I0O7pk0U3Q68HHEg+gTzjQp4D+uTeJZNw0lpIDpD6SsNoETBbF5TW9SmVvoYFw
FjK41yTDqjYadbMqY7xqEevJp4pQTKEf3BmYRtZ4/XHLSJzFWF4kGiqV6XTTQxrFPE4bwyLPbSLI
XA7G7syBoq4DcN1pq5bomj4dPSjuCysbtT40jMxmNHGoDhi90s/09RwL5aNvhIizstAK73yHZadf
5c2kXWm//heoN2SI34+P8KgKpJoK16Z4OTWMP327SGhjHujMXBxUjrkoCkHrbdrWAYRF6Hp+mgQH
WhPbd9NptYXHESlz8ZqjVuK+8D9GTJiaELltWjX8VJ8iu3M6c0cuKhU0e+XS5jNsiuJoosAXzdIo
KX3JmDV/0XZbZo4Vz8Mfs2UpanC2MOa1qlZjLVzAs86wcI6KTG3WzgMyXWNQ7GK63nU+R7TGbDzq
+9B7Sngyh8BeZOhbp+kBimhUM2iIwppDkx1D6CBf2V3SNHl6aBDLccm1uLVnKeQ1dol4MFC9ZWiX
UtktQFFnw4Xif+0PKs+tLDR8f03xXLgkwwUwk9WTzeVGwgMQB06bQE52qWGvrAAE/jZcIUvVfMlW
2UPB6EaxjLYWEuUID+MfUglNalPyCrwAGxE81MbhEPl3eWHijyTrXe56J+S7Y1QYvOlZK/jH+AXI
5yrVWp73K7R4w1fqhuMI9C6tHJXwGiK8vpANRbuwJ7IhcxTqiUhFjEkvtggo6iZR6oHLyM/T4d66
Os/ALc0yXyzrRXu26WLKD66/BHI7AvUoxv5z0VMfHXh84qcUe0ZdmBjj8sDrU+x26wcgxO5A0Vdm
H8SnaKsKqZG3UgFA3z7il5i7kU6jzoon1LCbZ4RfkfS8HhAx/2N8H4WOlrPMddHjhZo5jfmozyay
ceQ4cHPDsgjw7KU9C/BZdXDSMOuLwgwA4rbyZoJ+6OUgK/B+VdGf9VfooU3dkpvavy1AsCGWIuSr
tnh0wPqcVwCueDF7BUytUfZ3ZxIW7cG6JKvXWeaorwJyRHSgPLul5PGUo5xoL4cd2liAEfUXgr+/
rfCMLpV0OUS1l9PN1aVJjSfb3aIYRiK6ThMakOKinaYRCyK/OUrwcftAVU4QCmueDVy7miPl+2Ge
5pklCnddyyTjpHdfmIr+Otdx/XADP9aqABnGIWjkjiYK4/GJ5cad7aIrkEOheUgX3ssM8YzQCRdI
65aiBV5VZQnHMhIdryc+R2vHHSc4J4jvstfFns54EVMaYXqPvjhPXulVq0fgpywMyE5vWHIx/Lot
bLbXDJsl6D5+o2dEZQrvUNRi6jbMNryhN3/gBjmrmvjlG6N906A/bdX7D0to/1KmcNsGhWLh+IFp
S55k2f/afZF0WXGis7AOarAM9/rNgsrevFh3lHm3kmn3OMMkSC60YBc09xcR1fAdrZ02JXBSLNwF
DCOB/+TpvpOIJfo2kBpqrkYWgd+XfkrKymzvFZST1+BDpcTHpUaQKeSZZ+1gZhjnBiKl86UcEDeh
f1/V+iSe6LBorYCbZxI1dTMTs18tHszss2XBj2Vp8G9kTein2ERQJAq1dEU1GuSbla0GR1Fw7rFl
WAY6N2SZfbFOKrY6k/VarwdypaQ/q+EMV8vXISr28ndr2OBSwwmom7gYPhJibH7JYEn2GH1matfX
hH7ekjaongWtG8B6ft3ik9CZNN7NV53Q2lU0PHI8385Qc66inkrtTQ+74P3kwU2De0xh8GENU+0y
ylcKd9VyFyB2HimsiVaLPSdzKZpdav9UhbDZ7QufUXR6EBJQtAgmuEdGo1XZFffO7z+LY52ix7sb
8BmDRE4seuGzMttPXnuBklEa/0Jt+SL6y8ZKo4AY+4RGbjzEwEbnAHJTw9LuXUKaxMWSKleD04FD
w7vFVCuyIo2ipKQo10ZD4JBiOIcgBxD+8XP4luKuzbBrwG8nVe4hHCV9KynaaMcPkbJpzXRmXAk6
rIa6WQqCNbIdl1HSaZPh3pMrmIUFClPFKmdsskN5Grv7SnyeilbAaSFRsM0yKNlRceSUZTG5vJn7
Os0XVpL2Feyb5XH8vzL63kazG/eQWYSVUo79bLUgFJbc2UwrNL8Z92y77xMDvNzlnLJR5mZGmsFe
IiTViYCjjAEB5YqDlMLE/z9XRKt04ZKxmz+uix3yTea09cFO4/ryANxhC7mpj73SdTSuBEWx8SNG
ulLT6u45a+YizYxGR4S9mnsgUEXrisbVUq2ZQgqfWxxjWjxeSUHQ6SE2KmTUgHjq2UtTOuXwCYku
9PTV5NI26aXFL8zb9+yxz1NUQsX5IaLsQb0QRB52XcqtinmRDxg753AbqF2SimoUZYEgk5r2g27n
nM9f5B/xmOZJzLlzveQ7mIO/iHG1pmhr31Tvh3Cvau05ScMg+445wzWj/Rs5JjBLEnIgM5Bw0oCB
45KcUejDZgokx5iAuGzNEXdCFREXeFUeKzkyVCLKR+RPEFKHXcrj+RxNOX56Niw/Zyg6Bs6dheUc
WR3Jz+CdxhgOJcQe48m3rbad4l6DzzK2OWqqL3AuaSlHnHzQvKCmcIv8oPntUgO9Mk4qsnanEoJu
02Cd5/zfCJc145y8yhA0FON4mz2gzsFSbHYQff1hZN7orX0d8c9CNIOHqZb8VX04bxKUOXfaVN5H
H+bkCxK5QL/hzFZZPK/83YXn0nJXMJ2v9CNOmbpWRRQZ+NULmWuxGih/sLajPMKuIQuf9F02nMpI
OFFqGFbuyTq+uWzF7Pv9AEOcWYZqXHiG0EHZmsrWZjmGUBxqseF2nwX6VerxwXI6Z5fYn9kBRIrm
tVBp+yvH7+Q5ccHzajBuJ2jAtvVPKlsZi8rAJYpOYAWPy8OqFi+Y6jP0x066stWCYhhAAkDaNsmg
n4gnbIv4Wl+uYG+ZeUxlkeHPoXwoHsuJkxlgmSVc7FHf7CW5rQwscu8QmW1JloAUofi520pqPs9F
FSpiVF7lEPbhc0rQ5+kbhVwjtrok9kzyWF2CNWIq7BwwWcqmfsCvrKSjGHuKn5LtzmCkLffMHpKU
Y3jlxlPXOCMQxPg9k2fRdYeNd9lt31b3gU0F3kImMEDGmvbLQVZ9xMwV6zLJSajbOCpbwYA7gnhH
XCl8QbLM4FUGVG5mLjl+RVKYHcztZ4FYb5nvetiiKeP5A4bfLYTDXskm/x8iGPrnkTMyyk9a8hch
ii0ByiJmKyxh0oUl96jquHc++FQ/m3C5b65UllVp94is1XyWePJD5qeaO9iOjnd/t+/7aPOrKlAj
0cZrkaCyiHamAb2650iwxyk736d518gh+ftBzk8/r43GyOb4FdONI2JakSaysx6rewDBmocNR7xr
PH9oYx8uN6EwM0BriGRD0m8IbaDnl6uUe1YBt0ko8kZPGvdwuTLHGDzLKoo1Nk4W7c4yJRtp+CND
5zCjmuisn35fpx+2w2oCyZw1qfXcarjf/3ERvac/NOMCR7JFchR8SqIOK52vHP9n/Dcfe4lMLjZv
hSexcd9zAutoF/xn97KYSJjQIOD87DYXQ9kacFQMkm60kCCdvUWVLLAvAzg/Kkh85ZsySNVGLifM
kepomYtGmtx/HExxuV7g3k3GmCXGTOKolMIg9jgbSxdSUEyWJkkPPHE0HM703ZrmcorDlWeWYTuZ
l/dRt54pvWfUIBvTEcJEmFc1zqv//c7RdGoWuyktcmM2Ofj0b/ZsZfbZo6Cy/TfxxkkK/NfBbhm0
RjnhDCRFS2fNCgohpONfbp25cIuQ0sbXT0b2f13ovDyaTwiKa12EzZoLdqH7R5i7Ix+AnwqzhkKM
rfa7fyYo/SkhjZ1VXt/0jT3p10pgGmpoqSVo6JOgfO2HRBjQM7GfHvgiYJsqeihv7qy02yvblxN/
9CFw7+/HEO/4UNfU3pzltQ9V+vdqFuTx9upmqsNLxWIfIqHrAO9xQ0KqIVmqB07i2OX9m4DynnPP
nH/vGinZzGrWU27vGo5y3HsNxPjS40psB/FXfeHwWkB1FfJ8OqFwQSDFG1ZprkS98zIOABwdXMRF
gfnz3s/hbjRxuCtzevfMhWjExXx3YAsCefC1kfQRPcpaUSZaJXd3dpdH3uw/medHzA+omEXtW0G1
HyOi3v2c5+i5Bg3n53ps8WNM769V9Gymu8W6GGS83pJQr0sTTCD+xzj6j/GjTPMEzDpMXE8JW7Uq
HoKPlJMhn36q9fwgTYxcaEnzmj7ZcYzOPRA2AOyZwHC/Y2xhFzkqv4OIn8mEfvHfndXkQZSnr3/r
ZI7y063CqFve1GpYQse7mEyiyH6PKY0sm4UhuLCjXm7X0JTartjVJTSrUtWHpP29VVewq3gCbC3q
3jc0Z7rin9/IS30cV4Fc88Ztuy9f28EWanMdLYlqngMtDQgjJRKqjqijKpxIZw6rByDm1mbWNpfl
NGwP5/rj0+2zhXz8zn+e95Fg7Iz4hRjPMx73w6XeVh3VUpzQtFVFMjJOqF0ntKrJkoswOkPiveFU
edj/98DtoCyutnWBpFn8ZvxbNqOPMbkh+IfjtUCFrxf7+eP48HQ752oXpYPBGkRjRDteJdx4MKf4
ebcB1IbLmqZkJ0q1p3cHdvGVHwPoEejIjJCD3kEp2U8HUxspA5ZUeXwJ94GupV4mCkftrwGSN3aT
Jb/b/uXd/sgUTW6Taf32thsWSTMW98wUHr9wjByYAkF6Axj2ev8YC+FecU6yL06cihH1LymONDsi
54R/H0mK4ET83AvvS2rsAjbC0are8Ni0tjoQ3RMVZrisf00VHXuYQ7at8Zzr2brs5Srz8LtNPe+z
Uehc8COyARE/oL96i9FwQ9kDAdFmCOKT5smWuIEpaQQwICvePpLlF40T+a0hWUYwgmvfJ1MnN/YZ
0eJSZyjiim90xZgA8UpC1WWWPKtyNTYaG0e5JM+MzmurJXnonmsz4D941Fe53ZWsbT7PeZdE3p4i
L3OB9hnphtJC1hiUluQKJpy5+GpL/NpTM1XhzR3zy+WlnIuXnp7jc024ftUfkqCYRGP++ssdsS1Z
AdtzwOttct0qmdgE8TwouIlKSgsdbjGOOU0JedIkjHLtSJAxOkV9X8dvCJM2rk/GfN4h5UsmW1Mx
slta8MIppsb4rG3H08c9sDBDf+3SAQLhxgfEfkZhFRM51Y5QKdAiK/68/OgwNcsnATtK7M3LOBAn
i3PDnMJz/3q+tpHy+H1IzkoW0SA6FEGHxT6h2qPPM0tj93ZD05qsclf1wjiEneyt7+VmCA5yC7L1
tGDEYUdCMS/xBoCLso2xYhHUmUi5dOZs+bK8A44kMR0/zoA0TXmG3500LSkp6vcmInea9jsKsemj
vZ8qooGG+ANYPGrjzMOKF0aqNvUsQhvF+KB5gsqrI+uJLzDjgOprscEVtpXm3R5K1vpr3YjfQ8yq
XIOiqQtEwuN6s+2Jiy6Hl3mPVIe3f+R7xw/NzQ1M269uHSIajsU7hbqNohRThgJw1+faFIqgObTL
6MwHAZeS5pvtxgMfv+O3ZgJ6wgKhwx17bYex5UrW9d8V41M/q6T54KGSBk6FlB9AxYx0rlrlTqDe
m8hFMrIY8niOY7tW0ANi5DgWP9c6iljgmu257rfjOmIt36q/nFnmITK2YuF6aOpDIlynHtfzbXYQ
mDSyVgX2Ksg8cxUHaPHMTX4Ba6fJaYzrpG4E+xM1XbT0TClQTPJhylRkQ8o9R6oGHksNmc5GZBC4
SPMrCcFGOiz4Hx6UvzaDO9lykIHYtIa5hNHb63uAd3wvKParLzqR4fNuoKSSyKWGUKBvXUjonNWR
Rekmf6LACx96NUYcPH5oN9mKhtAFdPPuqWn+/JnTJP8lY2mFehhhP3PGEmzuNRa1dNn4GwJ0JhBX
LPg9mewdR+/mG11rYW4AHXL/cEyDPgPdmsKcv0yuUQW487KW+4d4WEkv7MP7g3RUDo/fkS8cL57a
RrPabUYDhULFVehPlrKD3Nga6RNAbW8F1ISOHsHcvy49bEGimuc0C/W1E2t2YrkXfETlvoB8dcF4
AVEa46dI7MWfOqLyRB1AEO9+RBj8Q289GSQP8UxB3Xdy1Bd6q7oCE2Ar4vuo/04Kgc+U/annCxAD
svN9fU+oPDBBBw5rMtNygE2H+jzAdMYtUMzngQS5HotNn+ENlR0yfTPjm+LVduZExEDxQhAjxqhJ
8ZlGhtlcKqwAOJFFGuJfej4KVVrPkH4xibrah643AZBz4E/7mPahKDuwcuWPqwcSPOQBvcRoQ3+q
FMB8l26J8FWnBgbbtz3mKkr4gtZOMm/SHaqJR89qkqaWk5usiBL2+4/X8n66Ry68FUJJJog/Z0In
Z5xn1bd6xcuM5LYiViRiCwR+x4EwHiGdSA8iDkLc9K23ka9JaoUS0GcJ8G5zci2RvM/BbR7WjvIC
Y0t+7ACIHoIdUEapSppUDbRhZhqeYpSVokfIG+rsf9GPCIgPAe5x0lftTcQ6bdcUOJ3s7E9bCYNz
Od9r4VVwOTwpLJgu9KcinRuMKtaKS4KgdeETv6cQfQ0gBxwJAqT1AmlfkAzXWbnDzQWMhnofSyTN
Nplv0I0Q6RhUMOfyFhGBWWLUhDe6wHzvqeJj8QeFFFqpiyOr7T92oYfXsguX4cbosZZ/IXfCw++p
Dxv7iIezx2QkkDsE7IR/2w1yyjpIZ4rbCrNh+6GTGICcfVP4i78A/3gy3xXzGgyqwiOb/4LMiZwJ
w90ymFQC4ckoiRz76H4clDHnYs2pmQ44eW0KL0n6Rtl096dweurtfwrVzhZkQyR9sw95ye/3Nv61
LfB1QVa+YpBKQqiXnK/vPwcScv99CkNdpNIpXU9fT7xNgdVTkj4ryIwhBOne+Pe/ApwWAoF4Y76S
stryEKM+0jvF7UhpNk8oJtrydai5vIBzezBPzxNGSH8OI7Ax8/9iek8JQoShtS3Eq79TJTgquy4v
3wccrzkkVF4+Vy635e5zWJTZ6p6AmII7RXd5iPPs+SzFzdK9E5L7al6FS/Hr/ij0XiOMlARs5uzT
+S43j/+1QVecD1Lpdrs/c3OkF+hsSWzmjgnAyAKU4scnMp7gNlu00ee+CEZPzbijSM3neuFpXFZm
sZB8W0b8vmFeZyhUoFzV6KEeiJrI1aM89wT5DKHDZux/3QSNmYbXS7VEYkkLLSBh7/LgvyE4SHj0
w98k0hCM401KASGkoBdAwTZLdSFcojWBGdD+tVyf6n9ehvRhPRHtygVj0gG2OO7TCCJIN9FIcHAe
V7GhDB12pjjo8Segs15KTYB2EiRMggayRCP534HgAW5S/fczxCPQQTaqf328AxJjh0y7KphnjrHv
TypMHUfLy2scm68Vwy0qo0t961UhRzKLr0gBiwa8k0Fpb5RgfdrqpkByFZifJhOlOBr6Gj+xsCsH
FehtAmJee9LPCAbxY66z3reb/tHKjmgHE9z9IAgwRc12O1UhkMG8Mp4rAOyStPgp87tcN65RWn6w
BKEaYXQ+cF4wBv5VCDaCj3OrTgYxZ4qJVUznpBpVq3K0KE4rRATq8A9Zl8uxRee5sZ8nWvFlplGt
goD6G3PImCObCK+rQzQW+3xygW993t6vEgJjP9QGJUhaSWBc4m+/johtaVFTiOLRmndfd2eWAvwG
xGAOHthEUNDjN+kkU42UzFMEwGFrfwlQ5BYtBzvEU5BSYD2eAMHUHMtLSO9bdv+6iqvYMUW+oAvE
Z6VHvyXdoQUHwsSEpNSidudnEQK0eskV0vyhY3HZfsQLF70jZKpJVzMjyHzdrNjm4eWAOrGQ9DQE
jRDItuqg3b9u0yyQ8ux1dMLLridd7EI3/o0aSy7RJ9PKLbxJmrDtXEOeRosYeSq4YblyUo9bEHI5
mG/4fpoafdObdm6u1/omEKJRStcEOzLsaqbSEzFIn5lUG/lkeqsfhGfQAKpO6rbFSZr8iR3EXgyd
ibhkda1OIR27Ny44/16ufBdQHrjTQSgv5nDV+FSAZ4qd5IAglu31Z+t1bOTZ/KGonoc3AK4p6cDi
UJ0LKcth9m/WobIYWDVu2PvRBX2GUlNXHVXIFzn4LGJmuw21CIYlJlukzNpb3JmQ23AWHDC1cbIo
K9GC5iL3285cfTgcKRL7ezjeuRs+lLiJVYq9kO/fklPZHXibucfre71TcBfSbYgChEancy6Kxk+D
kgVyWWRblgQnoLCsafl6txbLgX/ztUBAjcgehtWkvgFK7VuscAX8b6xL0HBPHDo4YSGoAxw9FP8L
3UfVBy4rE/wzSYrzu6Wd8DIFdGDubjiHC6EWCRi9dpTMp69eYemyzxW3MOvSJ0bvpDO5e7XFYkLg
eQLqD1ybgeRw3cntG8iOqQnWllS3UC2LDTEHdsSmLpKkJZz8mFd1WaxeNl3II5AX2ZKtxK1Tyx7y
tzLc9fFl99BJfpQ+JeZII4iNlHbfk23A1adbzJ0fmVT2wA8rbEax41zAE/uaXsbtE6q7IvC+LG1J
inAUBOcDNbxycGbj5TtpS50jkKcwT4VF6y7cSzhn4FB1PqTYE+1a83NNfZvyMooxNinGRervclCX
YS316/J5DF+OG3BnsZTSHaDi4pgD2L8CPfzgEWol9i5eiGW1gsT6gyfAgDsc8GKj3OTfMQyW5UbE
/UzVbJuvT69edM8cTj95TpLD2Uzx+BLPHnAeHf8ZAicsyu4hXYfPWyaP+0snZgz1KXrAfBm0KMi+
glc8Sp6vFyzghfCiPeQValGyZJ3UAaHxnz8u8gd9bMBycInozrI6RDGZMqmeZdcWrzANHKF/9Ww7
KVYrr9zuwZHEKfIFAxZGVV4+SHsXF5yDBSTgIqcky4F6ioPQ2mTU7ivXtIsGZ5n441eUNkYWwB6m
ykiGW3gH/wqO2L1Lz9YYIvffbv0IJyaPrH4mlClJc5sFXMRHy/w7uDHSEQtYlJ8Oj8QLiQGsnGxR
AQ86lbzoT52xbD1d9dSh3dXh9xEZszD9oOoE/139W56ZLekETZwhPWngkwMpzBxW8vaTlaBGktR9
ee+2ewpZJPfY1ojANEGoWQSHXwZZvsJX0VPGXIX0lmzU6+o4eJoOyPW42dboDn8eFsAi2chOxk+E
WejEu3WD5tA9M2xCblacEUki1Fd0rvKyivJNka3UkRtTs9HzWYRK2mzGmNO7iEbkpBBTAfaQYdN2
cFAsHaR3uHksr3Wy9rDYXKzp9vBc57DbApIklwxVOi97FbNZ349Hew0noKhWZI9TPwiMqGlKwdNV
+0/EqbEOyJR4QuRv1usdbeTtft13EUyrXjgFACmaSyLa4OCdTe8LQ8GVOs/D3NSRFmEril4+3nHU
e6+enUBkWExT/VRsa3I3vY5VIeQXmTU8Yw/hxDyZ5MI6e0wQLpGUQ7nco/qUvfOLgmYI00c/9iUu
GD2A2Xsoia1AeHJGWlTwA2wflokfG7HjU3zK7ksrS+SlRhFQJYlzo+bM9C2ISsS7fnZsE+UkwPo5
U6jDhPwtmBERlGHVK2Fr6I5TzMJLb39wpH0khlrvmbMQfLwRoGBpQJUJll7AFoMumJqutB6ReN/p
7jobomQpxXZjL3ah4Ykl7nftWW5fzXXsCSq6BhFP0SWiYHiLQoxADvAnrtzc8wJSJVnrsMudFOEa
JqjpI57+sVE/5Gb+PW/rQD8l8zoNtPsEBTQ94mIS619q95xVXEnCK7MSY5aIt+5Zo+VvCv4LpEyZ
KATmwaq4HrZqoBIEAiQHfn0yWBSqylSnop7jkOCrJ/bmiIrxuQM5dipPr6NvTb0wN2wW90JvIhcm
NwRX0msXn65T0zvjSRQoywAqv9JJWDtlbVXWn0kdqPhOA0UN2Kk2uj6USiNanfWT54nGA4qlf1Pz
PlljPe42k5+HQmd7rrRP0jlgKNYSv1wM0GcoCIA/Zcy1ckcibL883pJO9Jr41dPZ4s1RMvdYzSLE
38buV4fAK6A9WZLdK505ZiKkmonpnMRUQeRRiKuvVD8kB9qW8f5RnxZmr4eBCSk/0ohTHnRl6Qwm
RMfzzDPJVc0Bu5VD7dI1KZo4aOUDlm5WSFxNKx8FaSnoIxot4zFJFPyw4Qr6gGiqKYroa3TaC6Eq
VGb91hHOM1LHWqjJ0nb5/o9F/0/q24VUdbLSNK0ZZflLW9D5FjfkVpjMNd2Oo0H8/3HZ3IabXOIE
xcahhrj+5Ep8iPK4lUOSCAa6XVMzx2NEzos/0IvHKxxGsL59BwNodMuN3YsNRp3+zjxD84IQaJvy
zoKxPorzpylHj3eMSaIQaFNDcznmKtx9ZR97UMqcJCjKuwizTU4ADOrFtt8clP+BzRQOys3m577h
Xs8U/trF8mF4q6/CX1hPhYnNsAfYpP0gTgmCZw36VGPi+w+x7435lMTk9B+Ajd+7o/B6QzOWFVgP
eio5kob2WeP7js5SniJ/8JN8KqtICokNgXV+cwv0ArE6gqt9unCrMlGfX0QhHySmRJ+DXoK6SsJN
THgyliCVj6nBOPuGG//BETTxk+dGryUgTt+Zbi67Nd1jUBPzaSTFOFb6Q3UbCFsVbHOG9AhTvAwU
bE9bOHm4zDZFiON/oeXSodBWpv5ojw4LunVMNB69c3MLy2Wyp8vrmBWe6JNCJzVGpNdPJ/vqAl8D
brfnuW8gytFYspbgU7Gy4bJVJkoLSWdW+9Zm+p4k4C1RV1crqKJaSScQL3tw0tFw4I3RTnRhByal
j7M+KLMhuY2TOix1KTpdiftxXGU/fTkR+FZZxD5ipqAUO8UIVerApaCMsPQJq4+6O7CCUFcQGo5I
3BXBWahzZnHwwNr6mdOqXmXIq9iBXB7Ls9ScDfo3jOfgvf7YamXNg9lNBDX0hquiFneOYmspPT+3
oWjdwm7YY8a4RG/tHHICmVHhrif4MZOu0oRbLscklSyxnK/bOIDO6GEOB7FlAkkQBEraci39WRUS
XxPWxaPvMo1jDqqUxx1hETbBwdKpwpyBzuVALDs2CCZrb0Lgre/KLE71yZSF+w55zj+mp/yyq/Ph
DtY8dbuCFU3yXPh+w6T5VuFqJ45ivJK7d61gWw4f4c4JiJjM4+iSzy3CFhkxJKuJMK3LixSxtlvU
0q32smtNmL7h8Mu9Q2Sk9W3EzGoYyxTlJbTelUBSGbHg/hbbvTmkrBnChjaV6pDZJREYj0yXodaR
BnAtcp3NtvVvZfgyBBpPHKyIascfurBISsEPxl/qNn5KD7gCiZeyVF/DtVtntlYKa378aEGjJ0F/
vkzRDNpr2onaCvpmYFsKa43b4Pr+pRt4B91JvDdVPCWOHCI758pRsIb8Y2IgNXKO7KD4m8aUzy+t
Pbuyx305j/13GLIflKjssmyRxWxFVwWy34AwrKz16BrEEUAJVXI5CPlOpw6Pc7lFmPdPMHRo5K1I
Uv0oD/h6zNIyCMcrnN8jfoVqN8oBin2065L3yxUxloM42Iud3SFQj0zJw06tY+gH725Rr83QzAK+
CdKwlopqjSwVZuHnP0qHaLjvua2yFfhJ5tFHH5LUteLe+Xx4OmcXHVIIaoWC2hoCni8Mg5/L/ty/
iZmdNS8yIQ3FvAQjSrvovUP8JpdPnaShncgXtgODg9BJNoxSZHx23RHjvsfiEw/4agfOntvI9Tmu
9I+AYAp3ILaeBGJgcQ9J9iNUwzTj0d+YSt82otY/r2BpZENeembW3Og0Gpn7Hi7Na2RBnO4wtYdL
y1FvWdorOuydJNF0UkM2l03cE6HMuuyf5GcZCaOwt5mtnaWGC7UZPqVLgI01aG0mZAYQsuvKN3Hc
Nma98k0Y8zJP6CpeVjj7qj/vNN9lPjln/2o1+RN4QWISiemPMy/yXPwvNEL4vGj0y40nYq79HVMF
sMC1tICfYYSJzVx1m0XiG9FJZUNDyEJHlV0QabynHTaAFUTnyiVd8dlIaG1qCqbMr7OdaQgiM4VU
jyNNP2g03oWRS07XZaqftCW2T0iTYe3r8l5spzY9djvSjtmP2AU6MPseUz0/nJ2b5hN6u4Y3VSYQ
SBFey3/1YPiPsDMzqymCz4Nf6IGcfpNshnbUVDz25MXj+iUiOJRGLPlRIhP4bayLxRWnqiYsHXa6
g3C3DgWfqMeGT02CfoeaGJRk8riVxnCZtNDNOPpAvnpA/xOMNUk7rXspBWFV/mtjTH8qjI/OGRb0
8LAEUez/2ZUUQe49vhvY/qU9N3R/O5xQmo+v+kF8fM3ghdxk9xvBlOHlI2RZ3V4QoEamRw1yyIrw
DD+ITYVk8bMLsUER6BI5MOScN3BFKVjkKk7yj2fNvK0S3Ky/peBXKWQUzYynCdbh+slVQeC/KvI/
e/6l3Y+n7EYvrpXekqhPyYaeu6T4TJ+0bNMMX1iC0Lm+LfDlVwXTO0+B94DY3LPAhEeSXRuw7Zky
Ij8fpJiBs9LUQ025242RigtySgUr1+1EEk1wtfYd0oGBJrGHgI3v6dqx1zj8PrOMGRq+HxKds+aL
bxe+LTQwKwLVTiCs9mv4e/SN+6+HLUuPVGFJ9d/nzmOIUKI105KwZh/GTfLSw4llKw7zRRMIt5uF
kJkNzEnvzJ/R+vDRCHkQ8OxYAqzIg7NLCng4xS13aVEWEQmFcFK++nBFjGGYwsYMibIJOaI11Tqj
cJ0NvXHN6aVaCYaeswMOhu2lvdYKZOcbD9gwP7noQObGvl89QTexliFL2LFn7JeT1i6Sf+pYlGm/
QJnkSpBqAHU5SaFFkYeruPYN+j+PBWQfc8IBu9zQS1h4JRolaPkIbtxs9wa0T+nDDAVGS2DrA67r
DVGwblcjflJS3ommWfU6n+NVrBIDUjVN0jqLl16H/mUh8mfBe1Zz/A3H1q2j84sVMIYWLEMss3wQ
QBrfqUGpnGXScgQzxejvvHMF8EHsB5+rmpLtpMKuYWLtucG2tB+MLvWKMu3+RRuB659EtEJfpcFr
4cirK68cevrHiZIll/4vvVHmiPa+OUoQejZMhVLdlX5J6rO3D3gywHIVJ2ycdViW82AcdurHPTjP
aKIYfsYTu6GJeWgd+bHsmwt7QnpIwTi9IG75wpgoUi7QZHq0gfdD7UaASeMp8h/iqhE+zOUJmcL5
IvcWBjq2dN/SNXAjSoAfxsWemSmKtZQQba0W0My5wSFNF9FCYaoCefYXKpOZvny+zU76KB4b6TLX
no5EJrq26XvPfdVrqDmK2xkiiefqISF9xgWF47jdIaWCF27uSrCsErvJXzNbxRxb9gJwxIaR8fVT
fB9MRJyrMTdYkQFnPqaqU8m3I8dTQP/zciqoFxs0qho00ot6QUaF4HbiyLmuZvR6CXkURzk3DF7b
3wfLRf++E2YGAArTulWCucrWZ9te9QZkESEJ1ct+ool1lRJjBPcXDZ6FtLEEf7LxJBnemfT9u9N7
t37m0IOup8Ja1rqRgXNj7GXz3HS64d3BPy01Zh/c8WWqTKhIVKtBCEQVHIb9XNzXLhOOwbvTWITz
fyOzab+5volXhYdUOyau033z73rMNy19ybWaAlQRZxRWqvxyuRMj5MXU+7IufckFZojnGkPzyJpb
TM/vtn/7SXhefOtrr56JuJ7F35snNtFkqds7ZDNTdkywlo7E7VtDdhR7htUTwQYrHgZIxULXqymX
6j9yDGWhjNXRqOx8jUJgYu0EholHbiNiXl146yb3futSYpuL0Y4jABlS2uIpTPT//Wpm/8vl6O4n
laNubH9Y+AXL+8VJk86WhvSMvR0G91oIIqE3HnGY+5q0cs7pLDAzCVyOXSTOEs0n0L9Np0a4hWS5
7cqUaTsgxLfQsHuZlD+zhtRyZEMT0OduWB7yhhucrUMSC04YNKdQkLskaujSP5lFu0bspPRsl+xe
jkbdV6MOIRblyTY452uJ8aGd283xc9MS3V8PCgDKmksZnmh6+vOehoCBWTAPcsNtlPrnTsK7WQmh
i4vgsrE2HAyGGLdP/WWBIBcd5yD/FmFslpdFzomu4jXutVboCD6h0D7CFeF/nk8YzBh2lLAdSEDv
iNOQlMAM3hIdc2q4mK3v5Wu/srpLYbdhv2hPInQ6b5P+LDFK7fGCfYIwnjowtF4wRrdKNnN9wmZr
sZqyhVU3DhJvhh0eNQ44ZekMmb+lkJutADiNT1CN94G4HYQ+UmjWVilGl22vj6R2qOPnGDdLZcgA
bpZw5G93H2/oXj9tes1PvkhgdO8703r8uiXCywnwmgHNhVhdJrU4W81ugs4MCzefL8A9l6CH/s9e
L5CwuQMMbd07gsC6yiYHv8qq4iv4sATM0F9VtUYGdiB/xmqhPMclMeLFM+4Re3Cw1MAjBkBpKRVj
mFX4/q83P4Xl9F4fsu0UhLXi8++0stB2eY9lnDjEEGR54UkdX5QU9nnOW4kIiD72WtwuTc+cD4Id
U4+eQ3OYLZ7St6hZODbSejVjjwoz4vGCJx4MfQ9XAlej1KP91paiC2EET24TibeQgA1g4SomXXio
C2nHmGDSZu+qekDgdJKW8ch4w15uAqcfh9QDHGiw73zhYnO8Z8MGXpywiW+9hxMDkVO1m78KIl5b
j8hfzW27ruhSMaBoaVW+HMpANZMx7Ft08iXrk5inewlWr8Rk5o1OMVI0F3P1IvabEu0II1P9xhR7
v2IV6z7qpMAZeTybEgxEPbv7S031dpY/JTyAcm8x/RTBO0Dax9gt1zsdbYWBtD1erLOCOvPzeHef
ueImwUNaJwkGtOJxDNgBV8O7VG8o4WeqU6g6H/bA9BvEMlZuug/ANVCsJ7z9x7l7f+35LrZJRuns
LvwRE1z+Am5Z/3wfBNvWMfGz2blnPnFhAp4aeCt4qtiRv7dhwtM0PTL4rxhoE+91v20pw3eyxpWt
xL4yMzSfv9Jff/FBZn6rNa1XCuS/56ATeaKK5beTd7DIX8sIIyzEDdjYyP5al/wMKy7z1wbd6kYZ
wZ1RBXAxtYYJq+7fvjgCFhI/qTIAc7L01Old7FK/PZXNAfR2UC2wdmTwcEu9D80LLd7ELijyBmzM
hBbfvAqCeJ4WstP2njMp8I48KBEusJD3T77XwYY7g9aWAZWxt2AfndMk1H9a/EhDdO3P/msH1Yus
nA2Z1Fcf/UtvuE7RryfzI0T+Hbl2uTOJRaGcIUmLspJ1Mv4PnwbIRyN/PLSd/ZALd6N+oKxHvC+N
Hf/rfW7vClCq2FMPEXvPUkKEXFfqbK+D2Bk1XmYus/BXHiBFRzMN6YP+sXKfmjDCKcUkdioVtgrk
RcsRkwex1SjjBqxbMYRrvS9upEsG+SjM78JwYEQwpB94ZEE8fyn1ViHFww2xqR9fLVV9+SwL657O
6vtqYOHurid0XPO/yLzCWIW6wob4Dwfg/xYM2jpAVKcaRTTABacnNgZG28ObZhF16xEv0p86coEq
X620uXCr2dQPNYqvdaSSH8OEm3U5Y32ICw+gTzG07edZl1NnQUVRO+tmKdxzBarhUwL5hJuD/OqS
OtGXbt1BndziviPxf7nVwk+Us3gFjIsFB+bKrfmujODdwsZMJN76s/hGRoSPPWZ4bHCvvUB3b4Aq
boR0Rn8rVSZ1v1LhCoGtox+Qqvdno4jaWNcFpIMcpj86g8zciYhqfatTDghxDmUdW5VPGfNPH4CG
/pUyxPb/P/S3zzQy6UiiGgCswDOvjdIY1QK2rUoU9QVhLOH7YWflSO+Awph2FAATHAZygISogx3w
TJE2jba2xKU3E8NcUUhR2H9CVZemfVDlyQCxGPi+Ub+XLcxqLgbJ7eJYfDP/GHqlRnswXlWPGrZe
uvlOeKriUzpL9KIQTfyYBeScHYb1dmIHTbkn7xwezaUxgq/gMVlSp1VRpa0JRmdRp2F+kOyPR9Po
UX3LPtccpHmQRdqxnVnxLRiguKUDevYjwuZ2WzBUBLp1WZLr/PIZ34fAtHb8BA77WxNpFlqSQoHP
kB5lUwFybl2hY7YcF2WA//0Dzuzx1payiOTXfj4iVmA1tbu7bC+oR/lYLnGBOYJMomUuC6b7DfwY
rZ8NrlgOCyz36umQwCFCuyUCYs4mEkSCgEq1jg8KslscMnIyW8hKlOAl/VgI96Z3BX59hj22z1i3
vmxQjnviO+djHNNYoJSaTZq4AdUaNzHB/qJedrtCP4uH/cF7TcB8NQIpIq1u9i5L0yxAKrfzEw8L
QsxNK2kYAIJ9fDOL0i3hpSY3JkufUsY0Q4Xrxhu+Oh6mijQWJQBWS5sWWqW7kmIpLMmx8Wh7mdta
W+jBwbBxMvN9CexlHpl7trf4sCDU1uqxIO624dBAkiWvHmZmwjJX/Uv9kM2KAI3qIKthUo4zKWr8
4zAch+hPXbE2IhlCTwgk13+j5+/s6H14V+oqytaZVJ+CByYQyYs8a2/pfS2pj1RiDlFLC17r6z/k
vPf+L/jttkeM6OQsme/J72cEpCdt2tFMhLmgI1FczY4bm8yphJ18PEBmnLYiaPYdgAWgp2sEoRg+
rfWjHj+QAEoFauppniaRg6UNSc7gEITap42kDVS9jOHWL/XrXTACNYmDtfy4z5EBmZBRSLm9F13r
vrjWwB5MMfumIThWLWvfxKMci3QPmbm4FgV80c2XAU7Vhn2Cu6QIiMu1urygukLomvcphEKe7mIm
aDw2vr+CAeA7FiR8ikyUMYC2dHJJTh1RYhhpkNP8ZVrQrHMm5BvAgv5uAUxywUFPm1FwBoKXHi8F
orJLbh6nw6REZCwfge0Ui3ZUXyE07HFH2Bh9akftPf6GZOw5kaH2CkoD1K2daVonJS8gra1iRRVr
q0YL9d1t1O3pdlhibgZ/2vA4y++oT7fIKcYRo+OZ3FLyMJyWFjKUIkC8lS1XuQNL8iA09NdvGw9p
YN0kQ/v6H48Pjny3QONkcToNOaY89FPgzwSLIGrAvWax4owLhI7ZRXEqaOaxrIo25Rh8upxGKSNW
nEfVDMmP2XFjyAEwmjOcCnefnn4SbLGi0FiVpPKGbbI6IR1vr68Zb+LKiLfSOPiHoV5w1V51yp7J
xPAuoS/rA8M1UZgPRtl2whHj5mcISd3YXo28DIyYBo1oSHhCVyvkBGQh+9/agz84cMVALqkjWdRt
72WkZxkwJFIHJx7a3mZ2c2Go+a07UdSB8BzxvUY8EmOiU/sXrV+iBUeZvsVgqEZw42Vs8tRgO+Ae
8FlwGTPD248hJaMRmklpRUs5nBL1Ndg/jvoqbA4AP82t+zg16T/Ma/CeEGOeHLafyCx1M/h2QaBi
ExTRFs4k+NORJMx8RMguShyB2INlZIhR+bpgl4aL1IZf9YUHVvJr3iZiDeWwg/JNAv4i3iJv2BuE
50GjB7FIeYVcBfHfix8H0UeR3TDfUSJOmILlEnS7pDqW+OFnInKvJi/75LjuDgGNV6Kpfw5jAn9q
0H7CFx0fmXpvjY17IrYYhshfC0p+pTg+rzyGt3vIE18MLUCWl7igaumDFrwdClhvoaoJT4Sr5nAg
Ek9vDWdrvEF6bLJBJX2Qp4CRBVI68aYhHnK0D+xfMsQLbTQM68F7F8u2bjDSemifZXWnOq1G8hyu
FmiTIlEZd09FK1Shje7gUKpkC9gjyK76ajVT6KQd/bcS9m+kcnJQk95/xAzN3GIaYp7nrZHoGzuR
dLgCE2Rf9+MSKR7KpWI+EmMmICudOyN3aEQKwwymy00cK0H0BFwpRdRQhRcpScfkgHIw6Ufqii6m
Koyk4ITcYrh1FuqJ6N23GcA1pHZQI7ppgCQ92D/rcoeL3JAZV/5oNw+QvWvu0kYQKRivXhGlHmcH
BEVlEqHFaXPALyUfdvDGTcJaTRl98EOyTwrr/PyKoFKWHqGIBV+mYoBhOlclpI0GSafjUVWWW7R1
HsITgfUCGKR+llvgWbHeD5sOTzk9Jy+v83x5AQI8aLxThUP+8k7Zida3u4WIzfrsUiVXz8/R3l4+
ikLSLoe+CscQGEOS010oAfVDInBwSpnqt3XVzXSkXlaXSmD+s+VTJQEXd1u3gQ63GEbC+PjhkYQb
/VmmA0pgpuVMbinmOE55OrhlbaAbbc/uVzb8eKEhlfGBjudlnw4mHY+MlI5NBD+4rbVAdJ0VidqV
EQHHP6H8f7b5SFFndRm3GTZs+GNI3qTYtClvXY1NoHZu5o8YLQHOvh4lthq3Siv7AaQFkL7CIRoE
wb/AhDZKeOfHcBjD6QYN6S+YHO6vaGzkcXjcich6+Wpx9qTQacc1rIzu4Aj17pbflj0fmd+z0Ull
O8vx+N1jXTo4B4r9mcFxlxZZM+NGcAOy3fhmSfRZlW1V7Z1Bsq8mLMTSxbZbmxl63DN8/0ueXDkq
NKsX2pUPCnc7CqXls3Ni4yc/whOTZ+gUKSQUzhsRk4u2HB6x1gVIK16e2nrUkFgpO4wyC5nfN2+Q
7FkYVvE7iA4+pP00Bt3hWXFUu2a85lLt52PtoGesEeMu4i8XQ0O5zYArc3ORa+b/XFW0ivbk/nP9
J1wOZjl/cXAgq6K7CBd7DdtVBjXqFjIjWLyXyMGUgTi7tV7iAiM3M/HgKX7IU6MYtGOVB5x3JTs/
cSkhh4iRELD74VGTM+XXkNPftNWDF/Bo9LAMuIn20O8yLRz5DfaJT4+HWyNzQF5tk05O3bnmF+W2
0qqFUpBZHUx+kSfE4zfk8F8y3ornwTiXZbsbdKhKs6/HMAuw0IMyu8yM9XX4+TAzOuTauiW3xHmz
ABFJybsgKUceY6B5YVGarTf4yiQRATZFInpUjL1KzP26QcpSwwtsyb1FBES3yVJCAxXs9UnzdJeq
m+WKxcSLMSW0y0H836Ryv1eUGafmEc+6m7yZ3ja5SV+7K5cIeRrEZm1DnGoQXbWynB7C6/9VWjsN
4ww0HKnBQnj3/vWHimZkGz9Cj/Kr/s5VY2yRfV1FEghUrC7FlRISYA4ASkSRaXq+7mADPm5uBm7U
KJ9wZc9lN4bT9gDBYQM204IPXiWD0A1+gC00oEVgaYakNF+2RA9BksMZDGZpWsppEoe6G6+O4nz4
Z9XwYNfU/l9aiPQFQ3AtgeG6hVtr4zhmh609fzorQOTj8fonlkbGlXfqeRCxY7aY2oZ4fRJEZkMo
9e7RvAiB8IIcmx2e5Klgzg+6ImFIt3HyKh4qgsALvw8/fJOguxbkZNpFaAteu7nmr4FXQ9MMOaBh
GEoIFX6BKBEpJmY14X2M+/7dRHg21dyJJZn2yINYLhrlUklPOKS41xAyCI3N4bWI1O38aQP86NQK
Er/ijwtdrycdGyvG9nD1dcd23ROPzpD0QnIe495Ht/3cxv+ROn5U+5H/8xVb9Lm8axAHqQ8sBmOP
MhVbr+pJXotaqnLj5RUzx9PkCW88bNPoeQ/VL4/Y0l+PwjyvQDxsPgwyq4sjI4KbKhBeESVB8sfj
D65RJVs7nbC7t1pZu7t97lx2sz7WpkkXSIA25M8uPAGpk41t5tC+4oi2VHVAPHhCh5cSzu7n9LNR
Ok1eDdLPdwNbIk4BZNmiBLHTQhtxC9uMF3lQEQ8Nrcwy/gI8ID9+c9mInDr3dWlMOCs8xGVUoF7d
x7VOQmQsn2IcoIQerLHQmykmqG/EnFfOozBoq+kSR7X24jJkNlmiIXs/pvIU2Qe3lMrnjFM1D5Xv
RO8VbdmxE7p+RPyUhErk0BD0SeqbQcKFURUpFumlKUp+eD7qZJ6RGO6FuChQDgpbwNzIK+piqB+0
+RPoDsdf3okKAOEjKjd8GBwoe5FSyOuzeZRRK9T/60LEw9lD7Zyzd0d1HbulYFSTckPPt9wrwdeR
4Qwss6gdLSzhZJ3DoZfQnuxcsTjV27e5Ugqjn1xtbl6r/f5I161lrKNVBPLLIuDR2E384kAxK4WG
mMOuXrZNiR17NTqp7EVHufICEzn6L3mjKBDPWJyoDqqRcVWDC5vRa8Efp6DMafyAXy9d3XNvbbwv
C27Ro9Pwp1O5RncKAIMeORFCbWG4p6JDscymhn1byWY7uiZu0D7PGKeSyu5nK+M2sF1en2kYPbk4
YonFeXZrHtcJUOZdeCy4vRKaPD7zk4pjVhYW6HtMy7vZ8n4Q9IsltAs0zI/uJg/rw3vUCMVKYGBc
XyPtZfzer49rPDu/kkJbpDnbsM+ZmeptaTdCxbaLyAty1ynUsd01oNbzY8E4MET5aQCszsuGSX8H
fW/8Fpo3rq8CxHxX+YTIEgg78YRPTjJeQ7CQ46tItKwBdSn9fHYUtlh1phPs+3DVoSsgpmTpJXdj
iur+Wp+nxNga/D2XMD9xYWajlYXduJuxy7hYKm+wBRfOwa55Uq3Cjj2EFOIKUJ3MwbOjV/3EcX47
aUYQ/1g9outqogaR4hwYEdv7QFLN2owRP3m2qFsAhlnTH7DvMqaa/lyMgfU8LA2/6NdRqEtumKSi
G35dyO/K8bcKgQasphHzPnDdBq5n0ePhyjoSems0DuOTelx6tK45OHTq2966LfKEUL3ofq6j3KlR
9Isbxmg0bKWskAGXQ5IinvRQxdAbQ0dV4yt3BkjUZuK3MfYIpQSqLLtMmlqla39rv8d/qYDWHoGd
ckEOqAqoSX79QHWQjm2xwUgX+/RiS40TNjMbOtFFboVsZZAOfJeTgd7If5EmfK/zfsdn7OpxTur5
baBZbQPM0ZniGmFGt27qOwVS5AMbs1rO9MCamDpfilYPFKLo8uO+7VLRMzte4Avyq/zQZaADuApW
1rzaACwpbt+5m5nVyactJN408vP4PEST29shzfhx5yo67sgnp1oPRs+WC1I3euo6I8/EYChHZW7L
j797bPNC/PT6BVCXKG7gTF91kFLkHgx67+teB/hCF1Nr6YBmfza3ZaoQpNyB0dTULX/Adj0AYTQ+
+tXgtouDFMafsfZng0HWX7pFfWSRYxxJcTHAEbwHH64dZZ/eOHTxVf3Tdgk3ashy7FCVDBrO8TYg
8y3EXUdW0mSyqeNy+YJwFvSqEm492NfXVsUutGhRy4bsCwv7l6F2i4e8JKkXcYV20su6ZF5XNJfn
lDVTFcRonGH8C4Q8E7Qj0TyQsLJfdVvjXgYEqB0qhNlq6Y9jMtttvwWBRk2xapy2qlDKIJWuxgIX
fSSmZDCZZcGetjk3lp5oSA9jS8v+oR77ftxwz39m2WwSip97xsFmZ22BxQFjO7l21GBTbEqTcIBZ
p22i+PMNZ4PjDUdkom35oVkVICRINnro92YytyfelQuPCyBszOKiFfdd0h5u76nkZsExwp4zvp4a
Sk4yviTR1slFmePfbChjtkWZF7sZrGwbVhJrcJWaJA2aANvuVJKrS84WNUSdF5iz3Q9D/s2m2xp+
TwsR+K3Ci/QsjPTrxgzE5BdXRSHpaCJnEAYsksA4JmmazNp7aWtgXHx4YneuT8WYD4qfhJWjN/EN
vX7lh85ZzDGXM6/MUhezgLFh2ppD2Qw0SOlr2fql9ETQFeRY6OcTiKpouVhhS/QCpKroqLQBObHQ
OW0pfNDtvj8RffmCTUq0ZAEILV/d76dzi78LinXL2WIm04QXa6nWF/a5q0Mj/dC4zqlegeL+atCz
pF540yGjIBFn5p6W9xKdNfuzT+5Z8I9SzbiJIA0VXJGytbPtwCwnCgCdbUSRsoKZAjpJqsXy/mjg
7TwHAjtF9rzfRyoTIM3LVB+ULPkoHFkiVKrNKEonQ+SW+8TLGp0WDrTzdzqDRdr3Z1OolsP3HPgA
X9EmoUeI4gZqdscHifFd1+ZiHTTgwhNRlfttCKg0VLOuZtSpatn5KxeE8Dark8mr5pJLoqA8buF5
P23X4WgWpv8FvKLonXDRWe+35v0YCdeds4d73R7kfKIlD5lGBvTyzSqQiyu/xfI+giMB0qPw6TwG
H3Ca4qsuVV8ePBuXrLCvc1rklK08v021VeMPP8/cdluDU2/a9r9sSFsi+Ox0d41rfb8J4tqtFFj8
qzGhGS5H2phI1Np3574neWcm68MudZ22zFi+r6aWYTF3+j53thj8ZrJ6zwyUdi32rwDWsL3nc/5W
/NrbDHmyRqinX2p9R93zgVBVhLIZAVrFS70h3rniGI2oHAyzA4ZQwmfm4zu126s0KZGqLH8iIVUR
M6FLl9gDu27XtwlZFfOBHNk9gSG8r2rbez1Mcb97h+E9eIyN5Ods0T/ldjsCYF4+0iwOVJMJkLC4
nkZ+j3WSUu5kzR10grcN8qm4FD+RxupvnpCTMMxFzRZUCZay7svYFhqJcimrfMGKrDgdpgLHq/rn
8bWBbRk1P169lRR1OETv1LKzIHzpxuZlO+Ars7A/HVUCcyFTjSA7gIr5F4ISGqu9v6ahi9LXOq8Y
1AM10u6D6XnbUuF4gUcZLCs7fjZHsE2ARdWRnze5YPXFLgdbcQJ4db+q4GFOT6HhoUk6aiP3bDhl
qG7RXUEe5saaDXFLV6eWdv05G7vIJfd8iYzhTPxrwgE38TNR4TTi3E/SP964roxMhXk4jeqgu1dR
7sQiQTlDEB8sH7mkSEe6r9/PuzIZN8BASJcH0Oj95HhdHzE+QSwYRy+EnFR7OOJPImYvZ0DHR9KW
66f3yXUM0ugOprCcOjqaGQ+ZqYUF/HM/+bSOiAOOjmKWXVwrxzATUkNrDLeOi5kXJvCZcGCID+HT
RJCKMsrHdRvJLMfmm4kL3LCk50agcDndD56RKfX6dql1M7EC1EuUFDmsWRtGTeMX1u2FrUTWsb/+
C/5rQHa3xsHyvbnYurH86UL8hH1iw9iigfhLwBGCQHMsuIShpNhMDI/D8foFupB4m7OX+R7kahN/
3/Y24IuO5mfQ7NnDAH9l5dw/hqjQBPRg0ERiUVVFJcrPYQWc3Ww5cowfK7dbSY7ZImCedRhdiq73
va/siSwK7ySJV8x0qg46JBaU+EStJQk8rvwpHRxxPsBUKdfHFWXGtwoJwUSRrczZehgeplcBoq42
fr2/zK/ElgAyK9M7diFJyfjFsteEBprWdQFcwOwjltdgBk+0/EQTrq182A1Q97Cis2a1nbxo6Xz2
ZqzvCTOjE4mn2WSiiJLWL4eO8Np+eYHMgGksnQXwhxCHv+hSfRygJw0FYArV6ieCTZGibcG0nph6
HNd1/gFIFGW4uT8Y55dYzzNIii1VtrWUhjJ8FDnxIqfcfZpLCSznZl27T6KELHJuUL2zcw6mREGL
wZ7Fq0bUCV4KJdJGke2Ybrr2Bs43/bgYjrIBIyPVvUkch1hzkxZd0+hOVKNiFJ0ZPK00sWJWgbEE
YSmntYusmL+d7fz7uPPBqBP9hhoqe86AxNy5iOctn3m4gHn0ahwGrtKfZ4qzLTrzdrX0xKpery9M
9itX/wjMGtMwG66/ly3Ru26uPeW4oB60IRZKvLf7UH8cmO/U8zk5Sij4dDQYOD69BAafha2AdUgJ
WuYJDaM9HDzSTcHY4eW7kA/ql/fza+Se7iGbFVqAqzFFBDKfaN73cf00s50fIYtPW7yDoh2wGmdJ
6jfEwwYGCVb3PkWVy4MeKZhAJdicpj9/Jo2BQ9454D/r4YQ5SqIDJFkVBD9U8CwDyLiUtEC4PvZB
O1gBS5J0NQs72FE2RjVO9jjr8LllxAinxGlrfNq+FvwSBEEdyRhWG3s8fnY5h5OyhNBkVv+s72oE
EYQ3PWh7SCGSXoRUTLaMZKtzmptJDU2tuWaT8MhKjNnOV/1snhyXXvKkrsETziP4BFnQQdYLkMiu
Rs92e5d231fF1pY0mMwpJX/A8qmmbJ9ftxRnYRr6/iIvEiFDlf6vBLXAWgducqiKErbFR8taZl73
DRPYpACG2gN5T6MFu8YILC6DMMPRAMVTJrlq/UhAwdL4RuMD5ezJh0nUyGMnYAWRLdSXAit2Z5V3
+sm2Y0tLgygncU+fEfNdPzg/q9qA8Vj453HC5rVPXG0r7DMl7iSjzUYhj0XVG4nsyxw21LKCCu2f
mqUVS0LMW1Tq4NESVLVK5Z5pYiyRGBpG5gd8c88qKZgCY3SZsUCp4WTtVGNiEWZrzwYR8iI/aMYE
Lz8PTXhA7DvInRStbRjVb1eCSbu4xANkBbZBKpcCMORBAn5ANSHzyUYxQD5ETQTpCiH8qFcRdNFj
RemkLHSLj60JouoIwaWUOuqOXXXMfMqn9GSL3aUXDJBAAbhjpR5QUF+FbjciHGl0kvSMoRZJw9MW
L/X2qO8/C8EE88F2alzbMjp73/p+zxJx074pNnKe3b4Sk0PyuKABMFwdiS5AyPLtKFtBtbf/TmSP
PUkws//cO/QAmJRADblK4L8rl0C84VOPdMJIjCK+bm+PKZWVfHgEc2ZJVQYJ/CLBOO2RHfNpQRTf
gIFmdlJ+SI3D48/rEgjzM67DgagyRVDUk6PSHFf3GdK01QVQ7ong+LG6QzBdcRpAoXb6lgDIiTrC
VmUznY3+izkZLHeOtBgF6wfjh+RlO8KWx2bYDVcLVmn/UsZ+KqHQnMiR3HENlpM9hZ1uQbNctz9S
jHv4aNnbraQoRfPS3LoEzOt6BAxm8GYTi9TUpUHPYNcdts8zIekQPqVHpxSHir9q271Us59C/qy1
6C6RNRE08py9xHZZFQr1tUKLrHFghIf9foe8WGhJNbEO3E1qzDB6MLqDxSMFuf7E/GXLJSXHoJIc
5nMRntB6ERpEb772jcMjy5lgVzdVcbgKzUBHjG/Xx0uo1bt1Lj3xS7qhWsvW3CmSrWmfqWJ9eRDz
0ZYQQ2IEW37j3wHAHHAJB4C1+n0qKPdn2fzUgARbRUYJlS84tH6q8HdaJU7D9/qY/fr9hePtyHnx
wu0qqr6ook/S5ptSrMf1uJfvEM1gWJNqLsZgajVVilK1PRYNtt2GFAElR0voBZ4LMVvzkEqc3Vsc
XpjkgWmJzp+qq6bk23HuL3ea+KwJDxlo3LzhOlCg99nrsO+fjtuWU4W71i+XZrjfto/GkNcJky1r
PMq0rQX4BdifSbIZoxrWxmOKvgE9YeHdkAK3nWGQrs+HYMOI3NcCMbMo5IwDo0TsTtK7R2tw7ZcV
9DGQY3wjrU0pJxzsvCAyuB7rOXjGLw76wk/nAF9lJaeA1iumH4dnnVljLwP5Kg9f+wLjkimkBa6P
sYwEJUoTv7+tonKaIqkbGN0y6fybEHkAk5MvaV8Yq71vWaCbT/eulJgvm4xWKwaR12atYm4/XIQ0
a4g4nLkbDS9lK0X9ePI9ahgRp57tX9+jG3jkICZYwlEbmSIm1emuZPoD6/eGN+ukde5CDWhiJv8T
swNFM5R5LtF6M/LAP+z6lA+EOuSPLr04Qcgq6k66I1awMXxOV57jNArLuSTa/+tbVkmi605pHdP4
UJQBPWBrFD2sXthwLAQplvI94x49L8jr+pwa5L2VhM5iHkqlhPrhauB760r53vaLJZ9kJjaxBmWt
+sR1YmdQJ5oHpteo4rcIq/Zt4YpRdGa/RSGqAGpRRX7kNRm699+RmGQzxWrXMacf14pt1njmQSz9
VXO8U0M6r8VuILf+PjWB3nzhbyOx4QesXFQuTIQCRW0eweA/1owZn91s0nfJvQ4IRD+9Bj2H8AVe
qYhlX1iJaxOZqFvhykorR62SiNju0RDVLGCUI4G+TfMB70qpt0sz86RI/BYeJVI8TWn4vsQEfkiL
iuAsXi606YwDwfCdBgsrdfpZtGDFv1FnlQdU/casIo6PuDTBF2mVqEhovd5lMfp5iLjKqeVDManR
wKl1+PMt8zaKGehCCrS9rVN3uR6yHs9SPYTio+1HKR4V89ZXp8JKakflujhoTy3EALGZYP8z7Twm
egHEmGzgs/Mf/cbNB0fSXw+Y9W4h/i4LmlP0+hSnOr5L3CQSQYwLq99bedcXfHp49EVVFnjk2PQa
arDsRLAij3zhx/m/WxJOwp/5uVsCa/S4tkvsneSlkehyoWumCk5281wlySRTWjbYq1nB0eu0cxwn
2lWW2DDPoRbkZtZYFzbQdjIY2Od27Mm4BT7bdBIHW87nJjZ+hJm7GKIIhuODb9UTVvZblLUeDhUC
MWhqhUcl5aXddSuUoj/uUfxa1iBRzB25WMIkeNeYo7GOXx7ISeolwdPSzg+8ppwbTVXtKx0n3caL
7QtS4zII8ZpH/c7OyKtzm2yd3eTm93Vkq+KMdH9BykzYwWmZdvfqx2a/zfHQ08TchqJhzbuwnWlp
lnK2v0io/EIw//tyEgk61NETIGyLG8s2UOCA1p+OR02NS0KWe2uTBmWEqu05X+rhuIro9fXFa1l+
AcKSaTVQ9So9drsCSkCeXrCichCu82yLcdGOa+Iea5Tb0eHQrrVNcLsJUQ4rFsEA/7PAUMPSQiJ8
WWvfXqK/Zd64QG0yeAga+OTu9F5uX/1wpbSKrmD7TMJvXvEej0hE8McEUOvB9fOUJ7kQxKehfPwV
UGCPMB6yk5ay55t1/A2PDTaK2X5JKD2sbI22+RfssZVoyxL81BhCQ5MZUFNjTXVowpPQI1A60A8Q
FIAaIs3ql5po1xMWDhLZRrrKc7nDrTEADMIe0e3JqZBq5+xUriUEaCYMFwmQ4+6kTAV/sRsmOsPa
1jq7BT9ISuKfetbAirpM0DSyCTxhcpgcFndGeMY5H2qiHRfkdK8k245dX77mbCBz6oUa7aG9tZGR
tZC04mxYPEp02KMZQuiMGI/Z520044LqXlAKScjkHrC1h/U83im1l0xFkkST9+6jDiSW/NekxXJg
EmB8Ncgt36gRIpd6SFvcAKvy8DleqECWk+KhBXnqVnAZJzO/7To/vQFUjvXguRIw21wgqqhfOBzS
fLcdNR2WfsuMXxGWXdMMSTy8s8gKX3JAWdqUyM7dEJIxKwfOkYDurwCs332Cwee/UwhtOgjC28Qv
3kCJjV+9BMDg48q3W+KK/5mRir+UzhQdSie3sUU4d2l9OmlQH0/XKnD2xPfR4ukw7Pm25lgx9YPZ
A71SWsC8fqfQe4Xi3FKdSg2oI6jax7GZ1HCci5KKexaEdZtpc3MvCRsGW7U3Nml05cQP3y1Mhw9S
fiBhK8HU3m1YUZMsTfFO7cKrCz1A2YzXSzFeYTgNP1vr2oTWT3HQ7YQTJj2srw5yxOGWI4ToT955
nmR7wtSckMjNvTP5QHpoQIZbVOvOpr3OM/1lLhfleegp3GGcCHtA9YmZRsmWBGcJCnHE7rZxashn
7BW6LIP3qQZSIjPv6lfLnXUQG1FcBHCAm4zNIacRYJAw/0FP3afKY4w80MLQRtiHJgQpZOSJXXpg
T5hZfYW8iPil1P6efYzDeN05StHTjzpkUmSCTVN9VjPD0z9T355Vzj3iSIY7VECwlF/ymRMYYLQ/
KlDtYErh0PykB0KhZCDobQfWXJeiCYjDaVzZ8iDJSPUNCRIOwFqxCDO4NUXZuxFZb70Sj+LwqHBT
laWQucrmxT5y87NQqh5rhYdArb4YdGd57dbJvWs3BR1Yyk8PIRlwUCfGRD/g3Dzgf/wdlUtxuzmc
jtR6SyvlPURB8K+pTonq7uErtfGfrdPJgJdRn1D7lWxufcJs82xahZXnLjFGZYwQQazallX6aebt
6BoPEdKVGik6u5Fao9UaU/BjkHsNA/K3XevvrwFzB7mN+SpWW41bmGHXdV6EkXjtwm37y9pPp0Dw
BEwjsxoCzZ0yps1fyxkTPvB5tTAV0ul4EUaJ9Oxfm1LY1BRl2xpegG3zJcajCDwn8oYnvvxV94Bv
vjg//uPp2GdgE+TFjrV/iHXuc+iYSZ6+2KOIGxxKGM8Q+Jw/mi8nHw2ohqzV/FVWkAlGBLGmc4hw
x/OwiituP4m+uqu+4FtYAqXiAsPBJe8I6BfOwYW9yatUIaCP//wjxKzAvgt/u23eOmQW9/b71Rwz
Fsj2KMwTmTJCD+g/OR0i6R+ztjHlDORi+ZvLAhFEngOg0WLMUGD+pV26bcVy//mJDe/TRt7g7UzX
8JZYi0KlZkJbsWYB3dlC4uv75dB72pM3sE+4HNW/V/N8yHiddZFPgCzm72H7BRd0L70s8N+XyIGz
Ouux193aC50L3LeoKN8ltjMhgEYzMyJfjYd6KgM3n51KZgFLmPU69GKu5gj4c7+uRrS6+vwDsZEG
jIa3zq+7rRkmPI460DPZW6Y4cetzILiHxDB7zc4jiC3MUyXjDITQ5cvcRwPbqYTlX2/9lMaE2K2f
gf5bu8xZkpwrjtugSWeRB134AHsHdgQMeBou3+T10Sy8SwRNyKAqnAD3M5WwbQCac7gZlrkOzlCK
YKQ2c8biPX4p/RMvJgb4WwEqXaySGEkBULboCOkTMjgYZYGerJGqGDDIXtQszw6KDGanyxhDVWf4
5Jcklc9ZkmBjtQkySGxzXy/C6kho2nOTUM9xOOZiGoBrA2A0w97DfZ1JPhkVTvXucFmLMjiG79Ns
aWP/hNTYWn5r83d+SZnrZdCiqzbBJsWkuMzRWWwka/UOrH9XKJKYkcsXM5EPrinPC1q+MHSidDt5
5iBfZq9o23cbpnN0nJKidAtr+dFcheMmtLDrB+uFZ32TIjLGDmbOhwoXF7oboWtyZhRX7+9+KubR
5HeRuxhqBHJSUj29uFhdMsCONyDFyJ1RQcA1nkNI0i1PJJozXG9svO0xWjJDxX5mjxFz7/XOtw8V
VlLyojoO0Gr/7dUbDJBOWWKf6p3rkzw9kjCp0hudbT+51ZvCUw5BgribUyw+eyPQwpGM2sWJkDuE
hh9hgZmvyCrCIVMIOx8UGuqmqoUYl/GeXnC1TlMSJZvCAQof4HIiYXhKU22REDif+umgARNmKufm
NWm+D/ETwBeOXJGJUNiy5NxFtV4GWxPiUaOe5vgjfAVf8899NerbYBZi5rlQxEpBZhZ8ughnE3m/
0LKGqu10ec7zNN30J4VldjFkkGxwInFm/FxdwQaLMBVnoATJG/bACvLh4KAJHWCCEqJmu4iEnFWH
aH6Y47cvcOIZ1XsBd3koj8DjdCCSw1IBg7EBRnTgbPAfelzxVuUthHZqP1t496eJmYp/X3VET9PB
qSVHtPZgMfoNe15IL5GDYkspq4Hz2IiA0Q5Lp2SBrgWgocrHpxQyw6nwOUypegAvEd4vJ2QcaS42
uGQF1QtJG32Y5bmryfYJ2tqQJdrorOSsOjFg/vCsjQKGBFF70OVh85bi8cvnYEQtd9D3Z+/I378o
Yi/R5Bed6IIue1zU4qXTDHDGpcikWCrdBaDNm3iXlhqFbxXBgNV/8o6jYpN+iSoOt97u0tUE96q3
lyGLo415yPqGjuhm9joUn/gXLSePq7lLsR3AoSqTe2Lv3TJwMFZpOqa/cY+E5Yuv9JKSXid3p4zT
9m+vFPJZEnlurO/tSDW5V6NUHsrB3zagiz0U82wml6G0Om4XClF5tcONC8u8shsWzNyhDYT6fhnQ
C0xoS6raI/O9NpA8B4CrJjuOJVfKGv5aEJcbz5ed+Ca4ZpaV+V4VB2jjPJiEDbnLZzIL+XAv0Ghz
DV08lWOeRhRvGTHqcbSryJnshB142s8YPFAaboRudqQINK3LhIfT67XVn4lJj1yL2iYJDFsAmcZZ
s9NlUTWuKfxdnDvW7rOkw00z/whyOCLY9KcCF9Cc3r0tVR081gUa8LLCietND32tYo8OCiOrtIv+
quYsKtowxTt4YE2LG3iyYWEKhf0drebrn7l2/RmmyvA3WRed7n5az6T5YhAePJ3lJNWCXu/lKkfw
ixTaPQCzDH07DUgEpFIvUVz1Cm6tXq09g8VIZTbIhu6hQ8gHjhP8CxiMnSdp8S86gWGmxyoq499Y
EMVO8eWyG6zIovizmeZMfi4wBROnXMs11V/7NK1yvS2/wUU0+3eHWvd6jAiuNXSQT2dmg0P1Iw7B
H1Ju8FcFv+KpLEOPUiFRarA8KIlIG/Leq16jT92rhdWHiN6KK77AcivyNF5NwjWfYbekC1ip0XCe
vrJSyKzlDsIb92wacIyG9DmX/SeWJI4bxZf+ucd/LZUkx5IjUhVJ098DLjIwMeOaMTHI8ipnYuRg
Qad/kB8zIudB94iZn9nMZUzfJnKyn6ZM4kdTuE1ZHq5+nRS6io6Jic8uGnDxxOOD7tw+gTRT1TXu
vl/XaEbrI9OxoTpBCGnr4TrGLJveiubTf2Muu9+/G6GpLClmEeX70EQXjoscUTCKCjdWKPFCtPNW
+Cw1w46IwiNuMZnD/W2Z5ljGsCrCfzSJ8DcDHA5Wf58OPDkjfoZYYqmFPb3rmHtMD4F2hPdXsQS4
OFjzwJptp8jBlfV89WthVeYn4piVZG5A47DzAc4bNyi0pxB/jl2Y1IEk7Gnta8gYdbOMOoQTdGwc
A7C2yKHaY9NXZ3UtdN318fAhfnzePeusmF1YDqYr1ySssXu3xeFz9ThrCti2XEaSgDLX83zVAqtk
Iny+OFvqvTY2WqtqUdKlsQ+GGqFIcj6AcXA3QQbObo5IK+7H4LiKaCLEWVB72Guqwrx+T1fBvXyi
uRk4LSH5A57rrFbUTVF/Jf5PqY1oRP1W3E/EmmslUYkqss7g0gDrIqc9p6/qRT0VzKn4JdQH7k8V
HOhvzDNnyzpvwfwz8HdQ56pu/FThdeLZ9ff3jKZ9PSyMIspbT1iYjRhgZ/OCUGyHZeiHEi9iTGk6
ZbGqukNU+NRWYVsfjiI6GS51ghlTVi2yvaMI3cZ8Lh2H64BdBQLnFmGajslGrevSX3KEnj0kHRB8
29fVAn+fgmHQoNUyZn3Pw/zApSyO04ogxFhC8XeA2ba4OrzDbO6wX5ib7s2aGr7qMpWYlYvVETPY
J9JV75OUPYQkwzTYs5fboBmDkzj9TGQxK91HcZ9+f4veBw3JpEcjWbSNFJ5JI3JFYqPbU5qWS2Eb
cPBjZhmDpgRbwuAad8RNEECsRhcP9KjXLOOvvHSwnRjflaxmyHHWfaO8HhBUUENTLL8l0xkyv0J0
cqjP1qffmpfkFgOjgblUWeRUoKkoz60AbWhgmbOsZkU8npqdKyRePEpsSaRZaslLW2T+7iLgkI+q
6WeEX05D5YSmOxmJBVeDG1hoNeiThj11sRN9l5q8TNBi5gifSwfTrxtWJH+S8glbnetLKjIAMe3r
KE2x8NOCJ23Pjx2JgOKfBFLIX78Uv3XmgISWOluXDjbm7OSLM59ygkxy1N56nYoht1B5eiUy2ThM
5n8ghkOO2O6849pakRSzAA/kHnMHr63acBqW5E+6qK0CqQI78/crujGcN1msTF+l0OyIGBNwvwpB
mmHKlPzE21wFH45s6QwG0VgTmOxe5jT/7t9tz3qmQ6PqbPpdqzYqoCSaMtwr6Rp/D59RgnkWj5/k
nKu1J7DqmUcIFUlKPjJxfatPIq13ha5ofYVf6SvuDhrFWGuCYxmaMafgdlalSdRC54aRLZz00IT0
wjia4aPFF/IVrkDE+NmykYKCvJNTIJ2lhiW7ziP4G6zz+OA23d76MHrbBC5i260PsBwqCK4ZIT5S
wgAgRTFbsrsmsHVJWpDMB78IstnGytd/m3ELDlOshEe19mvLy5zoPWT0RxvwSgo81q9a/iIuOjfK
qdUa4h7crZCEeDt6DjSqNDe9peFvj8tRVazWaA8HskEq9CVPQohi1FVk4HryPcgO0C4eDXuckITQ
sA5gSG5N/hWeiHlupTqszwEH9AnpdrPmQIDLzGCyQIgGV08UWnzZKjlV0XgmD2aFqf1GMJPBc8+R
XtzqbFimzeQfibkmourN/1lcgwaBdbEVHYVwxGNdKmlRySfAhwxZ5bDhdMfr8FSbsOruZjvVb7+f
hc7qSXK8BBySp9ok6JlAyrUy33zRuKMlBCSzVIRchJ4vVL4uIR3PQLuVAQG/uF1HwSc9R66GW89o
PPBmEV+dbOhuTeHSH/WWvQeRQeqPppp6U9VCazP76ZGSq0ZQTz50lRrNuoCvC8H1X/DVX6r52gI7
aSHtNSBYThNwiy/F6xRsNZStC5unJWNEzZdRGTK+HoU3A/Iw2Rna+Lz2ahS+KVXmWz3fvYbH6mzZ
ZLZebcgrdaPJroOG4Xx2Fx2URtU2kmcVPbegzMS9v9mK+OSdLoj0bz41xYeAlbh0J7E51IltA+0p
5uzsEvMuYqT/hTX89nAgExntO2jP8WlwWIPqwLm1E0ibfJCeX0543qnbyJmNTJ66o+imCbmqwYhF
fAczWnwHIR5AZsgNywtuLzPlG9UEo1/E9tsXZVhQ0ncDx+LluB9pbyEHGpHfiawIaiUyRsrH8fLx
FWiAiZVxa4W1sKWSBGMhzbyvwotO95mq0eHGbblmB40vRMcp0XBvD3ZFiEJ1Wqe3XrkCL6vsNQST
UZtIZxx8wTqc5RYJxDBooqEbHFG2v6xF6E/fgCDista24pANUPdgzEY+gz9CqFgkIKzW0Gx/UNLz
FS2DhDZL4aZQPXIuZaAmVZJIUbClvuywRX43WUXgGJjuKfesR0PmChnbtqiaPRNOJni65uyoPbLe
5dgeBMVWlWBjHi/hnJikh+KjLXeei2PUdoaYD+t+RIBazspvDUKt//Npihc1R+VaN8rBlaaingYh
vbwRGwNqHzx72d/6P9W0scmWGFVjegdjO9WRYV3PX5c4uKzYOT8+Hr+fs+RBPN2ad3KGJp2F7b8V
VdTcFrDUQHD0pk2Qn6Qru1K7tsG5cpbZDjU2CK56tkn0jixDkfiVpVtDCS/qCKaJZcBU4rwUZTvH
xuheEN1pXRy1Fd1jo6oDMh3MiuD3+ULTn2g4eaa0Okf0ZB+TmofeFTa8JpWiEcCHKoLoeOqCfUaA
fXGNcxh+YaAz9B5O8BuNrozAHKvT9oq1gOgxJCL0FoZThJuh1yBCmnTEB5EB5l7JsUdn73mxoSk9
0ATSlpHJYMdwhgzSmMXmPVZktbZ5VeFQBnlDiN5fMibJR14l3vv/KPDqgMNZyTgfPYPp1MmGJYjQ
jUmsKez0oGnTKVhQu1v4Hoo3hsFMAp4cb2kr3skphLcyMuEM+9EyXuRugWUWTed3i373YiG+qQYj
C2yil/R1bOV2AiI9GhCwZ9xhyq7YSAioML1DYmndlHzXCbOYZQ5/HD7agUTutaT4u82NlzsKf/VW
K+f9rehMdlVEEAqgyrz6UA35eZhQUuoqmEDOFq+L9wmhKqhtfgT7DT0u8VnyUzoxtCsTQQtp/cA7
kJANr5tSk0xKPPYLd5tuqJWBMsUEF/RlJqwDXVgB8SJQWt0mJqN9A419zUzWG2Kz5CMYeXJeDjbK
EQc7WUORXd2qxK2jl9vXL0t5M+7FXpgCSXnxumNvlsaGkhTAVWN+vOkLFoeE6Cj98HuCmTpGrSt0
OloDyNGhenqn5/xgz+cnJjyFF7muA19YO4bYv0nLW6YmKaYmGfc3z4DWLvbc0vsPibks5WQAjun2
+Uhm59WOJB/IlE4qb0cEwcL5//kkkbS0pAfiCQNuSqpDuusEyFjrc7NXcEgvLay10uPjRHt6m9Hd
PRNV6LHMriOqOthGqFRVGiQRB+feNGNToSWks/ZPF/7Snk3zdKTxc0hp7Mjlmk4hgfZaaZtkBUEX
g+ZJiCWIA8J6yw/RPEf1cYziZio5aV6wZRysohIwLkzoi7ejFas9tDEcbmC+/i6ife+T930j3vol
vyaCC2gxNfJYcqnZQulsYwpl+Npj7wxXukwKmmrSnvJsB+oMJCoNanzPGOsCIGY56cTmpYO0Pu6w
n5A51VrMbAFXNQ++qE/eUCCHmf86vmEsV64M1Ju2xNqRiH7TL//Yq0XAY//T75LVu0hOTw1c3AjK
r1Z2FTMlRdfPMyLEJesukbptVi1HTncYXLx6eL8Nas8+skLDZXMOA2zV34tLibHJ6oJwoSEMjfX2
qAZWaWgXg1qilnNkK6q8jKP90Usl5a7GBllqYOTpTN/vlOC5k9MUvPEwS2fp0iyB5U1/nQzFAZKN
Bp+GmPEs/q/ZX0WDy8+N6cb2PJCV/OJYZYr96+lQUyGKSzq3Vo0r2mS1SLJHSDI20mhH4dkiFieQ
Gxx7XwBmnDTi1lqwFLXVyyqM89ZBxeZhL4tq2mIGo+59+Qq1Ib0WDC81gogSCWJBT1SlgsCt/CfY
BFv8vabC463/qEIqDAjVr/uT+cm0FDvT2vnp7oeQh5IzYhdRqX/rNCwKVN+Q1AbjJQ2OMwtfrvWU
29lalOTpQMVdNiscZ/NpOY43x8kwAq+qSAKnli5rpL6/XvTkcr9fyuikAHPW8W4zNM/TPf0EhWUK
Uz5Nxb8+GYYCNWsRGA2HDE018ydWuMqFM2uVZmZxlfaMioJtCUr8X2SCet3SIUb86elW6JQ3JdFN
jm/iJeIQ4KmXOpojtWLoq6dzr2AMRqq/gWq2GfMtnWOTOrGAuRrU2Hm5G6MQjZ7U4q4W41ZeCalT
6nYkGaAfsbR4YA06J8wwl5PCK1qMQJZzZPXv2HlqD1RqqK1/4PJH2hR/m+HOUFXMbwrbkbKgE5cN
0n9FfJ8jxUcn24Ng2g6Q4IETXC2NUbUPav9YHSKKOpSTs5CrM2jnjA4n41ATurg8Bk7SYG/aYYBY
or8miGZzTaDP+w/eBujsjH8T5QESc/4gda0sHiWjk+mDGp4k8G4EMalEK+EslmggfcEN1DRStQW2
WRG8Wmi3v0i9UqFLAfH8BfgSW+5lxmzQSqvsDy+O6hBxBmWL1hD7FdkWJNlhmSnbxIEuDoTCKfvH
PNJBNobEmQCKflseft2Dcq9sFwfc01oh7DJ6Np3tZ0QVG8yCYOXtpd74x8o8oeRvB0sSRCmwSc75
TBhXMKFDuXw2s/XUQ2AXE4ffK3U55jbl5DfqBCcBAQFkpK3dsDVs0amcrTJew3QTwCO9Tq3oYVqG
FBumdQOieYQ1ey/MvKI12ht1ifxtnm5plWF4hanFbzSk3o2Qxp6WbkzU3w4GBqveRmFNFv0zvWjW
zbNojGrwa+0m7FCF1r6sl7qciADy2PRtLipQ0vHMmto4kYlginTlZZdDhIN8j9uj0kCrW4301OJ6
cr4GkeTUKiIvxl3NDqNOu6HkkRS1HXf0O4j2y4P3WHnbdlcHI67PQMx4pYLzGvsgQ+WBP3hxdnP9
4hjuSFeVjqypdCMHQ5jTVSYMK5QQmniMHYasu2hpvylH/wshA8obmt7hL/WnIsx8pYk+Gd4+dIYN
ADQnHLnUrHLx2DS2VLkVn8ZHVa1Q/9dXVxNNTIXRpNNCIRr2TblJlg+bEfEMNkbWNMTd/OZ/REl0
Yg6z/CqIS/eGj/YBjRt1XM0T0sfszgtyYjY5Dj81BPm3/3eY2MI1HIkRSaH6UugPh/SYYcRgNlcU
mcFhBSzzmknG9wea0fwu9AEaNiQAfIlXiXGsAVNav0+ZbKndbyqseEvj0Jjc6CyQufL4eNP+zFEz
dQr+/b2IF/PzIyy2zckKAsQHfKpWw9PYM4+dQUzPg5Xc177LeC9JskZFQIKgvolxmXxydNvHsNaY
v86fvfyFBVext5lkkD0ng16LONWv8QNrpqsMbNuMMVdqJqMltqv0pvyT6mh9sgbye8kcxw7+aEbt
w4jW7VwkdwF9ujt9bkKzPdxJYoRHm8U6MgwfaLJ7G1RC31mSlq6Ol8pXwrFzXPncPk66y3/f7O/s
wL1thYqFskMZlP5US74YFbvzPAvvJUXR950Q/zfMDpr1Z9x/utCn7ZgNalUetp+1T8+5US9GGgaO
PAstnBqjAXgf3w0K+SyOEVSnSIM3KGMLdXMHoCkbdM2rDRXxVMU/qWxupzs9JqJkcAru1UMewq+G
MQJMGhMZ0xWIvKvyw4IhDN1o1lotnTq2dtV8p9v7TEot9GV32AKAe+6R6aAfxoH/y0B/cPodf22s
coN02rWYs3KiIHm+3PGVR+mWV7TMGGxb4xAjpfAjrUUo4gkH9rOpAxBXLugXLKIjNasVdq+XaIA1
RuuPKgEsISIzRfel2s+HwVS0fI0CQCriSgR+UHoz+voSYhHM1kmg2RNdNjNu+O/yuVDWRgVHGB7D
ssbB88eTsXFKjb1FHoh6T9bxZdF59emR6stihkWy9ph+AlDyPSGP/HamZV5fbJt9q0FsuYK9YKz/
4NR7WuHvBgodRxVucdc8/wDj1k8Vk92JffcqF9ujc3NbVgbZ8kOceAvPDjIWisQOnarKjRL/lTGn
xciBmdeHHUpzYjm79mFvfqnZEYS47t8a+r5a4dIHsL01qFnBgcvqEL/e0J1970uaQbg3d7w3L2H9
+Ai57fMU3UFaLEL3IzL9j8hinXYmQv4ZBmeyljF0M2kQookDGY0TdhpwqQue+GA3UapraFg7RlGb
RdeKYDBsEdpEHXa9RmLzRtiawX9XSiE+RyxSb2IS5n/CfkKib2nWJUG82j2XTcEQJIOGHhJPXpSs
G+o3ZAaJBuIFcI43s4P+WmFAt/TP+S8stvNkgyclLD3PklgekRT8be895stV0yvlb8LBXfYcBfOM
1TsMwfP8RwCqmsNnCEmB3MwBfMDgzXgjyGjZg104+qzkhAAjd6u9J38Yym1KFP5BUSnkCA9JjtYG
0/bppURySAXpDD5Ax4rfDRvRIi2rD6EB+UG5VAmvwHYkSlFOasVx7asDDNsZsJU1maLXD2qLs/Fe
BZf6mfNSelGi+UBM3PEopuwOf0sQm480pMliT8JGPGMMlLBrbqk4C14BI+X1amPoSeQdtlJ7MT4N
DIDIP5e/QFONwZbL+Q5FJr/fmxGWHew/NLcVVmlXunfrvNHMguhP0+d0f5izs0AJmHSnLfNd+g63
YjKtrXTkb1IO/9rGOnljFWLvIIhQ8ex6GswzKBcsvRMm+Kky676GiEifyKlJkD9cEs521T5EpMCv
UEhFZWuhO4ltr4MKMAXkRuXaTY2sBLRUiSwhhgRetfJ8YB8K3dfuA1XM0GODZ433mRGpOn4z7p5z
5e1fnNS2de4E+bISaLRyz104KQrxD/03IcoG3oQXiYnc7HgGeNnut1uaqmPTt08cGlzBbTuD4+6h
PwezPZHirWHK8CPU3wCzmrr0SttcIOxYgctlkJtWDRotkBKPhNwdjjjDB0TxY7I2a8g9YBdQ5ZEU
cyyP6HAjYzxPKjqGcNDihINx8ClE82mzs4UGhPRJSTts6VYbQM6InIAjElMW/CdcBG4QIi8oVbU9
8gYLjVKbKwqW3RdfZgrqCsSg97EwOyF/D47D7YRs9YDVJpR8hSoaXbYRscYDr6W+MHp0yOlIa1Ub
scJPEyKKsJDKVigtRvGqX+RtWekPF0T891MSdq8yhc57cE06aT2vBBpu468ZCag+fyHw7h2JRb94
I0AQVu9u39FRp4+FrpQfvDOgsclRilJ2L3vSqJ6CXsqWxzmuIqBYXyEJiyS4vZ5GvP/a94sO3KDk
MUdiyaL/7cqGguO4TQS1M1UY5etrhVFooMMpynyWbOMTcqx24FFzyOB/QVa4sItPn1XPcohFOuBd
t5Jnoj9XYHmKADTfJr4v0TEyDWiutqL1/5jx2LsQBvCN0oFpemBY+GnFLl2dsjHTALi0B6uxj2xP
nWsT/nMWXw6wmFRYwpCAaJ6oCF23QvXHow+j+Pa1WEZVaKVaulp4Y3QP7cmrXHB58QdEAZUu9eay
98eRhTdqbtrFsffZtgB7XsA6na1zTPklksTGuNCTfQ07dBxpsk/I5g0FCOg2ap9n4iwuuEx9jp4J
BhkHhTYfDQGhniRpnZ1BvA86ff2Gf/0eTYvmujhnS25ZuGbv8PpiGf1wBmcj9Tm9lK06YlGyl72I
yeZj9gWl0YldR8aV27T6K9epeF5qzuIOMnOXNffCphSD/VDD/tYDku4yC2V513X6V/DNhUaUGafZ
RBFCORTEMV1q72Qa6TFGngPiqeOE158VBVkHXvbn0Q699cNXFZammovqmpNumPloyNOhaZ+Z0A+D
27nT5dactmiIdhCG/clPTcIGDyyfYzubqDNjfTvi9PaB+vXgikOPZdf1TWDVcwY0t+EQ6xM8/y0Q
E6MckyjZXUKRAz+Y1G8ZdiV3V9+P5vPrlzGdCXFLqskJnXYG5FGT2/LE3cmD4yEKk+2osjl4EGKi
zDzbDr2q0lNgoxXJKxAvkUPYYfsfLZ31hZOMZXufetr9xSX55x+kx36bvEZl9+bJWyqKiZSPj6zu
Bk7Ck1ebcniIiq8aRXmHoCqgw7EFuPUOP+TdR6lp/Ekmu/U7pYigDDWAOrdaffvwIlH8q8Jtip2E
h7jyVxnekRS6iGIu6laz0KJQeCP+dAH0+VTJMAdVlGQ1FHocQBm+5qa2OHiA4CaGDfkBpcy7tWo+
NonrOQXgEOBL6uCNe1ICppzt2ecu0vyyJJKt6Mo15Ln+vQTHqgFhyXfYn7Ib2kY4JV9BxNlx0LRi
CJIvBKJEUYg+8bp9GX1PGvb2t8c47uPzcZosQGt9QFDj23JdPGzmQcBkzioxsPV9JE5n4gKamVAc
ZnKDp46/SCgLDdX/CxqZsW872dx7pcIno1hF0UvB7woGAhhq+wfW6+8/cOlnQhg+N8puQhjoGoDr
kIIzLXraTIuC6PyEzeT/T3C7NS4efFDraYW43KyyZRNJ6YVxuAS+sPq/UcwOP/GFn1mXh5oa2yjU
g9tLUlkgkPpEA7L2bxcDWnP+xv+fuIGcfGG37HY+mmgaEAERuMQBnXXO4K4UJRa0SlxScy0rgyOP
oKCm/yhp+ERMjN0PPhRAz3WyCfIt5ZOP/e5pvSyyfub1xteKG5Jr3kwunMyyPI4YBEeXvz4Vg3IW
rsLVgDR+t/mgI/Tzbe0gPHBoLr+8bD33iG2+kSkN3HDbT3QAKw9VndQDh/a0tUC52PSe7TNa2Iuo
ypZIYIb8N/62GsdGvSg3xwarzXmKeXhheNisUn0SvYhUOVBZjf9P9DT09krRsnAlZoD3bGTYxt6h
bMS3PME/W7ykGBHKQki9aHAIMFvnBTVRPrfNGZFpAmHs291WS8ekrBTUNS4AbclnKrxtMJ1FenXl
zIy5zIcFC5BNWKWGlX9fKfAFSm5A2D2rN/VPWj2erFbnijv7jgwQ5KrqK2lCpYLCNd6/XqXUf0F6
iUlh3RRVk6rFYBN1rgPfhhXoHwVZOeE6W8r57DEdMk2AkWJuPXQvysb2EJ44Z+R3MTT8JtWnlXHB
ZtWvd69dhkep2MQzFoofpBu1hfJ79g4p4MVcxmnLQAILELkqzR3XIau43ERAY2riyh9JNPA/MFCA
K/iAQz1mdekhKygSnxd4ExKvaGql+MCE3fkzDu5fzJNYvtsJ315wCBURZtKECoxAH8efo6GiPLcc
ErdSC31vSDtqXuqNvKGSiuxmTGfP+Jb7a+0chvRhD+GOLLfHTSh+HOtNM5EY1yIF/L6SH+9SvNmz
OvhE+yyFWCjAiHH8uIvYpzPVlBdQkFtPWTZHRJLzHwgLn0MhPcZ7yLyyd5BPonH019W/fQNyY6Ga
ZOGeYd3BXxYJhwI87UsRlzSGANQ6GjUSq/upvD/4f3Cv7eawET0OHrhwUu9yJRvDygFL9pE96rw2
6h1WDEQvrryLyHxeIAIsjYCObfgJ6AZJIbyBpGjopDhPVO0O9yurgVlHFoH26ODwtdlgerj9hlNP
3hq7gQOoncMayU8p7r3cPDa0y2MCU/4TnOJY6XUFLcsk54GcompIVVDVUh2EqG3+SUMQcdWfMW41
GLrpzECaxsM1LLlmrttjrj/b70uW6T3xI/NQ5FGvBgWLrk5HMd2PB7Lnfd015xHjk/K+0oQk0d+r
NC2nZjwT1tuCUZDErF07JHmS67DPVkuwD/bJ71W1y25FB0ZcD9fzo5IpS8XzX5CTPCNRTTFuYDPe
nfXRArZD8qZOjIou8yuVnoKG4hkAGM0FJb/BWyLR2RR0Ow8q03FFiOw78PkcHv5p7TwtEy9C0aJS
Iio46o2FAavYBl0jmGXU+WTbOB33YDYJSoEJBEgQ51LV69LQj5ag+pzyadDvqZllQ5sE0auyyy7f
rDCfWTgFqL6sEIyaz/fwpK8HT7mmrL7SnXG/T6ATtAmfVTRA/8NibTbvlKVtJ5xpqQml6s+DmbSD
8zMGSWTWgNzS7a+SH5TDzmHxKQ6pSzfsIcP7LFBXOdnnRrYh8jZMkPBARnptvfElSdQcC2H3VRIF
TIdFReMjK/c7ycdzzqdbChwEh9LmZwnv5yZ7GY/OzHUER9GQCcUUsWqh1TkOHFu6eakv09h5dCjR
V4PtAJ//tKH/rOzMkG59SpsmxFVCXDnuKxFfUrC7U7srxUMv/fQ4c4Wuxj9Ciwpu5FPLCaCaZPlC
TNdld7uRJCLWTxayNOt+NK2SCUUDMyHiXMseG91Qx+csUMzn8L5skXyelceg5cZLTOjjIztb6MDO
9cQnU3TIEZO/9wP2AlRWer61hEI4Zebn4if6reytDafz03t3EodX90Rll5V4eiCsivcIIzSYyK1s
Kxe7hOoVuHKdEGgmKXFH+qanby7Lf38V5+/GkUxSIKXL2GCKKfiN0BKMN0ChdSeRtP6/LRmd4q7o
2NSrTWPQCySWfAkVrJuncw8YIwnKk/JgeolbyJwnNDdwQsuNhDEScJy/6+3lAgkay3nt+KY+PGj7
IgjCiStkhbzTsL1bxxBXXVQkGpbEyH6OXZHl3cGX9MvhViaxgthmBPoLKXDJiIKrZvDBE55Uyoc0
gJE8woRBgJRGZzdB+FbvskFctssfQb6yT/qGLvxYOfb+GvN6RBodYXBOq3OJXpK+EbczPG+kqaND
BWhp5a/ZB4FOM7M3o6htT4isfpbU5gtDp+JTK4BL393w8mCz58hJGJLchdbcIy232lCd7tpOLNNK
XrqMiV3SZEaOZyag2nYB9JpAVKkaPf6i42vih0CTGn/kmh5VvJ4PeVk6bWqxZ4DJQeouYZ7J7ZWc
XIfg8Rn7Rq99njFEGwlOBMCb84MLMgLwdCWefIapQu2VOb7o1QTrdaj7I9unc1GIAIOI57kXtw8j
JBt7gTo6hFeGvVBOyEUb0NrLbHMpgANTtFlB7R9ANVvg3zGGx0WHxZvmlcxRVnfjZLphGsTX1GaU
p1oGe/GrIcKYoXLLNnhcedSOS2UekNzn+VvPi2fw6P4ULIY2JaB25pYUiWTbApJZWteaO3fOP9+6
Bg6pDjhjMWB4CCV+NwLsrKzU5r5QooQh9bFM3iLZHLK0i2O54CyBEOErxfOQRwDj6hNxIXnp1zZZ
qNvzv4GhUiMxFx03Lr1uLcHI/O7BDmJWDUK52po3Pd61FNTZcpxTZJ1N4xUmDAMrmX/I/pGofj5Q
RNpv2K07nsWQEaD6zPSBNwf1Fq2AFM/BiZnB65qFMdKFppoXwwXZt05odanLHjLEGHjg2UTmYt7/
mRZP74fSpDEH5b3LTM5pgErrO8IhRib2vELIYzqIRqO+tf/QCVRm6mmwWd2qtfso6LBckBGijbKr
TQgfjzF+INB1905mvJRdsxpQI7s7zjfGYk3RlMou1TYtunIulav7h3pnKb8HTVFx7cKsWiWUCyci
esulWbZ2N+MlMHz+GaBomO5zjBv+IW/n+ZiHZ5B8TFrOSdg5/0OHoYXEXnvVa1TAK/nOq1MaemgE
rO8JaeoJEH2f9OQd/HPs9tHPLZ319DIWZ6gdpWwR1gzpqwoGrGoYMxCtEaApyOsYIYepTX7OBWoD
D4WCQH/toBPiPZqdRlyWeAwmoNccXO/NcdEYlv4c/H7fLBWv9UVphMhRzvI231FTyiI8xFtOTK6H
UkzCvcnFqRlebdiGxCQQFaYbrkTuWgauV6of/Rh5nKQlzxEYoE74qGlBPeZfjSupQNRmf4nQ08uS
j9Xe9baZ/bXILeUPGVGGf32AOuBO37sbHVJSbob9/5JmiUwBZbmV/6qIfX5Dgb6DXqm5G6n9a06L
gC7Ez1wD9fLb4a8CCXrYlW7H2oTw+GribM8natH1+tESiUtc8wu2Hl47DbTHkGWanxGUZx235MmB
rRaku8YtniCUqqIk3OJ/G9kZuQYVeFp37gkWc9p+oZ/O+9105FsXQpJjcyq/oNuctaOHq4dg4CDv
j1PewUThr8piePYiMCQLLhMGe97BmtyYDOM4qkiOPHG/3G7+9CwALdJcA+WdEytTash7OjqxbDo1
gH9wKnNyECHqx+vTTVOEK9oqpblhc2aYDGpd5CXsqgcvl+L91I4PuDPSuG14E1zO6iJvZzR1BQDa
mPPmAtAZXbv9opmaqII+OFKGuCsIhX/e4msFgEmZA33h9NYMeHyiTny2SUYZzikphRN1oGmcYkzn
B7OieFolyq/ihj5xX/ngyAXMeOy9J1dP3vdJMT9i3hpU0xuMO4eTaYxmjiYAHA8VlezK88jDtk/5
zlS4P0Ny04aJKPgJgpVjw8kXsfIMbA+WmmwUpJRd+VO78hNBaSN1z/oE9EsNCjwtfiBqfDtfh/lA
3+e4GK7CusP5n6m+437HGrAzmYbqsXjja8mJ6jUQpkbQYglUTJojpKAQrnWlbiIWr3kG4sgsBkNV
yys9H+tzqtFaL6jbvqFtzWr5RQnimaSu0ahXLXmeJZ21jWP9ziw1LfdBKezx6rDhMWsttPcQg2X4
N8To3qs+2n7OTjXyOzZKUVhss2jYF2Ta/05L60WqRLMiYAoOpq4zOcxT51y+XACoOX1z0ZawT6jO
PYEugSQh95QREjdliGf+NaOvmIlqeIz1FkC1xct/q88DAx4a0h1fEL57qtTtYMBmgJap7YcJN92V
Dn0sFRPoLNltxP87bRSHeVzA6QjqZ+59E0TgH3EZyS2RIvgohS3wHHVQ8IES6lvD0JI6U7cP+1cP
eWHYoo0YVhgFqcTy25xRJB7d3yIsEDIGvL0jhqcrrzS2i+smDtsFy6MbQtvUEmK0oEzaZdQQgOkJ
T4WdgbjLicM4/8UZZ/ucPz0XWb0K1PPJ/nfnQHN/Cg6g6D+iIJWJiaenthtg6PAiJqI6jRa1UDtB
z1b+dmpjbqEHvPw+H86VmjDGqL1i/pzCWXoJ95Vz8Aml3kdzEhlGt/x8RyLvHrL2YFXl4QC/wN/d
q+2Kj1NrDyANq4UtXRraubJF8Z3LVnphfr1ZGWE47p0GDiKFozD6GG9O3Rl04F7HyVsaD/nzTyQs
qg+lcdWW383X/kQe+EXPteJQ1hb11/GVp368P7HE6oq1PLok6uHtrT/qcW+6+to5YYLwhZvybD5n
EKnLNdnb2rY2cGEFdnSMsJa3YaxO2Dx1QpTslZNAyL//lnfICz15LbOZXa482k8Tu3UsQ9u8e5U/
c8MGL0/emRkxJ0Hzi3cW7XBUbt4c3qJawnR8D7MQNnbNoHts5KYhOI60GYFcbYLm+W/5ovtpXvFp
v6WUO5XbsIi4NJfJbiHSvG0gwfae9Pycw54NXccJciCiagTrcf9r4vvTCZ8DlJwaAwmXUOjr1Piu
3u848whiKp04C6apyEeioJ9iJiT3pQ8BilfvzPxbGNJYsmnAY9VL6XNVvYYGFqF8NiJc1eoOE0BY
pjTT21M8zixfEDc3Sk23GloAmUoD1SvF6ByNFm7iWR5rpXxeEsu2UfQR+TKG+sjbaqMGJsyv/yUQ
couJUOpeY20ExCa85PemWhwBa8VWYJyoQ57Xs43cQyM99euLZPqz3EOgitxK7k+2RL5bfGhDzxdb
KnC3qokmJzZKIt8VShyhqFYxb/hCIiVq7TWH9QPq+9tbvT8SgK4GnujIkpf6VqIYUMZymKXV987V
pTbEO45T+ijpJmOSVHLdxCZAl8bWPTVIWtBhE016kqMDmXu4xzIa48NokWLWCfTm5gejbdU95s/g
comQ4h3dlLK5n6MrJpP7LiqhxoWpth5AF95x7l9nAsFNcpA5VaxBc8ETabSsDNfnQa31Yj+TIYCN
CNakA/hvq3jaUTGbDIdFuaScres2ElDywCIINrwX0PGtpKxFbbisyfGFxfNqnXEQl7PVzlIN1GDR
Jn8+grTIGYu7Hctzsox0pBPr6NJ9pxtYP++VEm3bPAt2wSjEB+cl+ScSpwZiq6wrBmOz5ECc7wWu
J7T9BCkhsPO31+Ay8u8AOkjux2vXyWsxvel02gwi/tP6S2SZFLWcQLaj8e/7hReRO6F8EOQ7ANAI
OZaxFfgqXbee4XgOnq3UrEivgBqIx/YYrMA/QYdhbUHVXhr/rOYoW3AA39EvpwGzr6rJvhA1SOFm
hUxYMZ2iVmxYM6ZBuSxzqThNPvPZj9F0NvvrF4KvSbCbJkNK4LgXYhymgMmnXPdqJbcmIuLrl6nQ
7VhlamOzi63gUer6uhZqdYDFe9geMicOgYDf3ea/l/r0dfI6XCK8YDtZZ+kzs0+bmwvSi6X0ur/S
Qsi/VslXvYsz3VdekZ9V3WbmQyltY7h3Y5PwAEkCAk0UbF+Z+8LWLS4dNlqZJS5eS7iamluVbnbT
u6MqwobY2ZwnNu1I3qec/r7sroIaVemmpgx761iWb77nu2if6rbp3p1Lw4qoZcZt0RsiPfvoIlkO
ISy+2RFWfFd/A/vu/5o7yD5aFFkn+FfFY3Cja1kluM+CXznosUX2a+9+gI6ID/BFO+je/e6pR4Iw
h1OBuTOf5KTjYg9kSCk+iGTnXkxnk6pL0hpZOs18nv0UwpMKZZZercKm0rScw4Wi5CX7S9i9b6FM
l6nE5dPGqb2L9ZCgrrXPKfKxHea+0PzeuBFBW+ci2pZOPKvQAby+IJE9DO2QZze1wOjdSP21fZ78
JSrVSwLUBFkvbKeQ4m5yf4uQzgGRd27kRw2drsXdtN1egji0qIpz0O3AbPWl+JkIDO7nrbGNttNY
88XLeuOzhy9v1nU72N2Q+xPIxebBP7kYvObgIJYZJpongh5mM9Dr0hZr0et3y2mTkazu9nPlJcdi
BFj2GKQIFtNsYY75Do3yibfJMn4BG9fqfLgYLzaTxN+Vs4yT9oiZ9GiLPcxTEkZ9U2RVR+YkCSXw
i2ShzUgAawaHSKtzc3y2DnZ9NyQY7tIuxbtoHGm8zHCHJQgsxvlSv3yEo61/2sSRbN7J+M1zT/6d
Ylp4piiC8nmzQtekg+YJ0Nz8VH1cQGuHrKxJW+OYN1qetFe9FUPgS9YZgYNCvlaYSIrgwbiH0i6v
IliVE16iTaozG992ci6mcrQbGsseJkvYUaze3J0pbcRNJzNEPRGaLIyQFetLE1qXaRb0DnUEhbvI
AOySjmIbBwMg2lCDKMBli/RvZz4P0pcySCnbWI9VwPHH47MVLmC8jpLtkjn1cIkhr6YHXTHHfd5N
2qqQdjYjI4FVkwijmlLe1zLcyk79e+Iw0obaNjOnugvQwLRkejEgXfaIyfC75J9XK2mhy5eSlRS8
mNkoEJva0/KGFZVCcykYf0MJzkUZ/BEpFajMYP5P6k3f8PcNLxpL/bklb82ewY9LaaUVPsnL4LX+
yZRF8tCadYxwp75Q4SirZmFKwJO8Mjz//gjoafv75i/DHoXFPpSxZiBLGt8+MXVsyW32DHPIKH5Q
aJZmEmDJzLiuEaYorP8cISRYVQRcXUv7n9BL64667EARC5eTfQjpHQ2DIXpK8it2Yd2al4/br9tD
uNPBFLc2Semme8bvLCoil752htL/Q+smghDun887MCYU3Kt2WEwkuZW4YtoYCZKp8YWJfz3MBmb2
/BcdzJZ5HWa8Q1aMjI6aRDx8qYqHu9uzOYcK3nXLn1U+zew5VxChpT/ySaE4C4ZQm5sipkpt9L88
D6g3sXdfm3xl2ozgUVGBDuHwGS8TJGAIN0iPkpGUAEQS7hbgMIVUy5tAherw4cGf6etUGnfkpPZm
VZLNqeJdrllKpHr8oh+UsCUhzzXtFx9OC5VluMsJZHT9VcqZElvjdi3AYw+k0cokkjJ3FlId7ZmW
Ddhc3u+D7q9XUd0xgDmWUwGy+1FU3gLViJQreAtCzAZZ05Te1KowVQYzYB1vl6ln5or/nD508T5J
awrmq4oRztq3jngMEJEIh6LgHlH+usxm2KRzSPzRQVkoXc+7n7aDUMgwF1wH7bZG9Jhg42mAMlca
lw9XI8+O33RiX7JR+l01XkVBrqZvhePGh/uaz1lZn7EY+djMgZ2aoPdxA+I8aufMDeE4eHMteiNv
gO/ys8yT29xLH8jq3w92SbrzM2Ol6RBGWlr+SDc9SH6PH6/m9ppqLwfvJwXigvZhBENtuiwCqPsH
Y+AfVsxXspI8AHe+LyFThAvwD2FUCOu6IJptF/KZrA4/Rn7AQqFl3lq+JrMKe24OqWs5Q1aYFAbM
169r2jqV8XJZLLL3PoRKd2aF3AwvH2dwlvtNL1Qpk5SP51234379pXLcq+9jJUIgpU1PkUgFcnrb
HPaW8McmhNDxxpO1GdaK9MzkJHvcIHOrn2jRwzWOQrdaQYiR3QYOPYqJpbcx/IHBUespa+N7Wm/P
8SkrgGDEXMPXsGxB2CV+/X6JJ6Pk0i7gjJt2LUX6xOTb1hL58xVPOuunfAy/iE9/QBox9bztx7LZ
CR/NWDEzovQW4P+21hGJTpzvNi1oCS8M41JSp37Y35NtH+0lrkzNm5wtMyhyutlLLSlXUdb8N/gA
WHAOZpD/WsLRvLfpeDB9S1hJc8Rzi/jpm2xrggrXKL+A628LVHqvPF8wL/2C8Hxb0oLEQzzqS2K7
H84SRfZAd/GmEP1U/nH1pWC95H1J5SsGK7Ec48HT17nTVtVgy6XkpfvT5tfxAaQDD/tQI4Mk+i5r
+efq4tYVIHV98whYkVa9MyJoJEqRbADoebDLeynI2GHwAVQabA9gJKgVANQM6BxsyhA9IUZh5/H6
RGFn4FZnrKz1zY10NSFsMzKUpHPW0qy/UWe+bW3G0aSHtJZEarEh4y7gHp1v3J3vHNK6dD8mUaAM
MYygEbvPgtlKG+NeqAaqIAHbat1Zez0pCnmMfsVbl6zuqbEG1h7AUSLM5w1RHfgjiFMOG80km09/
v97DJhzfCXbKH8Wi6u0Lr+L0vWwypjzf9J9KZtmydrpOeft8KtaA8mgYlwbmTDYb+jPLLWykcLiF
IwoUxgfiVm2aJLJX9Da5uVlAQ5KqfuKV2fEkRSInubOSWrXOWzs5QeuJbVXumcF78d/bQ+D/35DY
GAZKIeAtRsnEb0jqBDJjyuw+G7HRoeZdFmQoImd01CUWei72Bx9t2UbInodBINnw/6rNlWHcTJ6q
TFlC2LKcc3BNX3Jdmql7/42lxFKqtaRNcrmMT03NErbi4StVIV/1Ehc9ACSFEVNFmBKCjeLwPtQV
yPDgxBqmzD+ksH629MkVNBePxpHWdJDjqD1F4epNP2m8oLcNnffuSLrZr9RYQQswmnBOroVhEVBF
3rmFN7lc9Shn4Ef0GXb3j5gmRKgJ1eAnWhWZPKJnf2PFOPb8+0180KyFIR6004Q1wzZNSfa52543
6T/kDG9JMUldPNY1N+74f0yhGirwcAKwO29t2ZLBlKm0cTMwSZe2/0F8xCzV/r5aRRrg0aqFBvDV
60Je5dDmofBf2o54jviW7OBnLY8gPY+sx9OKsmlv13vL+kVp2ZbFeCOtk8aIMEPqM/zXa8TRo7RW
u7mhpxa2aCackT2uiHjAI0jiAsYFhaDKnQ2GnIizR4f5vxoZhCovS4uUfxtCs3Ep12tO8vCcOL/B
Ef5yms61GgHkv9HdE8/7JbtlAwJnPgzv7K/DgejR7bhzgdSUjYLrAV5zD9IJz38ha0Y0pLacBjQp
W0BHH+MDL9zJDx1TImyZr9gyl4pt4xox7En6DdDonpiaXs9yhCvy6n/AZCjM3xf/RvCcuEVH4Tbx
kai2oINeu1zzUxe4LXxaVMjKN7mY2hwNb+TUcJWTXEpLjPG+0E9/x5h5r1bZGKHndxJ5A0h0OLNP
tAGHw7sl87GetTfS7dG+lnKUdJDbL+5VP++HaKkL6B4A5NYwg709I+qD8PHtHSicFAwJTq5T4zDI
OEHhj1mbhY/cb4CxM1YFqqWVA6pTb2ybW8dHFAtsaKkNu0ShivOt5ujlRHPusGgoz5cnnI2W/R1s
L6ePPEJGT0kbu2fEChO7rZqWRvt0y65U9neiTrrAVMDjq3nH91mcjL4qdlHj3e4h4onrXOuQz5BN
sjp5237RldPiBlFgBgxhAOGPjRl+LI5WRxDyZTzVj538bn9HlzcbadequAZcnDLEXUytWF1jcBE/
qyHx/7OI4BDqqVHqEFnLTTRbtdWcmcBw2Su78Vx58/v7+a9yfcl1/hX4FlAmIWGMy1tkfrGNL7mw
xYTY7bOSSlRoV5Yh/ukDlQ5eFoGz6M9jSSwUBuCqWETkJBdTyhIgdRX+tqdZ/rawFuflSQvTHNt4
neLpt7HZiuHO7gOqArXE6Z1DcBLylKcBxfCBfK2Ie52l5Noc4B4K7qI8E0SAxR/iMAxtV8pFc9H+
Cj7/FfPIKRR3mQr8yyo3tGzA0PQJ9aiLECrD+kkYTAroGgmRHa0H8dmUfa+QZqhl1m3cLakbzA1Z
jNTTtk/tESXUnTtYOSOyWAHWqcNgxjtJj+7KNUSzKpU79esNJPFoLz0gTcFZTPFEEC/T9rD9NoU+
T71WL8lPztU6OgTl+8wD1Z5iiDXO1d/uye6jYJ2DUZP8ZlLGii7rXwSuDT6i/Zn/+cuVmvPtfT1U
Ak+gh7dOlCMelWbrObLwUZT+zHp1Zxbj+HWY5ZH+ly/B50Gpy0XJJnN3/J6WEji4QA+QWd/TLz8z
qvD8ky/KKuL0ZM2Gq3ImJrbNIasMSbLJXSi/aTZJ+MfCiHUiksYHAzZiv7dk4TsClx3yJdHUVMWR
0IzUho2PnlZcUoWHuhS1VQFxJ045P68JDTgU05QYRTr8kQnw/Jlw2/5ISTBmh2Dc9E0gx5swlr4B
RtOOkXc8e6VLi7EWT2EzKJbX7zuFlFuEpdUHh7uAdEEYZrMy24eNrL+l14gQSZlHAawTqpHU94h0
7wYJunGSRsulNGb1KtorbSf4l9XVTERSvmWIdSRs9zJ0ViXQbzFBDC2cFKRmej+/5EodpnHGuTbP
NXDjXAuAMaHux7Y37ioWKzA+OdOXDlTBgrrgSiAn62wtwWPZCraXlUgWe2f93FlfC7uV9lCiNgGg
QqUkLv01lKywTJ33S/N34x65W+bUtJ4hCHlLYi/5NyF0JyQzbYBdtebMt6JgUjJ9B79ZR0ZcF0D8
arCYxbDw7Vdi64dINCZ8J+pNuXOlL2EwUnvsFo85bQEOqao9ECrORLeDtDamc/lgW2pPRj/BPthM
Tj+nvpcE9yhy4D0e1axPgRk600OgJC+4fkGaYUFT0jtPCkB5li6ObxwMY862Vy6UBpP26lb5Y4x0
aOjpjZsha3ry1lfgemRzx3pmQI1PjOtaA6lPepEAZJ0e3cbvhQXqk3CimItJMssUBQu/8kSBCsBH
qMlN17yhV1KhJpHCG0WN55UiF3ZpKrcoLbA+p42p28pgVeJkIX8HT5N/GSS7TDokNEKPASYtdHTN
zKfiAJ9MLxHCYdF0f5imCZbKb7oKve3V7YvXwYyr8TQ2ZCrMYPB/HEzv/lE30T0F9O8/PBu0xjGl
ddZCmIurNcHsMUewTY2GF7dsuoaTTFMAxfa6UQdofKv/XEkpzEWpvul5cp6oGjLQ4oRpBZqrWMQ5
2bpcin5NQezMZfsYWo4ID4VJT7HtVAeCaaHiCutKuqUQIAdpfFtWNrf0FZ5lzo09X6nkIbd4P2Rq
mAmopUxctDi0lwwPDnFwL3Xwh9FwOR9YUGjvXcwrI72tFABXV1BInLPwBOVPfRi7eChvUrSkNhUm
xI2J25yKgCC+I6kUv9TDCQx8V3v9kRyxbUPIuC7t6rUYC1Fy6k9tcnwoGPUdfquJUpKHuaA8dheT
rDxCTiUnslhgfuwq/02YDWEHceTWyiztdkkdVG3S/avyyEkeJznRGtNuE3NKAP830sEm3MQWEtUH
nADEmP4jm0CXwsym+gcRopafjm+HHTsryWr0gdnoZjGFFnXObVgP9z0fLMPyK+CO7IRZxm0vKDWB
dTRRsWUoTtz8GOOgUt5Mhp7XXv4I6whcN8Vt/LTIU4NXTcKSw8QDbdHvHbHpJg3m+OisGrZiUyO0
IE0UEIkRiev4TWLwzUHCWLPG878u/hj/VjSBfpxujEH4ce0f9zADEkUC5l1EdznqVe0R29DNh7C8
ZcOw6N/ROD5vVyIFRTjOOywkjF4bg/QRxG90vLyVdF/qoNS75EV1iSzwLw9vOBwdTYruWbTBryKk
LElN7hv8OjqpV+8pM/2Ypi63/1/B1E5IqXr9zYq6wZlJRbel7potStnaYf3gKZ/K3RroS+/ZGF1c
ycB3iRF/kEebAB9ltwdPV4PAvbACDw2QQ9XDIyfcR30IygCIH15hl8GKcDPF+7GPFYjvNRmTJU3Y
Q3GkC0yOQ8YbycMKu3vCDbMYAivGudu5RaQhcXSkvOLoJNaA0RLdaB9IX1sHVevGpeUUbgm9dcah
GkBejYPSwow8XFqpG/XgXAdR8EUW7e30onI6vYBq2MO/Tv36j1hBVNdmnYPzncJvOU3gPFBtk136
SG+8ezxkNc5cKUyM5KyA0QY1e5OgADTJM0krA8sH1EmWKMym3oRN3paa4npWEJ2EvWkikiIm5AuZ
me9J8GIhiqXrO+XvbXY7K3oVF94OHnq6qYacRfbGf7ov0Wd2sZSK7ty13QJTUrEzH+hVBINdpJP5
HvwQjTLtenRi+MbeuCNKqQmfkquCS60yvxe6R4EryEMSQRTnHMk9iFAWj6H1FiI1SzH3NAYvIJyc
/RrfCHXqLmx79bx/Xkoldedz1Wr2voqsS7MTKGPSE66zTTKHUPNkN7lmH7JDpGSvx6egQPlo1uoF
J3AcuVNNgXUAd0saX/11DQmImGlrDnREl0TkvhRrI78p30sT593lmLb1yOng2y+CmdtvhYx9h7Va
ZA9FJe8vlMKKuPXcT+naGGwpFiIeE/X/QXa6+4bx4RJw+NCSlj1Jrs1Y3+5vAbloMInbicB84WZP
agY4rPEzgbYWWQChG/r4Jedemk92ZOeEr4ZPwrcPzstzk0CovyC05arbvpnuLG7wZMIEL5Vqt5oP
xPah6K7j0gkpgFh3WNgd77MZCwI6+JUh4vXFje4NdQWCZacLZl2u2ISXEDAGKEIjtoUyDaa0r2T2
cEiyznMdE8XTC7QOFSK6zXtB7v2R6holcUZ+n6bMajFyHVIEWdQh+9Faa/U+EHKPB8Zors2TNnNQ
lamCJvBZfAL4j5+TQvbwlfxOvzHXBK9puDTGayM9KEKWzmM95AC0LB4V0B5luV6N7eWq5mt21Onj
1uvPvPDL47Gc78AVtzeNSTvSPh1a0yhEIThn1Ad7aSXUPe0jFeCIxe4GW1lVc5bXN6iU70961jXU
gZEJ5hVK0q1x4hTCJERPDm4Q8mL4wuOvkhFoikhoK0p4IoYzLnbnGAonSMs/b7cj0ZZZwKJSp6FF
4By3t0UqKMg0kvjKl8jtp5ajl8EjMc+JcCugZ54t7yXCk4yi15nxXFdvb5u/mhXGKBLdzKUiDp4+
lIxYiN4lZ5cbaRd5JbSz5yRVQaYDs8pheR/4TGQwaOj0UU04ZB4L5l6tLj38bTlCCGXgdQk2ZMQ3
kcsBz3A9iLPh5T6kGVbsjypMBP32HTuSo/JMOxGsFA6PPvkoX9YVqv7LSPj0OVh6VFQVy+5N8DmY
QF/iURsjPejAN1wJojzpIm//49K8nTApRTzJF3VrVaL0gnMphRcu/c33LInPq7G9HCkrVnf54/9i
RerDcfLrkasHc7ag09znLbeXF88btLMEXiuE1al+7/rbJfTUmQaTfuQEZ8Sb3ReuGQhTrDIEquGg
PTb0xDs7VFQFRZPTfHovL2iZzy5B3vWmsRhXlIxYm99HJpJEZV/tidP5mRkkvqltnmy1WdTsKDqW
Vf8FPIfMFfVKMDj4OkPmopfRpZCxpKs0i0ZFilysA8x7NiI/xtxVmyllO5O9771toVE3eIWiO3Ze
tBgRGxs895gzEcIxmjGb4dVqaZPj+cUnGFMFaigm5aqEg01NjkubjiFZcXbsr7Y44sauarW9hqgk
NDFBA7nkfK89gzv95ft71fnEGPY42QygVh1Q7tuAwhWhwQMf6Q8MFcIZrfeKzR4n2eb2H/05Qu5a
lpm+S55+oMBeCDzFymmEgrVJYnzcGrtaA7M1ykPugVOSkg6QaOhvNM25HP5H7IfWhmAgR1J1biny
VPt4BrtceE/9BcZLaZWPUqS0FfacHkcW4FGnU3TyvkmE7byPGrpOFwGYiAHQDNsuVllM0VeoYL7I
sxATXWJQ3gATTydWuMfyWqohdZ8sS494yYpfJqOR+8j870z2bWt8DEJnfE0vpYb26+xrl49M0E+n
kzEv7iUuleZ5V1wJ9PxJX3foI8alNqSpWgab/dTrgDAe9k5pkXOrzxtWFygeYxsH9/s4o5UG3hRS
okLLXWneMKk5saEJ5k+TDIUUUuGhEeTNILcOrjAJ0bAQnoPAb1dWCRj9BpOrwaKDIMgn7+pHEX4b
XjSWUcWUSrP76W6apaxMKBVjm/PUBLpauGIDrGvAZooeVJ+u2A4NdTtYggl1ifWtZD1PxJSmXzhW
HlWRo6GVLWt13rhR561zWPMk5VgobWesu3he4j5LMxIhVl9GUOXdsmpFTj+INpuelvINyLVhsOo6
z3hbz+PTdwFyH5OCcw8+jjq8slXKQrlYV3kuUwqytIRAEXGdTz/wRqw9QmTjkkEP1LX3/bafsAsd
a5pj7/yAb6enUijbiihElaHQ25zPFVYq4kypiOvwmA/rgz0UeLGLaXtC4kvz5F/5jEnbcHnccGEV
5c2e02+9ruop1ErLB1IOso2X3daoKdOqPTXPaPqJYf7PuLreBRlkZ0GzblXNNTql/ozCbtT7DsCu
npgZoe6SYFOA7900Zp8sz4RKxhLKtrSv6n05bUdzkd9qwdvHtZBFFfpkd7N7OkaFBfl1aDc7ouyX
+7T/Z8P9dHr0S4iLKOrmrXJ8Uq/KUeHJeOHOuviyl65VtDDbURk9VN4kFQ9aQDeJApd26JJuxGlu
C8sKlKQ22lbmxr/oIB61nggn/ZBidFrPybb5Au1rbwJBffpyeV4RIqMcBXbvbdyP5HgjhTUGEvA6
h5kk0SR8sUD83AJ/Hta9GPd4GDdogtJfMc5/dW4bva+aFAfIqpv2zMGKAcQPjE3JuPFukCqazlLq
WXIMwgOCbAridCjU35/dPJSUhfmXfzdDATxJyUP1XHzjCF5Uin0wA7H1fNiArnWtwIlZSDGcOnIM
TeQHVNg4VhD0nHmR0Fvd/SYEoGuyh8vtZyk64OB0Ayd4qhqhxa9BVENoSvZ4gZwviXvUgnB+vUlc
4snLHzxtkQONwiWy/1GGc8j7UffCGhDsW0yV5AbijqBa1EKMvzhxoB9qnvX4+bTOgc6DcJSp4tZs
9KXHLXyOQZJQ57CvfsfSr0YhbBb55GsMUns4cRKv/cDm0Jg+fvDcHn+aZFr+cvknKttiYaqQO948
6R1/Zn3rkS5i/t22825Vd1k13BgG37yPg3tptCWnKc0zSHjO1Sx8hvHOX0os7teOFA5v63VaSMcX
G2vWOegSrQL93hHd9DxPQ6FGex6KndprwJpE0Q3KBehi32cXXeuWYeh3MtxNuWSRFryi1P8MKRyq
eioJCx7uXIOMkYK77WTT+kNcsBdNxCiTWOs9mAxvKH9G0o9LQsWCK4aeo0T7lUjwLvyu2xb2Ka2s
t/KON6taEvc6fHL7xbCv9e/fhvVr726u8onqEESK5qUQaM1A1xkte2ECJJeqsEO9X/r1T9oE0n+3
tGVBPjnJpFx+8dMQa8xzAZ7k39FcOHPLRrfzIOMIh+iVGcMnEYW8Bg13DCuPiSZGtmYwgGNR1lwv
gaepbxPU93UOnU9gUAcE+WfSsegnIU4JboxrwWs6bWwRPJaWkrgDU6VGopLA0T5JXOffrvUJwkrP
rlVF2n9nbdSbk/ecFdr1Y9AvsMxqQIu9DpsP20rYM3/RzTiggpnlpz3V0+TM3x6R7egc/hBL4E7L
et03wu0Y5MUXOBX0Y13196mkeD1Pl/tliBcMXGsuYPQc3zJEvwqqaWKMCCtNJGASW+HEowtDL0pP
/a97P2F40XuasI94m4pDLdm2maE7wB93cstyGs8l/D/HQbQ4EGWbGiyMsKRiOK4aBlpebAB87cOb
C4isqQmi3QQi1kGTahgnRD+Pc9Slp5iLvjE3+5023aNe9wcy8BRCm1ijFbgEgW4gzPl8yzEiJ2UZ
gB1M+dgAfvh8iGlX3DCoKqKesVu02WX0/f3MmOeT4gqDtWFc7OqNkVOBXMremv7fJXOUu2BKJR1r
/yO3dM/82Ft1mVD4DYtP45XNKIWCVQO4yYEcyntf8eRLGrRE72QTF422ViJxt2TZHQpfOZ7yDRkO
zKpKY0yz+ExgaoMV1NiM4Ox7Q46qSAz0nboazW0HYVFajSwA/2j6yRs/+trO/09YJsqqVr70ag7r
/KDinuboaVv0WQ0fe/kMhNAxozFUQDkAOp+lFGRimlnbKbHff4rxDSQ7Y43Ru9RkFKN3r4I2t7qY
1TVE+qK//L4q8GRTMrOVVF7UqVfBA53/fCSWaJSNuw8w6cvKldSn63OkCQROL7LMPZDquQ4LEyii
L7DNafn6uuHwSBUeE9IzcB3xbeoIuV/TRRDeGHm6UFVqs1heJ0kbeqV0aoGTxroeqb03FI93Vo9p
4T8BB2VdrLoqaMgqTGNPD6BIxgA00yeo6D2A9uBrsRWR3qndhKbHzphYZpBvk6MXFH3X7e+noAlS
VJnrxERjuNDGKGXOjY0s0ZxBM5UrH2cSmuIONQMZDcZ9q990P/slVzOE5t+eD592yJGppVPoaFZs
ddM5GojaFEZKLRAO7TaHuPDeYhfQO90cocXmnPED+UL05Giw3UtD3zFdVi8nAGL3+ZVHHg0SVy6Z
Q7eo49NyASpjbn3CsGYOXSDLmtoVJOWjVPO4n19mgVD/d8EvycecuRfGg2PEm7Gmfc8CuwMMuc0l
2H37CdkOffVjfq32A/cmp7QTKr+qG6t2cWiUN5j0x/x83S8QDpteggRb2hx0uPxyy5obdeAEDvI+
qEMcClSx1uoOJPTOZq7WkLD9iQtBDtqY/llJmdPVUzpcrDdcz0pjZh9BEbMN9XJZWBZZAUgY1rsJ
Y4alpInKL75bqZrA+5XgU3Yxwr12eqsn/j0AGmA1sVKdJZHb2CpOTbWngq1ZOgRNI3IFnhDZ9b1n
qS5JU2aAn+Gj/8l3aZwft0C4WivF4YpFJLwztxNTM1bUq6JoJUMHhHIXf/L8ZivUJ6Q87ofoogiA
JsGQl31Uh3uVTLOkAfccLiRjHkBePXkP6eVbRM/pIqXAp+f3al5A3YOHTQ/qAAGxkQO5SL/UTGlR
gO9jRejaXLHWjGXYLop8tNMTMAmP5B5LuUGd4NDR9nHgnIOnq8PQVfsl55TrIYs/4jw2xukzBRzH
pT12QqppF2iSmldT9iWZ+w8NTI9F5S8Utr69kd2k6ki5B1We1k8NTPhvjhpJBheXgwvuYodDCItT
Ba2Cu9gQjUBc0RKiQScNQUFv7MH4dhQybLRzLVJpVgiRXwsEMmhFtcWICW8D9v2m6JiukLajmwhA
19K3nhwPnJWC6yUVNb/xuHwDGe7n2eSEai3xzCEwFT5P9Qu3WnodJ0ed2LPiLBq/GIvwzXEIb1u0
ZrbnfFJwj8msmxoqkOxBccYYN34BKjrWHKACrcbK4EUFxH47FhGo1m7/t0ssDZTl+DWXmABKxPgk
svhookm9tDzoy/LtQBna5Ion+gJmsv2BqCieetTJ4oIi7amYjru4Vd+w5BY2JhwAQ2hWDG8HZZY2
/Z7UHod7wups22Xgmk2Miv4WDDRmWV6RWWU+1s6kTWvl9LADWSQROLKvk7sa6hTv80MZgHf8KIG0
kJv/uFn5rZcmSHxvZuOvALN83ylC3xvCw4fqVqXtGC/pzkpNKm2BRQ18+Vcx33qlq8C7o3iGnHkT
2yjiA5/3K/T/7u+MV5bYVy2RB/27IlZKv/tbKmjk/v9wO649+OB2vMjqbff8E9ZieYkugyiEi95v
d2QggZNRpDzs+8+KRnkIcGfHgrBO8/zE+/hQnfO3mKpawARiqXH61xvUx2TRC62K/QT2iRRZeew6
whWw/qrgsRF9LELDCFVJ7RB9XiLvuHdVDF1Fc9GAGLQYwAPHaqXq5Or0u5bkCl7EFlwhjcD2yVab
6XNMYqnEj72aNoT1hIu1G08rwmBfklZgDMlb7AoiEPodYo4sn1ejOvvaMv/e7FGoCG2216ldrAcv
dKXu8KnYKXZtL/iXkgEEtmgZMY5NccTaQGLtt2thLCLXG0XNyKP3CDG9ixS0MTXMo/tR1goUeEhS
e2R+V3hcz1CZHEG5wS+Km/R5Zmqgu6JC8QA4R8GmCwt9FKF4iANq8iET1nlkuU8kdPakycJpe0vY
E8i9TTtxFJU6Soiwk/gFD5yTpwjbmdBwjUTAl46bAe95kZgXToxZatqW3tsu7fnnXzTrhF7HbiHS
z10O+toW0Rk8VxBfqOF/C5z1ejXZzjSI5kQ+1+JJuHnSNnz8G9tPz6F5pznTVN7vU7NzaTI22SKr
FuAdGTJfAjJgMpEdV6aCb+uFG117eqD3+dR1CIDVWSVjr0mDpRMrprGJa1NOuDOxg9WILo5kKsSG
0nkalNVs3kBFxWTKzI9RWtjbD2KfIXXPPWshVVMCnVmUKu1sj3vbSbXdC+ORc5wZ9F0R5caVwDjV
eFUKDDh2dFxA9IguoHYsRWlCNhyLwmZiNzcOZyc8I96a4iFQfX5kcGwOdRSiNPsWXE8cnmjFBGZA
gBsRLg0BZg9Y+wcmYPaUJGaC3jzeUCk/EzrInQ2HV3TDCt6eow+r09qJBiYtbe2Ahrdo4Yot5Oee
TPuEm9Mg93EpVoUOlPKGsquMOlhgp6oh+i0Wj8a5z48HAKFfNvqobuFtTi9q9wKu6QsOycSIg8Jr
AGvv+GTOdOdPdvEtKFeZEwX6fBbHepJ4uq9r4mhnowPYFRQQA/yU6tmN49pdEEoSBal0LBVWs111
v0tHBMWrMIVW2/oryBJwT5E+FcZOFHF8oynWH0juAEk246O7eUr5k0maE7IIlCGufpZBr45V0rbs
HHW5tQLBk5KKYdYSqa9mC/PWmZ81oJLs0+Rmm+sE+ynLnUqgVeTAC+O53X7X++VTeUmUeqNf+RwD
j00lfwJ7XcODN6+KcP6Z5qDy1guQqFe+PCzEu0sxwof3O2bwuaaPbfpOLTW3o63D6HfCBv5d0va6
nCoaMV4GjlTKZgA6rsOtTzYdfNSSbA55IwHbCHBLkN39xdbKzT7pD56/ShYLFKZdvCngh8Ixqcdj
IJ49vKWYLZvqkeHdb6gh/nQrEvCq8R432OsAaiqLOJC80pJP07u3t0SbcmD9m914ZXuY36VVI2Xb
hCQ1+SnIoPhswT3fd9+9/zEHXcRxpVMO7CYrUypKbP87h+Dhtu3yXfMn9IpycFrfbLJrYXjFaDK8
LBpY3wMMACnxnV/yTuKZ+cfl/MCSxVOw0Cpi94+lp1JS0as1x+nK1aiaVs6nZ0s8wk5U/2Z3+Vfv
NVYs8RSdLy5/nwvwk9jS0GsifmC4+UYon4vQkHGNKLwqVZG6s58pWln8MqsQsShHKNCf6aC/nu8H
IuyuxBFLIx4bFHke8m/hSAm8wGJaD61XEm1FvSBjgDPwlOQBZzQNOT5Old77xkROggG703PKpfWB
TIjBl1qr1uWxnb89J7uBfUe5b239IkLUpJVltMxrwtaWHkpWHlHqUkqf3KpdO3iZOrfI2Unk1Wyp
oyAWJXUSM3p1PtD+yZc8tO/2iXGXapLW8d0P+60uzI1nOEMxzKSTu8VBKcY3/cA67fIYzCjMlSdB
nCOnnF10rtItYDUK6mWJbaGJ+/Fc8BDgl2YiMUGPgoL+z/mxCbC6Us/vOHPrkn7+tUYiSLMN4JiB
MyA+Xe4gS0GM+9YkK1JY8VxLKSiP3Df3T/YmW7qwaRV40hbj/sxA/vEUJDTV+dMtzer4//beWBWK
ahTj6paaR5XUKDbhrmg+W5dizVlwYftibFiT3hW1xZCTMO+JuohZB3kVzUl/jar66nVoAkYKqjF0
nvkk9iXyA9mXmsDz7mgKN4YAUvMS436Z6sD8jHcBDukQevICoCDG4tXfpLi2P22XfvYSweNf2aOx
axBkhLh2+5eTrXNDy3y60yGwm2+S8AgRFG5Pd4COAgnsD6kP3eyw25TRL7JgtEwHxhpR4udKHH8/
TRmh6W96BJ5yl9SK01MXuaxysPxHu3ZAZ0QBfsg81zzh0zPJqlDpQyMnM6C5z0KWf2u+OjJrdl6z
YTDGBmJkxGqAriZmY1sEDX+CEvb6rwTZM0yDMe7Lx136NlSZ1sKdGiFCbj502lagiKwJ1rI1i1Im
cyNqzjrvfcYYiyb0wba0hEI1rRkWjRNSuVv0FhifC0ScGO5HnXBjUHCabBwYYfd3sOHhgYsoK4TB
GBLCjk+NAEY2OJeghgdJ2f/B6f5VSl482BEKkpN1YOUX2l7OMyKnmCsg0B/hajY75PrZs4RAOiGC
X01Y6Mmy2x9r3fB8v921ObDtrqQT3zOILkC71Q47iYpNBtI0qjJzlzmwuljWCLiasnOb6ANBvAHR
qFDv2AGQZ3v+Zg/S0FLkI/HHxGWXWkgYIEKavcIiePYtQuRwBAlbq9auf/wafMggyihISDRDXEKm
73wL5mJez0EH5fVn4gZh2ukCmDFNfAUOBxMiAV3H45sBX1s8t9QJoljsUUy7AxSAX2PfTbs/whkW
I6hcA9u1hbBr7bJoq9LyunQjFHZyBO3ZteTTry4riKYp4jWVX7M1lddqphuB6C4pR2/9vW25xtsA
xmH5K0dCHY8ViHv8FKoJFOyBe7aEXxRAaX0JjAUgmgTNe6XkKDLNZSPkEJHN6V45uGEAXX3ibp4z
rlmVTAOmIj+/8tbWr0PQuk71YE6M2ebglbpyC9VvaFykiJDbmARcYlhkiroPXskPZhhvmkUtputV
OT2YG+i0BdnN7+XHInUTP+6ZnSnPTEzba5LnXbOIv+M92L7W2co8MEayHgdaPHFQQ5D3wN1G8QGw
0ffnThBtFQae1j2xR9Qz8ZO1P7tnH1NmcxYBdmRHYKWMScCpMpr6xl2ww7oSoVHFA7glO+ZZosME
qMTkJvQ/5A7ece/eDvVu4jc4r+KvXANgV1lCUBplOLv/EFaKtzPz5PDX4VuwKu6+ngcf2DBImsdd
FhPGPDqxziNZSri4xe5kNoDXFHV2niX86M/bUpj2REjwbWdah5bAw7ZUcD1SjxTEfeP26bcNjZdX
cnYTqr8mgSB9AhhwwkEb/RSsLNJtXAr46pFvx/VJ0URT/hUpu+8kDLot3R3faPwpuIh1+u5xEqQf
iFhXTW/UoLJStdWxs/6khUrKXBFNM7msGyVxJR6lh6S8U/YWdc8IZlXYIu1jDE4rZ25EPLL1fpw9
fk1jw8ZS5XEjTNNDZdTC23RQoUNebCQhzNEz9qDXTaZmVR0MpYrZmlsIuRjD77Flem5cCjuqgEuK
Fw9CSVcGC2Vdw3IXFS0i1mLbildJB3/PGxxoRNoHHW1EGED8EQplRPSwmP8awmvBXhZirozemiSM
3+G8X+zjquPHj4QgJ/DJI4VFSh/8YyQuLSxCApWf+/tBswgsg9DuxNPQYIM4FeXajSs/fRelNvj8
7yFNU5rvlkQ8Dzl6Zxp7Tr3hKNHKBSzeG+/VIcMFrtWS6VXVF3UNqpamfa4+FapCFzZM8+WhYZZm
kIYPQR7U2BFYLQC4K4Vynf+BZpVn6EA9T/e6jrysB40ercBMm0hAFQF2q7mAeOn0phknR/7Ge3Pd
RMiRX9Pf/yteC0bcc1UR9YubejODUkR1zn7dpyOWYGxBtOmNqqD2XVHllS+PMfpoNv+nrjWH+hg6
VDhgVaaw7H1axS5WKc7jLvAz2Z/TLPiytZAw4qEtcXnWVrCwpz85XUfXFl1Q4savDvxdFF1ee7pQ
/aBC4zLZ8BVgSIkE0QNu//Fx2TiF8Kcwru82KxySsn4PakA7uOEVnSNdM8G2/0EQZjCApbdPbGyI
32km9ZvUX7lQ6hxzxlOTNjhADFJLWyPkyIVwu9VW73h9ErfjLNKEuNy+/kvaNAcDkXZYaG6EYVAK
sx2uObbDsWDNz1TC0TjH9j1E07oINKT5N17ChsL9vBhI2jP7gVFzL0CkUJdH3B5basoJoEtOWU94
KIblTxY9ZBLjaCCDwb3D7X4HJeZuWp56S+c0Fw+zqL8pj9gLiAh6qMpmHRpOpQ/QGZxs4RlPe9N5
vFcb3riRLNWG6W88+NfEnC2q9z5OcZR0TC3lFdHhB6ZsUyWoYSDJFlsnTbCjBOXR42TKq0irw5cz
jGbqqiPXASwANfcFPLgCByu5uZZdD/pHoRnzhOpixGmRf8v5r+1jS0yaOSZPdxEXB/JyH05J6uRS
99fTH5JCcG1xtBginFr23XUSeTjwEaPctevmQ9VfEweNeINPLX8vNQuLVHm60nd66L/2lwlMzREk
s7tQoSLN5K2rZvlWiXdKUFBkgpXJUv0doD64D3z7OUjb/8Zkz+97MutFkhep6S/DuaGJU6V4ZrI5
/L3YgGprmGq6evIcGgCeOszpjXnfzSc81CgERyOi/TZc+enV1acePqFJDABY39tWfyOm5po+LZpd
qt8iS7BiNEP2mobwQT7QjynvPTnBjF76PDwtZRovg2625E24AHOewrozTSG6fSJYzu9W+qJY/i7v
nRYdIF+c+8vsQ8Rh1wOPq6LtqF6o5EzK5LiGmJA6ZmxodH4Zp86Eo55s6C06NCjB+QKW/lpcyYj0
4v2Yk5O8/w84zZmGK00cx7hpoE2j/JF1ZrSzcbwOfkDWgZbTfaHXvoUTibYY2pLDhazwiOHkrQ8Y
xSv/HKGpXVbDNWpKvjc43VDNwB92DjJtkvVqpr/tNNo/7e1UXbMlZ8Meu0HT/3/PjqFHGTTE2URl
xivcqHVkWuJdDzNfUtvJORco08ANWeztuBxEiHxIR22nATLSQGVcApnSlhd9uJuMFkw6iY0NKzJS
kYyJ/tbQS3YxvDSiIeP1BWWyjDKT5C1FFv8pM9sXitsWlaoZON8QMvtTtTWSO+eFrJ8W9aFKv9OH
S/D0c2mvc4pXWxdy3zYdBzRZQya/UOt6YiZiISJcMQf3Uh/4OCbSQznaEyjlJ/QLZiVJOKTQkcw5
9Gi0MnY7VeQsUVmao2luEbR8VkOK8s6WbK8QovedmmLGJJ4rVNswVsu+mRgGlXDiA0X3bypS0eS/
/zNYG7r3Tp2VborzpTzGhSewvir5yaJuJBUqvWc1xDSxsEQDALWtzD2RGpkHKV6RG9VjTcpaOJpu
vdZ/wMxPFl5aFntgd/jZQdVqk+hWoZxjmX4Sem5cDQF35S3nuVIwF/AV7NGo1yXbCvouLoOngbUM
c3lQv+ywwMZs5FMSVmguwWyhetODs1J0JpuE+A747/T2U1ah+xxpYk6saGLSHCBd/89sJ3V9NOZa
JtUjW2U6UaTmEmy2cxmn36HrqOWRl6LWHE6GioSzC+y6ADjpwbKbbcbvdyFy4IEqxAabc/1XU5H8
qaYK7LGr3yOEWhqVHxMb4f87aAlNvOtKkov+YimOk5dLgSYUt5b434zzbUI/BvZ+Zk9gJz//UzBl
QXbNlIjnCLk5YA7A9MHIwPUr0O2VxvZ2qrGjchou/ZS27Ui95MxVFb2Q9m3+934wntFGtkWHUoSX
2l1tucM0kPCpc8Ba94X4VcBIcDqnppENB6hU8zfTmjNomeZDDirZT8BgxmnnAJ96ooRBgKvoFT7U
trUGCWCdlif0HvnG2aoCM/604WQITgKvpd2kFUvlQ2+3Z08sUF0FO7fObteqxX97GQ9t2hoFdRGa
/yJNIbVrQwUEEevpUQrsKtRPD01uxTSamSjs20q13K50EK8xJx4UFWbUALfH4gzkJcjNFxk2Eo3J
9deI14k8nyhAGScdy9VDuM2PFVFUJx5TvsinsdKcqcc1IglZLoiMCSnf6EDOHMAlKO079KNSBY8W
LWTYcUoR5qxHEBFzA1sO2a7snLNhAe9zZh0+B6i5JK1f71t5XlDLwExjojRq7hXNzuG3VgLV24wF
hjGc++BEh9fUUpsfbiw7pqm8aYBYs3wcaxmYNQsUV6u5CeUO0EXiFWSPneXcA9BhmoPiwhfqpxOZ
PbMGETmhO8NT3mwyF12Qne+3Kknx0IHprpu56+IIt7kjHhpDgg4f5CsLMd22TSYbUfNpAEIArGzr
qgvNAlkrydM5nXcoeOGRM7YOnx9VlD4v+mWbo/AuZY4znLDmS5PmGFbIfkKKIGGTZwNLEKeg+Ovf
6pGOs6ISiq3mO9vE3hUtEqJSWBK7nZAyYjHSJtvWKNEv+4HfTxZlueTkN/jggGGe6hF4PJu+md3q
pbryHRoUJS3yCQMdCcw4C62bLTsYj/NPG3yCLEr3F0NYqsggzOhX5xRmrzJn5QiHecE13qgFFSrl
YuFmukNTKJzQ315jyA6gyaE+LesLRzOXF4Ye0N//C/+FKmi2ZVNiGZuTZRQy9suETHR/qpOYAhQw
WUJlyhfwQBU1gaFhYh26xXlCPLK+UimEz/2AtIqcA5XuY3h+8BlWU6H/yirY8R/yhEYb4qkrO544
Qyfm53jrV4L4BGpcXrHHAMpPUTkm/S48RYNQH3dNfFna9iED2o9pCz+qhy4PaTlExnyCaQxIUy8U
8faQ0+uIwzIxO+M8lX8EM1vJq/oZEQVZKdahMTktQ31+0gx1IgIOtzDekSJSwHTXBmzNLz224Bw3
O2sRJuakESiYWw6Go7KIf2+Fax3jt/lrdBDx6VFItqv3vXcMVLQJ+bA1TfwZllMNe43SP1N2W0lb
AS8hRpZZEP8nLogvL1q9bLplJcM6YO59L1yv1qnobMXEE4JeJDIv8o/aJNcga+rjN84Sl12UlWJg
QIcK10XPGzvUv+fNTH+EnXOilcbQ13IbraNOYqpAREqptEx0hdMUeAat3Rax4YbfxHSOtAJcVjjc
pCa7cM/9HvPXrO77gf3ujbtSmwo1F+5irrJBaFdmLuHOuUInFXscD9Rf0gW7IWAEENTlsdxhrEzm
X36aC/6bBwXOd0UO4FkwMK9c7BaB/Dn1gWkokm10l1XVwBsH+m91hu6mVGQPHDlRcUVFO+6r9GL+
78UaTx+UzMBDQY9+5MY+Wtj5pSAPviAkkpX1PPgdxiHRhSRg6WbiHICpZ0repLVhnWlEBDdo8/jQ
uWRIXHloZXd9v0e7+7cRZQhxjG1ClI0ra7CazsxuYWWzbzF+kqjLhzNxvP9Du6Em1ITOaeVfswDM
vNIwQ5v8nWGk36TuM9ozd//3kDBf1yLCEW7HYNhA9bCeSBLUoGGKDQHmn4R9KL0XI4sWUgu6S42M
5l3at13G2lb0DF4NtedCXb32H0J1oPevPZBWHT0NUEsMJCwFFgEKia/wumfWraUwsWvmPiEQuuve
vrn1WV1iYW7jqnd/cxFa0Jstu1cYlLm3dt3G/tf67TRGdJZdx5A8r7Pe8n0DKXaDXbwlKubauR4w
mqF0Vq2kxyFE68mFVP2W6jErj2DCc8LdjHfuqibsyUo6oFNGrgNKpIbEnLMtq62merhy4nWemRyZ
DfrlbtJvuJK8pOQGq5Hp/Bf3x3aOnncw2HR6GVorBH9T/4HWHHbF3mZmGxHywaicchYUZAnJPER9
jga3rRDPzYn4imLKZ3ZQAajPuFQOmHmUlWiIPlsr/Uxix/q6ZcLsdCndfK/4rwfrfy4hj9IfVcuO
1gu9Uv74owVetPHSV70dpBSWZbJdVANmt3Cv5+TdNpPBxGp83VhdIOB8A0YAyqPQgdYf63Gg5OSu
GsP5tZ7n3uOUpr0yCkckFp1ls1ivuzofn5Zm3GyE0B70AgZ6gEm4DZfTvhe7vWDM4u0RQ6zlFt7L
EMgzaid9m5ymjCVHQ+iF/8S1ljC609kfyTVOCNfTAj7Rno1sBXoNSoo7z1Iav2Qkq2pReF34LGOS
UNayPRV5uD/hkHsvzqXtcphEMU1CD/lF+05S56l7jLVfQk4NfQHFTcR6ignLULg1vbqADJh86Paj
Tb9WGabDJRh0Tp1R5EtM2BiZdU0oQt18Ub3lBpqJ6JteRTSSQV+iMfnqYIvqGvkoM0s6jN76ujcx
KsAKq3kYaqlT/FxWOm+fpZligGMU64scufSI8CSzW1zMPP91MuKxQ3tqD4jmoHYDDg9WTvtU5Z7t
H1ubBTVvz5Z0zBP05yVVEZGW5ZlNTLT6UwAeeQpKKyWBM0Z2YsZQLTTquyO8T3MoDhJuDVhhjITl
foX+auP7qepoaizp49Uv7g0JFr5Q1t2kCicv7KbSjTh1J/ZCqkElBu06nNCIndboSUB3/JU6OCMw
CYh4LjdD3zkKaycMyqtIeZXiYjemfbnMwwAYenNmSSJfoGCesOq52vY6zITgksNLAgWo68LR/fUR
5bP17Ks5BUJU9xLsulabm8HEhKOfG6vcoYv/xi+QulpkGa7J0xhFhs1Kl4Df/7X1cjcmSwAa/0wG
rdYiw/wDqOFQw4shQpOggMgTaZpNWqCoIW6QProwxuzOd0T1k1NzZz5PGCiM2PW6qz1s2wS97kzV
nh//i4dIyfGSTRdM8z6adaqMH/uSqlD8HdewpJfWYShsAe62Av9yP+jTVw7ULyr0K2vLf2o2PNn0
zsoOl6WTo1P7IRVvUz8CD7S41EpIkKpm6M6OAD7MKj6bIyvx8a1KwGmF8a5OpcStr/yfPu5UeJgh
Oz/VqyqBXIKA+ZIkqPqXKy07gxXmUGHsJrHmljWzwO6axwq5bOh2TKItA7ngZQIrVGcBcGEnKHRh
WX+/+b0hCM1/HRH/82yP8AZi3Tb90uybHIxlHpj9M0RhHMQdPIgZBwD/vDiEI+mfTxUJv9ilnmSF
HjCyFryBH/bqSB+1333cDhjvh/7ad/v76gCG/09PbuitQ8tF7uKaGOPBNRV7SF28m2FOvkBealYR
WvxR8ulK1dwmE7S4pNKnV8u1WR+GUvyW5Cus0NtzKB8jnZsc9GAxTzvIMqqWBxWW2PyX4agsv+sO
ePQ/GMi6hBFPEje/9SpEbW84kZ2+ZXDKRUh4DzYfHWOd39bxrtzpaR3z28Cw8bHMDU0mpTSQiE+o
tkqNswCIygsYUTlDy4giMwV/4jjysHQTqFCHoKitwEoHZFKP7mVoeNxEHyh7ThjWemSSZG29Eheu
eRHF5W/qaDIGJPxGAmiKe2uNd+XOCUsmJXyhOTO1xqRx50xSGu90YLjWR0jLxoK1L+jEySC6KTrT
hnFXuJiJikAEulKXrfcL5pf17l4H2xo/tMeB+2KHoR7avcAWlWo8q2qdZCMORDqum+iHrSWHJwLY
S36Zm8NG8MGnVMguuT3HkqJhNWVWzpNeQiQAOGWIkqM4zLq3LcUqN5hh0em4z0cZTrwfhD/mlpyu
0xHgGrvg7YcMa+QhRL2V84c4/Xn55oVC/BydHyS5Qc54sz6/mKkl7cNplm0BIGbqIksJrLBEh7WO
LbxkCo131dQKA8QWiJJhH122+qLE0P4RQccMCDXYxfSmmiOZsqJ+d3nVwCgPm35FsjEg1iBut9oj
bJWx85wHzsfX8kGaFeO1d40XJ00DGRH4oKcvT1Wfsa02KJGgHMlU402zGShOy2c6pzXWm2vFu+DL
R92KZ13IAot3Sg9mkxK0mNzLyP8yrUymIYtN1R7voUNW4vZq97Xny/WhCdzgR0bdz5sV0PtgiJJC
FAAL97u2X6bT0lLfRcfkNPGnW/WU2H1+epaT2IO9jrDyeYGCRI9JDkwHuJeV9e7PmTpGpHwaEE8b
7r2vH3BjtaGghFbYQ8YcKSmOC7enOlup0ox592ZY0QfxYTtViQOIWtvU6d8UnAzrjh9+cUkt/a6+
vbRMdNUmy3C1V0DkOkXxUMqXfqiwWhP6h6Dn55W2pX3x0VfgGWy11gKB6fuXwzUhZl7bb6frTLdk
+hVOL9L1JJP4IMKz14yTdRekvD1oA6rZ32ekquaIdQGJMkrNRYePouGvQ5ZNKlD1AmYc+c8SYkrT
EswgEiJLcBAKe9/Bp15inS0X8R/DRA2J6isF1ogP9hcQ1WcxbYsTT882GbwmADMGNWkOQhkiogao
5O1y2ZPsTGyZoDuo6SqNRaqfmUfAgWx1+ZSwZFxUshgjVOn5cHHhENyeCWlFfoF43iTC/fXKpxhd
OveD1IQZtd8UEh1m0gswHN/qlcUq44ZnHivOCWYgyq5xktVsdVkysmREFSXW1Ibx9IpFBwQ930wP
GJ7DKcBVco3a7qP94M9hYYrgwYmAkqzqEQxxQn471s4W6F6Wo7UOKfqPkgeLeJrlNmCDQDgCm2oO
+Kq6Yydn2QJPunKsuiHzqWfR730xBDN44CAZPE4Q/RpE6ZABFdhez8vWXZgHR0mHokm0nkoYaf43
EPnSdQ9cZV/Qd4bsdvOM7Z3W5wV3R9CJkJAGBFW3NklN15dqf3EZqCoQqeHcQF4Pbf0X4aV4R6mw
pHo2yzUUPDF9+iOFDzqC2lnmq7rtUfRQITb7hh1Egai6MSqEBOL1IdEy2+Xzx6vkO6gedspx7WZi
sU9szLNDbxUDiPP4WX7gNapSjT3tFxGd/C5t3FYtCD5eiu7f/kwGZ2dniuEgd/4wsdOBEViSIiaJ
QNZvsaOHrCyYw10tmaljY2zkUz5OCxUFokD4ctXOasA2z6CmzHeG//UTaRm+AjgkTeObR61rSxIJ
IfOMsQcSiloIQIgs0SlFlO4zdEib3asCX/4NS+ceT0nvkFB44PELWja7cU6p2lGcVA04cfT1iGWz
oq6/tBM2mSLELinla+2h0PFqk/Ozgvgvzqczm7FHrOKYvdWQSayBdb4D/7uWtlU+vzv1H8cSSVnl
l9IUzdl7cnXffUc2gX9TlJqvz3x0c5OOZ4uk04YZ7soRamMS0MvBo6vIQBTvpPi94v3hsHIHGxCg
Q2WhWNllZWQAyy24gKXZRLYrAOVpiUn0p2gZhOF/PQr7hlG3RqLM9jO/z2asGrfwcYbOV5orPWqU
Fp8dk3zvl5qB5RPeuLrYVQz7zE77Xs7Ef8smWeAJzUiMB74QxwMUI+4DFXN10mLOJID8mYouNs1y
9GdKwnh2iscGd2xOC+VkAZ6gqt0revkoQcLq5FuU7z6/H/jTkEPXLt5irTepXR4Kc7/lNrTtSxYR
FSYW1/HIUqDSMsu3Lm8KCw/HGXlEjRfcWPUWqGfyPZ20I0jd7dy5RGE24CIiEOEnkB4ZfbBQ+aBc
+HsTvSVu6WPkvrwlWFL+8UFq+HT//1DAuIcu4eEpo+aPyvzPHf+GfnVFCFCNEFNwoVMgMlt3Hf4E
zbD/Vz64uVhgaiZ60h2Tm6L2qjvamQCjW89aFPLN3vibZ1c9XNbWWVgDTT+AzUbxIXZJTirVT+en
lz1eRzvWMGxvS+Xs3RStr1Oi4ZgwJeko/TuBlNB5kQUB5GhMVl2+j6q+G+LWevBeftGo3NV2YeRP
l+7UisNiIkmf+sZq7VNvdcEFcijZTIM08u6Igmm18SPV2jdCbQMPDVmipi4opI8KcVhCNHJNFlpE
r7LHZ6EEQuC1m1y/du7c7DTEkjGR+2Y7/zOI5Oiotm/Cfk4eqDuuUT5FPEFjw1d8A3+E2qKsqr0k
2L6Yxbb4Uq53ap3DYPeg4JDIkGv+hbhMppL4peSXjhIAqg+HqMg804YE0OAM/iyhDaYac0Oukrm8
nP2ir41wK1M9REYYXfxO/KrtX0Mh0t/gSrtJ7yzxY9R5yhQ7UdrMRNXASnqQMwtZFS8ggn1oIEle
LmeO5x4HCmJ6Oe2chXiScbErg4ATXOmdVHWlI52bGOGhxBY97jIwRLh11QIZSdEdkKxL8lzaXRV2
dlXg/wYFBf/FsT0gQY3y9fPu7YDUfX7yGP++NB9TceJ7KiEfsQk2/KLQ/+OFtt+NRgo89VnyG4f8
IbWXoWIuMYBI+bYfMuzW3jwWS2LCHkESZkwCMl0bURAFt6pyfLPHWYWQT9y0EM5r0vG2Kbtaenne
UxHBVLrWP67xQAgW3NQC55RwQP3owsIrcCBRe0M3LOPX51zPNOGNOj4eaczbFAe7A51vgoV1AQQw
j1ymNwr+fEJ18heVPuO71UMHLa1Mh0FPJY3nff0RxlV/DJlZfVtTU/oXrdOKtbRrMKKOCK9kKh/y
Qw+xul4ZDR0/hxXV+QQLrR8EIiy2j5/wM7kZwBqDz7VOo5wToigsO/esJOOxnll32tfpdald1+2d
Bt7eQztk7g/VkMYgQLSk7VcX0of0JmUHh6YBvkNzdRu+X6k94Kc7uJm5rrhKEWDzYInGF/+hzhR5
8AFNIHTYORjfowdbLhq+bvnr4o2S0x93YuJhJH8GuR1PtkXYOnoI5mrr9w8uHOAGsH6znWF0JF9V
ZSRHmKRnd0PZDn9pxlwiJzow10iAWtgb2uMBQCfAU8dy/T5s+6sPpSujcnqOkkfCKTvRM9a+T3dR
i+o5fP7+YTcsW+q3ZzfiN3WBbVjbWdVGtZooKnWDxz7JIC5XPesTaV+btJcE024T1o06I98UGo7K
WWb+5+TUUKyJbAP6DDmvUSqmpBSNNTZHQciC1Q2FGKx21QUiq19DVvrMvD+KdA9NKs6Uq6KW8mHk
aqeikPxI5rmMzG7aBteXnFHCvaAFpKNquu6UZ2cacZBDyMRZEqZPDAPx4Y+p/0MyHTihpAIs2ixk
en75H0+uI36kUIscmoL0qejOgpLuFjtllh4EOyEX7teeGuToTQ9ZgMnBDXLyhA7wT82nypBV0H1y
OAJmdm6MuuIFQ2evN6/TPoMKvJBVJMJR7TXXCjrwyvWQBR82o/qZxXbwfvXqn+EJCuzft1isk6r/
vZL/Np2gezJ+5mUi0ljgCZj2RTPsb2nPUkMz1x84tfLaiq5TlL9qUKiZc8+ySPxkEne+VWduroWE
CpitezAn3SdMX1UQx9weC3wxR6soaTwNlnIVDXMwlGjas1yqVba9jL1iupqKv1lG7H3rX3adr5ya
8E0IUrZWdyF8cpc2agnSHtWUQd0XGxrCrsyKfTqna0EqOSEKJRGt72qxdJsFc3pJUl6YRWcjkKBa
JOqqj5bq/7PupjfqO1MqjrYYS5mrnC8uWNGJN4+uNPasJorMnhKO+2iunPh/S8eh+ypNSoF06Rp1
MkHJ6wT46lzWJVJPARqUntAH97jj2XRmhNGFa8Q70lg1ZRJzzX1ixF/10WSetH862aNiMUeKUpJF
o1U84j3sbQnHGIaSy27SloMfT128YvDlfdWXFtr21MKV1hF+jGNlTVgbt6pbiK677/Kad9xg4To9
wSgv6HhNJHDrIDVgYv4iH7uhu4IfxyxdzGOA1NI8dSLhWZqN98Us3Z3u9TwI5/X10q6jWdGFoX62
4gghJWiN2Yx/R1eY3N74zJeh3xxR3xTWHJSX+hVkXNQizLAZp1iXXjnI2MMWaL+8z9H3pt+aLHum
Yy3NiTmPiCneqqmNObo+moo/LdKqU4JV/F4HtpzlK7p/1JuZeoV7OuW8f9xdgMVs2tSLGhH7jTQA
XDu5XFBsK9o7nQbhM/Pt9GTqDStf5ywCVwblQ0r4tPzU1d00cruE8Ci1c56yAfSxxFgdeLeLAB8e
zsoW3rQ5DxBNosyMu+GoBuFpeThwLLInpw0SQcTbDNT4MW2yA0Dx4JX+/4h+PZ4O5P1LkcnqlKWY
epLboPlrRFWbm+zNPlLnadI44i/fDE31ER3mNwABRlKjmlqoSzmOAQsMkcE27UbxYI1RlKqvmn1d
ePnCzvOSKzNlneQ5EBfvMk7JOlMy8puhw6dx455QuiRcU2CvDYCN5ALd71tzl3u3JPM5jQAsrp41
iZgMC51P9FRosK6VW7kSDh+NS8yTdrMWa93CU3j+VahhAUCe+YL5B+yINTC1BoYMu57NbjlfkO1r
4bcSsqG0dIEK2NAQHvtutS+92ofulTVe2s4namN5K0Zg6Em//nICh+lSuS59q4BnGtivwb9Dv7xe
r9gVcHtwIpY0cttsUanYEhA++aGInmMXc/ydZ1l/jNdBveX8eik6XbSk9ubcj33bkyTyVht3e4yb
lfnt8btecMILW0lVImTiZOxycLO0JaAj8D6D4HqJg6nl5VZAm35k7fUUs8g3XyZOnZ/VitYspA/9
fOgUUdpZV+N6zdDkKN1wFeR+MP6L92sAsut1nMWf22/sOtYmoUcp0veR7vgIfvB7v/3n2I96xfg8
Tly70zkiN0oD8CmoJTE5eRP2PXJAggmmvh5TgyLWspNFqaazNOq6X1KbSqoPdKOfaq+WCJXkwnfn
Eat71i6hzlZr57lq5VjVQnEMX0FhUgLC0ccj1kL1hcr+wYGVx5Ip8MNPYz9wtS/M702wFI5flDAg
kBOOOF40hsmbqLL6+sNYP3Lgr4vER6+whehMuOgEgXx7vU2s6aTIsnIjyi208k/SHDCL2i9G4h2L
KsaWic8pnqJUKAHGTtldCCnI3if1AJ8Cvz7bI7t6QsGPbtqnb/mq8JcRkgQ8VDQtd4/ivhFtvk/E
m7WrwKxAf1bXJ6SHNmIZJOBG7MwvVvxtaN/1jLF+9BV8mujpaci+cyRLBKaZ6htMnzuaWXsV4oLf
BsCOQRSqfrSWRALqUyZHIhxvbK9i6gTDeuInNV+g/IX0OclbI34Tx5/tRI2O6+fQbiZuqftTqOVZ
tZxcfFHSeKatS1p2Q35TL8TLRiV6FuPf6EuEYAsdOGvOEZv3l5/i7z2g/qaoZyYLgvG6si2FDeJd
dZjlmzKv+w+3cRYAn92lvZVkHmOx6bV6uVC/93exUTXAduZ2Od6Ga2CXJtvSg5jTpfmW9ajbE1Ru
xzPo20q9V3ReHnALcjpn5P75iKU2CqjwdKFl4ChxbcJ3kUPIBXMh8s7LRDaS+4HkK+74/6mUin5o
Lfc3XTZQKFzNCuCrF32eZe3VugJgjY1u+XdFL2OZRGGiUf8OWmcImir00qtrxzrQeYaDbjqMiQFm
YoE9dW54Q7GBK+wobQqDe1xgUVrUlTHg73Kip9j8IGWrVkg3Ok1OxPpu5bRrrebNnx3DIp8j3sAF
1enoFw3eftPwpRTKNt6mNTT2KXuvUoXEwh7ACCWSHY08jSvvafG0bYOq3FIcqZ/kfAeqgyiD71Kg
kLANrw+25Xo4k/vKu3RD9/8bDwwJslhGXXeFrHxvRDgGV8BneFqfROTKurUlNyz4ZbndctVAZAm5
u6ftRLqbybNfALJFazIG0/JtYEWDRiUycJtyejU6awjl6MDP68CXkgsuuggjQC31Yw+cKmX+xcRg
5BqHcS7WktpXETWAt9S4ZOhGLjoeBstANsBlpX0k/g3Z6DxRa8SPFMDeiV5P/FxVv9PGlxAr5mYQ
ETKWx2/QSvrAEyiZKVb3IgpFVQKMgy/qQx4dYJb23Qk4dyq8bYtnxFrFLV4aFHZz4thlzf+UeMs4
Z2twS0NYCIj2lLMmhbTPOYG/rIHFr3Ig2b2ErTpUMMGnDGeD/4NuTrLNOtXctE4b4PoQmuzrKkZj
S+obXUnqXIccM3gCz4B7odJToFqxS1BpvE7T8nfs1H4fyhxgtFAqWvQVk/zSn3KZNU4cDxzZMYZS
YemuULDwHfjTxXQxYY/g93afOinUSkuPuSQtiFP8W5NlGrGe+xojOhl7VlpamjFx2KnumQG8u6IU
P9pkbbjPl1sa46HiQS43NpEC6/eUErtYYYOWC9yKRu09W71arJRnHgpM+hZ0GGPadOa7YC2TwuMr
JS3hG1n8v0fj8nZwp+864e8rHezlM8Lu+F5eh3jg+9iL6kP5mumUpI95D6gsVwC2564QSgvJCnJz
zPpa8wqwGjGYEf8brM80vTiMCwKPlNgIUQHNvKyrI8iwgwpOgqLJQks6/oxlo/Cx7Ul5rGTrY8dU
D0C573D90J/iTPm4ZgXiDEO6RyO/wCAM++AqubgBEySK0FAlbxpuerLJOVMb7354Hg6oA100Bf/d
BHto8TXFPIXwdLMdMDKmj83lZqVFMiLMOSQp84Qpy1aklY35oLoQa4QT/XT7Unl5oRiFk+HtQCGU
kSokhgrXA89jgFFDrWac/IOulvVxN2e7qWnUkRzvZ1eqrCiVd1HW5EcK1H5oB4+aOVjSllRQxDxL
ueuE+vpUgJoG0Eu6rH0giLEXleoU+R8FIuKuIfbxys01DPhAYYW7HNp84o73tgoy0RK7c6JUoeAQ
woZcjL89E1+ngdKpVsaV3sum242lZk0EJWBskoTa5P3Oqf5+TlJLmSgrsrP6hz6DPXCgGpaLx4Ur
97ZnUUFAdqlLLELuMoA5fpreg6+Uhsh1sCe+IF074kgxdVdpKnyKhX6KJ8lYLyUOnPV+45yd2JBd
xWrWHU8826WydK6tPpfSzW05M+M+njOUNzvjgxihsN6cfSpSwtQFqqVgOjBDVqD2i5mc4iTpfLJ9
8NBYz2IJw+efzsKV3QBSJ/UcFpG/FsvX2IqSCB23pNU3l4BUDb7mquaSj5Om/+oIN/4BLiMip/Ky
6qe/6A+m7mFpAHPawITGHhzeLjYgin6WdwRMNc03lTOcHrzkIzPOASCqp342NqGylCtHrUTYkn0B
k5LeuP1lDxZcbTVwqDhFaAwz6ZjKisSVbMIATKGBMnxPzdTx0SHofHencbgujGhB1HsiBNOmtxTE
CWXOrcHYYCJhuBbkl1Yczx+laRYQG3y84R3CVtCCkTsTs46RRHbStvN1Cyr2ztwQ95mzdMKAggH3
xThtUQMl+a3iIwqpxVYRPtYZrdVnt2BJrcNhasDLTmYBNV4ez6rASm9lT6ua2wj3Y1rYCL5YfqWD
rQl7L69wA8ttgR+UtGHx3yBycwwgGu7XYcwBv4MHUh0WM4RgCbDidlfrArwU4QfRipwtr+IuEjBR
M/njep1pimBx32oPPc2Z01TgRFczUYgU9hhwagjZRAcMYo0Po/yds5JqIvHMJb3e+2X9U2xcZrfP
kGl1hLDquTj/1xrAZ4XR3DnYZ8PxkcpTRSiC1LHe2fgGUpvM2lzkt5lzGUfplSNGuaH6S2XH2peR
9a55wK2zQfuaZTGh+YNB9Lmvy9h91+xvOgsYVq8HM7zOutd1j2Gmsh+OuJR75nxCWKNFCtEKvSS9
evwqieQgjc3+uvKgMcTjgrmtdbXZ+g9TdV37HJmQN6Tx/Xm3UWa6TSal9cK8dceVc3VJHae5K/1z
p6QX46K3B/6WwbuB261X7HqhH/KFh06Lx6jgVIY7Fe5H601MaUhXCoFb/PuUu9aFx6q2utiOlQth
oWHGo8Mu71JVwo7V5lO2Mba47DPZbjKBCyLMT+ZF/Q089BLkm1DCTGQsZ9gsNWZD2SDvoqpzFLdH
S0IooJNKYfWsH6++op0oihFIvg5vQngTaS7XAoIYlHIyKLBO0nzE8amPo772NygPWJ+/vJaFFSDQ
kOWomwAafkxegCnteF5RFuFXEyD1yyVu681ogyyrLafXTuJ5FbUZYoa1rL8Gp4Bq0RlqbyCcYsFf
jKF/7343rCTmyM+bu9nI12uBBl3SOrWLtauhkS8jCvE194t9woXMaaBRfXJUEiz/z/SBMC6gyMic
EDKO6mpKmeB48l6C6y4EnbAYWnuaJ8hlXEFznlXnyrqSYLzTX9vx4C8PmqE9D1zfGa0lNijb8FG6
IutmjkLGrhK70LV8N85o84gXhMnoUUziUv4uT9xkDj6pczYpcBJo14ED9HgSlkyKIONJiZHcb9Hx
E8rEC1n99zrCtgei1eKPTHbd1R1BkpCnM7BxQ6PczPzL2Oy+Nk1cjSTI1XY6iNoFxoCi34uAUMBp
8mbwpdgsptdt/eXlYKw076+Ep0yPVUj2fVX4QUlX1ZIplQ5sb+QW1jq7UQrOAInOh6vyNZbUWMX1
Oro61hUwSegrXvzjd+NIeaIXU8GBR596gGKmJvn1me9Ccx4B3vVUCO329QQYPYDRW7GFi9Odqi3T
owBPHUK/KLiKKz3kIbb+ap+zYOZXoEV7oeLseMSuD72t8Pewu/YSov9LGCZwxa90B+3VIsIItrKh
6MMg4I6pC+fUY1Eo66fvpYZXtQ/o3yd8EU8InnCnWKU+S9E/Ica7dehhyg0Hq3a5cA0jKqgkk60Q
vmIOxzXZVAlXhRXYGWORJfy2QKm5In0ieV80XoEslqOpW2j018Z67BlXgxi1LMG+GlEgtS0TscF5
CFdnggnsJFeGEXLED2gBvdaIn7dpAtO7RuxHm3pn6SGm50xCRt/3mEk/hm2zdeG47jMl+965GZER
L1vSMVc96S/d7VZ/n4G8/fM6TUpA1mHyVFxVPEtDXbicwZCPL2vPTaXq+aapYYr3O5dcDzE2brti
MJvnwPAYW5GZQCOaaW+egecB3y2O/Gc1RGE8Q2w2Vz6qhmhcs1/AeQMv756SeV0pu8oVTwEb6Icn
EfOhbhE6LLY4KM80Wm8WFuLNRCBRTxcQveedGPviIkhl55OGg+sAVEABzkH/T2MAk/5QlMHs4vqp
fu23+h+4yhueNG5fbcY1vJPCTb00AU6kYQZscDe3qcKcyq20QpqyOzCCLAkuf5ZVElLiSTQz+25c
YX/WJIhVa4AZmAJQk83B96vflscYy8KBb7MRu4kGOVhcgtejkRbHJiXXv3IKOZXlZ0Ktq0JlQagO
Ns7jvtNbReiCVjnOLEpNe77d6AMTtkzsMDd8PhezwEMkXuEe9XC9nwi5QeCNcIR14YNMkulQ7aBr
2FmvA1t5xWJl3Vx1GjZbK2Qc30r6uP/gFvMnt0tyUkDOSZdyDiCadc3AvNEzsh7ZsIyzOGUP35ip
0G8lJmvvXzqm2K7bUG2TzxeWXrwU5l0hfZAyNBJvT79mZd+bq8JWWaZh5v2wLYlJBALaF3MGw0mc
U6Z8Lfuk62d3ygzRl5A/kmLWhh+CuVc4OkUUOlB1Jma0XUAqhwmQzbdOPmkPEEOuZyhHJZn52ux8
oJqZnIs/RbqSUApnnFRX1+xMLmVyKDXMqJeZ8MPJo74i/ho1Bz+GLmle/bIBGR5sLJpFqKNGAsLK
ZZuGLwcuaBf2k5er8YJQD3ij8vYVfMbP1R5CxfDjdaTN29gB4cJqc+rPsBaszu59xx+/lVNysgQ+
GbzVYhUHqZCBIRQvF/FrYVey893989kTFfMblyXHH/AvHflrPr5G7NAUmg/0xHtwHS09w6gSA21+
wdHboHucrKYehBgcSEaxy3yPmI3ojUAU37272jp5rUrVNo2gHmRiOBtR/KpHr3sGHnRRSVqXwDsS
Y8aA6m3aNlH1YZMEnaVaX/uQpjAvesrLhRtrmC8pide8Xb6Usgdi1jYb+cyys8S3uGATHrXOwzaO
31T7gWzQS89wNARFSpSx2I8kIBSjPqWYrHZcFx/s/qhTzV27hmrPD4oj8k57nkOS0QMr/45fhh68
UL5R6ghWCx9IBShZuL02ZIF1JeHz+j7PFKAsvpfZUDETWk4Pe/UkBIG3f6iHie1VfoLH3onWEQAC
bcbENhd5v8Y+5bksr5uaE6OD/UlTGIfRFY8BXFXu0rW+uGwot3/rb8UL4wNGnHaJ9nvkOpafhHgu
ak7+A2/y6a7jOTRLDarpTMcVfVX6SqP6beLgGLiYeeoqy5mqEACUedFIQ3+/hxGJzdbAqX8R04JA
a8MlYRPkiwYZVRtCzsfgNryTemPLezFJac4qTYrkQGnjLVrL9k3lsyzHre+X8XBMoqXXxB3YfxSC
Wh3l2NA8brF9YGDa8AEn/Wm/678y/oxdyuw/w5KyzKhQx8FmqUr1HGSq+pfeBjxkCzHPFyo/Th9T
OC/dhY+AXykiSML08/+hCODxLH/NF+ey+mB1QZht3cEvnGhsH4y3Dtnv35dIXuiKCe3O4KzhCxRE
I0nDC1LGcCvN1IWsKLUB+WILYPMv4DHdyQeiK+lfgZIM7xqyh5qNN8Bjk0B0WhqFNwXF2we8OJrq
ewSLXVblJkLu4cs4gFcqyyoY8gx6T7adPK626VWgD5NjcheiNHsafzITmVoJawjFVC1GsKVjhQQP
R7M4tpqYrQQyeuDXMYReQTFvdKKP8J7qtXkgirkFnil+wHHTGAHV8aEZQXOmshMld58iauuH8Kpo
nxbXr9W3t1d28E9yG7Vva7Kjj9GCzhGPqcABn+l337bYLUgsR4zHQhRwd6+OFe/rpVwslmKX4alM
T9FyjpZk6TvHiGfqrXjQ6Z/kjG7jdnJI1FwOIybDuPt+IImkdfb7mcKxWj/t2xgc0eoXfPgCfMT1
hsNlERIBye/MUGiGoaOqC3jZILMv3oUyvVFaRTnLuTvEDTrMnjBu+1HmoA7y1JypbRZIuQ90vkQL
JBG0rlha8PYcg3lgMT+EVfnW+H7wAtOwAiOQYGIxsNPCnij0UBMecCcOiL1UIX9SfauYNHQ45fHo
UOeuASBiISkST9MU3i50qoN0HEcdnaFG9PM75RkyvUWdU2FvMkvik89HB2Ct1lX/G6bMGrNUZ6EO
WVSc48QSFbL1PVh31YUY9957dd68jlgokju1SsEE4djxmH2/Qh/AjC4JOW5xhZCaYYyxlx0rXw0N
qekeNQfc8cbwGmXmVVQxY3dDG7ms0PPits46yyVYRPfgz+DPdaNw2RLtv5jhPtzsSI0QoCxPnioI
6TJatzHuJata4Y2BUUIZlVfBcMXPxkLVs8W95vAjSk4nyYjpGIrTxAvPIY86zWIagc5RCp5MZw+u
aTjgYPF+TwfIKKP6e1bDdDG7BWvUW2PuvFg2uPe4+9+Ver4XA8FOJ5itbxi516NZPEBJxjKnYBIS
2sec0e1D8V/xNjlNc7ESbK3OvNvlk0BjLLFhPV/a43bzDpcewYVlHMmAd+A/5G7w6cKQ9/EuiUU/
XPtHlV/xuZt+e3OSRIQO2kuU5V9ilxKK2/RdWv+YscFcLN5OpeTfetmvQQLVlQXRPpgboM1XbKVV
ygMm+U2g73Yb2zG7KEY4k0PM6/2YyRLjBaIe5UfbSOtH1tlYKyJVfcnEpm+d1FEJUogcyNPSoB6w
4q8RX+/QTo1xGdJsGaWWZZKpP/VkMMwW6M4XVvdulaiRkWP3TLT1WxbzwKrni2CM5C+CCteVq1P5
Q/HQ3CV1/fUojxWgShBsVOtG/PBt1ZouqTKJQubAjKbSA8wGwykDp/lgUFinXUUCheTSv/f6L0d9
5EZmV0bEL4kPRfQBjrnOZOpVqyLSrFWyF8hOezV0mNpMx3OKgpc0ildNLqr780ItDx+l/tkyRJsk
qRtau8+BWyE7Faf3Dt8a3uXw8PmW2o6Dez/UZfvEYJ86zZPn8Ts0N+D2G1zCOD0AF452sr0n4JPQ
F/LfdJHOT97x42YM2/qNftAHgkR49ggM4CeX0byhpqFrcUGoWBALvRmVw2Z/YnSX7UxLpFApG2aO
2bLoFOWsGpSW+2APxPtFLLNw8ERl2IZXmjwuFFs1eJ+gyAoCLaLqYmfgFlzgdcRHljFUS9OtCH8b
BEtXFljmBZCoe3zRKTiUW2AGSj0K9sISLcgPtTuTM9R3E8HKMMerjQnXJZBtAUaEUJtzcRXMg9an
fyd8l5VfEhRzVtrBPQn2mRis095ldIBXF2jRtXSwoeu5cQF+4/IbFcKIBG7r9QIMz+/eyqjgvwB3
CfTqOoLxSeE2BRYKN0CnYomJMi7A2wYnpYGkoQ8guedPOewsXzX5xyxLUKtEuiaaxWAyoKlwCnQN
6ld2VroEdJVv59wFqChfk7q5sY+OU3T7jQi9YxQ/sf1+G5Ln9+F6eYMQed/Q57DTnAEaGL57ohSB
AazSlcgahEGsRcEg0nur8L7PDDh5qksTGwE+6j4XnE4Xj0FG6UMvSx+n4EEiMzJGCoC0273xcSX1
HQ/0M05MEUuwzuM7HMfvmIso2xw5yKrMpJPtOvdUFv+0DSfaMAd3MxKUIuRy+iFrLQkIwKrbZcEN
GFFf/6JwHgmV/Pmp7vZpC9kG/633atHkYiFQ+5s5bwu7QCWdkOdniVdLDoaw5R64NUYDw9fHxHt2
oAeP8sg1/kl15I+zHiDHsp/OeFRoUlpx/r/chppEzZxG1WWZUUaX4Xm+SEFop1p8saHog6PZRw6M
K7LDn8C5Vp0AGOsVbVttesxDhEfqJR/dNYFZAirLDaY1FmktwAm2cGenuLkWD4hv+9pMAF37Xdyg
/Q9nUDpMKQ6rTAjh1eB/rO3iP3dS294tU41Q6SecaqA6qsUR2GrARdW8QRseiisMeoNir+8tNAnQ
up/nlDiCjrrVRxwnJcTB0p1dfTpfaXCIToqR3KUTL16UgONHQd9RHHCqeB6+uIQ9wmm4IFRlFexf
be9cPMo+4DaRdA47v+TjsUTsODsXgrW8YKpUqRMTV1Em5tcUySnGeiDshvHbyv4SOF0F//UR6Ttr
BYijBwQ8ci+t0c1/fqIaigwAPeLP2c+Kmhee2slRyyLdAOZsgER+o1OmDoCEOgXMq1tL2YPng0Gk
hecap3TKRiyKXA5Y1NJW3y+uB1lvD4+Ufpnp7KNZAuSy969aFM4IuJmqg41e3PxE77snL11cDue/
t54P5OyBQGu0q4lYELyxln+zIRkdo0e02iim5JkO/UgcttjfVYQClyxee5+UlWKaQUYZD49b6Reo
/cz98YPW/0LreTDFmoYHIVA8LYyVldUzCZ1VLA1Ofztl6cimWg98gvCbz0neoL9nfZBjgXxqbVBG
0EAod1nCCzLOguCmavfRLbMHhhowOUPZ45tJOBVWbnzC8dooFfzswMLnP9mYB7vbYynIrAMh7bUr
/Jsi6TkHykJUdXBH+XD3V7b+60YEQSWOg67tRflUJeq3A0Z9X7H6u8/2CQ67Z2X+WlJEbL8yywRM
MEQrRNGBX/TNX2aAhf60PkAM6xx8oYhPDT9PorrmWBoM2VoCot4vqJVCfkadcmMwxKb0SLxknLAl
/sxxyik1WHu+CiSVHUoLTIHcpJiXYoKXGg/60k+XJOZtL9OLCmOmGJUfKzKflN4YVk9KGXs3pVPi
KL0cdqPujkTYXvrTOxEDVpSvO0wwWstzbha0aoF24UzxRKGQdx6f4JXYPtdXzY8X4qcNbzELK9nt
cG1eVzF3XvVPGetmcUFnLF672OCUNPuVcNY5Iv5fRP7oR733vQmvbSKhp4IkdtCOdLBkYvSe3dVC
M3AZdCiJhMWwRWmADr+rltMnj+naK1/7D4sQQGnkTB4OV4qvPrOGLGqI4hX/CZFIpMWod1XAx3FK
WH+6SP8MQ8/OVA9xQ762lrby4rhDGKVkj3La6elrg9M6u+eBQRvAdbDRLhWz/AGhgrI+uEkQNWFZ
L1y3fEypf5EbB2X56S48GULhMWfdUC/W7sWd7dm0cXcvSGM4eZi21oaM7shreWiqNzoXiBP67BnN
aNrPVHYktSFvfGWG+S4zqiLziJPMdLhdkxXNiy1iiFmadqSW44DkrVKsNIHKPUwt09vQMIO/Mtcl
soUCWGYUXwArb4+Eh+TdjjGGTInw7TPUgPF1SfCepEJLUrFyAFN/0nWYjytQBgWlr6bEw/rDIo/L
o3KlCWlb2J+fN171YsYKNEiboPU162jKvolPrfDBop3dpNZ6YNVeo3AgQ6/GIdMghdKrFM1rsV9O
Mj7cr8X4FcQQvc10yrXGKPaIlgvP+TTZEgyhBUxB32Rfdp62nObUaNREz8cFST1xV8gv3pP4tB2F
zM7YReGzQ4PqkKzB9GcqCHd4PI4JV/0mWDWNRKNrC51EMiAB1ojTgYBOAh9BzeRzW4K7auX1oJUk
tyDV00KMidO9Qctm1jUTByo7ysx3MHQw2K9jzMYc007FNVuhOGhRz/OKlaJ5TWCcffKZVz3IcCpd
3PJz8uEq6Cyaan/j8GiuR2SZapWJIRrDU8EN4BetPxuj3ljzSPk+edy2fgjID6zq5joo5jNphe/U
B/Z17XCMbamw/JeFFWhFu28msEkMmN1UnY2dtqhQutx/RKy1Ht1bNeVSmwkx/82b8QHyZjRgrFS+
i89S1rTjJD48IAS46fh5/M8Mr0t87D9lvgCoEfsxQg2wF6lSIxiR9axWUpRTdKfKr5O1cgDeF+6Y
x99H4ax8Q6wQ0JIs3AsPoALsF1Ff/XjfbVv/wE7z9EsHL/UR/GLrrXJUzXPbmaodQK4HuI1vw6hw
glLwrbWp4soYjDp3qLiKPqmZJIUxuKLeG9xnMaR4QSukC0+Lu3c1lbKczQyA6PZIs4Q9BXWcO35S
cGXLvt/SrX0h0Qn4A7pEDKE34YrcnHeHDMEYIfRQO1p8WCgnEcZuIL8djIuCqCBR7jA4fwg9tnQC
ZDFVaoBHMPax2YcwJKxFGWNey1m1avuae0zkawiK0CU3xDWCqYgdIPWsXZtI6M9FBqNwns1/SMr7
5EVqZQhfn/LQs4KMvksPiOD3rqH3x+bypEUlOBgSvW4THUPVvO/o9PCa2lCI+CiTFa3SH7bzzSme
P8gutR2bpckXHNrd4UbYQs1VbBIvH+g2s0VOw9k0igdG/RZev5lye+8xl27VKtervp9OvRqVLbYr
wVAfnZt3+tKzmHHJ2md64Ul5hBj44K/oQJmYA82E+m0VR2D8+JKdE7Qkbt0vnoI6aOjrySKbWUSG
n+4BHfGQCZ4DfPwckAWXfF/ZfKY7VlKjvC0CA/+FQSRNEdjrLjw9UctBKZJF6MZMtQephZdT326b
+SN3WJ1AiHNQkUa98Ry4f636qMkQodEJhuTF/mePxpom/3oSUoSjgaxVKiLWDz1fZg7Dob8LDmm4
b3qnCvLJP+Ojg9C8VEeCzWVxcLw6zjFrzN5YETMVs+MzuCde7y2Y3ZiGAM4/lHS/Z7okmFgsmM7Y
VJ9TVWQim3F7bwZLbyT89To7ZPaDGr6EbyJ+6V5imKjtC30/VFd5GQikeVHk+d1RSLiFXfujXoqm
reQ9NleaIwswP2+yAvINZ4bHKYCrWci61TO4OuipBFc8B8OEca7O/nafIYxxL0pAbnDiIS/KZG+g
XVsVjcm8zvg1rKaJAFDntezDAAZrzVBmkUAW4JRVLGAzFowt4Iop7RnU13z/nJZ0A4MA1qIQ7B4f
cHj/mOVWglDbgqQTP6GUJtvDbqzX7Am9SwSiBTagymltgQNCkeYaRsvlpWdWiy6+2f2U+64+Wd52
P0wzlM4mt/Ey65g1aI5bpT39sd0csyhPSzfwvnIajrs0re6mz3mucYRKy49lgX/mr1jNVGlMIhGM
P1I1hnf/zhY1mileShaUq7kKgc2luhBXEU6choPd7QEiHzGBT2ANJyqMNJ+wvsDsetNR4vW27LOp
JLaOOoHRQIrbML2u7p8HIUeskQ0Huh6bpY7sM93grNDR6Tip4CDFqpRaqGbuAqQP/ypQSlMwkaSQ
LQa8xIORpz/gQbcO8RlDf9rHHex/t/n3917ulDo+grPX+9L8xuxlFm81yT8i87J9ny3PrgfD50tf
zl5F0uZxzDMlGa0lhxV9CycTPvJCxUXsSIsVYp5LbsEY7IYaoOXHisigTnGsO6yp8l/vUHl+zDrp
NedUtGtblNI6i0xI32dLwufnyknXuKkGfIrejfTol2VE5SdMw+IR3ZbO4MJPRldNWYMFwqffexz+
52qxx584v1qEpRGPwKgxvLIzmrui9nL75M2cxOOfDqbSRyz6eyqkXRnY3d7+P2h5p/SsVXsYQkXn
KP2Vo8tp61zzpKCzdwqqLwcR4YSZDdEu2xybOC7yeCfOHWhDpozjrXrSwqVe0UxUouQghG0aDbPj
VNcFG1M9GlepyUJUBYeHp4FBmNRvqIiuH+tcyKXr05XTjsIvNYRUoBSyAfva/J0oeIUu1oWjEt/a
DmhPynkyppHALuUNZubLtAJFjpE1J8VZH0+j3jbupNHPQqplmU3vZ0FnDD3H6FALtk1QJMmm7Y2P
o8ndGncQlkNZXuxJWS91kRYUuJnu8uLgBwnnvQRL3o4fzZyIrLYCCtHfFDfCgiWXOOFhkjW9MRDa
DpxZutE3K63x/NBewUV33p6zvYmD/8aZVAmn65Kcc+HuE5/QfFDihjKlGdqbEB9CLPSqjUQvMNve
ZC+4gyyUqE75Ke6lfNwGM5xxCvRIIuBFhKSpar6g99szDoUATK0sK1377aHHnR6qzi3VYPKNhYRo
UGbueEiBDYtSVc4luxQgA2jhm+Smqj2pyUF5RASGPvZPN/9u1mYRDhnJtpI7hwmYccJJXNlJE0jD
FtzwtQKPYoP5FsKTIw7NsQTVyh5grlsx+ke6rHO/ggEHrHcCwkqssaZ0M2dXhQYq7aAXvolymV2Q
U7FFGpGZxNWkRuSp8+m9BsggeF4ipS+qKVYeLnEC5tXUsSJsuAQXE9cstU+gwHamPO8neatdwgDN
nlmZ9zUS3oZlyggYnRszGwszIbLVK9F4UsyudbqpWG/luNnlkraAytlqzAACctcpzm8QgVVAZbla
M3Y41Onz8wXKv29zL+UufZkthqG4S5ItJacymG5iNlGY/prIPESGKC3x3m4yx57CbTvYoCuIAzPx
1k4ompy9TVp46lTkh3mTSE1FoBGEuKjM6KpHW1D5e4npCbGCuaAO0G8e3/PqXQRzTH5FhrfuN8Of
y4j0oSo1eb/KFNbj6vduWHYQ/+72ADCK4bL2peE6zbv27t4NSyjI7fDbpRXP3mL3un8yZ6iEMv8c
Bwq6m4KKF7diSZuUXFywlU5Sb8aSo4HxyYOUg9MNAl6q9/cFBLTgpb/hz5JdsFcOn6THg8GJ78qg
huUOM0ACjNLbvqhDnuIZECSLiP0XstkyHLVKPkdFKnMRnSkGJPFUtgFWCDSWMZnK3SY/vDToXpdF
SgmJpZUcGisH+66nY3mTVw3ej+G4LooSnc3wEDxjQh0SreV0p2e+Ci4Y9eL+z78T5uIXaDxFhqKv
zE869Bp4Q+XxVhmEIX6d6I5l4RlXV7j81m1lALzPRPFDnVqDGev8UN5vCq/+CNf+9V7dSU8+hx9s
u1uTyn2CxzLSlOD5TNu/R4O3DtrAxgVcKorxkzQ+70hwipJT2KBR/BfkO+UJAmqLKaElq1U9K7+B
cqG7voCGASsWysq7lFd31VFp07ocPdlOuItJKyI/GETjBdUwVRvpn16+DpyQR7B3BfKjbBLzqexH
l+gvHTwH0mm3KYVWC38oCWE3YBofdKAThWvyfR+fBmqmx7wyYtg78oyeH/Qfp5wCAVQu0VDgOwUr
G1FjxOaUYWydCY7OPBzsHjOZ2RcpaGhdFYAtxXVTA5EpcFPu+5dKF9VClK7cf8j54LcVWyT9QhV5
GM3JnPgkaErfWVr389wC6v3OX9LYEmiwrV/YmZtL6URITmT5XmKudleyxVDor1OzLAMVo0J8nXGW
leCeK6sOHzM+YdaL16jViNb6kZq2nJ7zOdFI8V0Up5UmjCXOnDNfkHCfA8TPxnMfA0GMdcgtTJS/
rf2ZgXKFpNJxP+FkT0b55nEPcnaJG2dAZufY5+uupcfK3zmlcC4oWFs9e621CAzHpF6tE73Pba+b
ebfqUKX8C42g98gPiImea9b7iPqyri6LEv0axJ93PJKRr2gNI2ebSgETuBiB8MAKSjzGN+rjfWfv
4ilZhxQZ5FU5U5n2AlbH1/870JThppHcrX2dUuYr5Mm6hcwm4HAyHESuRpUrYQloVO7/NscQ6Yk6
wTlEwZTpfif0JPPHUD/iFzoImSELCGKsUnyEMobD0DyWPdNzC2Zdq1tVWRNcAI8veMQQdTEX6IJU
PKbaQo/ASE1yUFn+4P87y3ImnyUBapU8xBdVBYlDEN7iHNlRigYyjxZ+lo8Cuy/V5i/8x+QWtyYI
ZoZBuXw8KR0LY6PnHVWck++FQPRUii84uMQZaZRCxI5QpYbhLZQTM7fe/f5TvlMkWomZJEmBbdHI
LzQjnHlTBAbGpyZJNZgd0i68+q+dt75fLXphoM0S0lNgOoCNZpwRJTF3ffLlcSdu0T49fJ39wx6e
KubFXHShr791RczNBqdJ+M/gYJLrVg9CGuZVZy2xZu6d768zH0nQrxoAkF3ro2SMqMeulvVmysfS
4QueGaX0taFhDCS6qXAryguNu5xwHrhL1J4W2LOy1E2ijhEwA1FdSaAKA7pVEbOdq52298QcSXZU
gaJYijkjdO+WiyJgtyB0ohAHa/3EUSyh9aZhpoJNHWI8GP46lvWZpLJ792aAoPh6ZRl2geE6UECr
2GkHbHCZmqiy+D89H/Su02WmHkK5lS/SkZ8OsI1nO/fu/SZjUDg47lr0NWavWRSGrsxNug1EXI1r
JUN3su4dXyKaAebu52Rb8E0tgjzS6kQQjx38tC8pVsBE7068Ixale3z/BjgKFvr5GErnUNrU3DYG
MQp5wFkKTBODTx0velMdA/lCWzj/hWnWqbi1Tv7EWaByj4ekZwjHCeY7O7d8N+twBDvLG7ZE3YpM
8JsabLsxhjgHAz1tsGO2z45I8s54mkMA6D7DHockvtAUx6ZbIqJT3sEfAoFsiUP/U2jh9G5Q981o
lqN+HgNCRq0fxw13sv1SWXD1qodCdYuJZHTD3VvRoxfbyKbLkFcXR29qB9C2mRYJPB+gCBHcp+CB
wr4lD906z6182cah1vjVHFEMzDUQPBpUGMm7exYQYe5Bqpz89uWwqzsycGUTX5pWb7Gaqj6zPqFn
1ojrsV5PLT7ZLOgcQRemn7EDgbYdmyKBgMJoOP486KdLPKSqRKhpKZRYOP2VMukfBLfYwzfARuie
6AcA2ECx3eOujmM0746czhQ/Q98Z/Fvy/Wy4Ku9QhqeAkfx/cVAHBgYdxLhVazN+TsNgqAWAxw69
BQSUQlUxoMYKNRJ6GAJKvY8U8NewahNyLsFUS0GvZC3yAhY6Kas5bHwMtutVYfv9yBXoRC3tvuoU
W51Rt2IJsAm6ElX8C7Mj7pgtl3yv8tjB/djU0StPeju4rnI8m5H5fysdVjxcE/Vs0g5wlsQx2SPH
zGWKHPJ2II7paxDgzxlv8TwCoosID78saCbHrYD/+z51FzTXsyksb8KNNmIeL7gJfwrpCpm9XHKX
86nCuEq+LlEYH+VzipWc+rLx8WEO/aVefaL2av4xcn1KFfW/jishAbw4lK0P2OXcZLYTZN0RsuPA
QhFJ4LGm+IfvB9AZUmQRNSelI+6Ywq83EAl+LezzpM68PCyNWExGI1ulyQv2dt48kV6ecabhEHuQ
uK1HVzKaS0Pa23Yp8ZAcrv/h9o3+B7ZlU0BwJ1ENGlHKRoPDIV7oOWubIEBOeXy04QUGnQs8FB8n
mbfkIlPgEIjJAWWC94g/L4RrY8sAZ9BFax1S0q+JYf3+knMMWroHAfvm6rl9VwHlCshi9Bc8yTA9
d3UTwFRof0lWs5msrmlr6/rXdqHegyXkBy4wE3n0y6jx59ChLHVluWKZuWXFcIDNQvsjrFyrrwkG
4A/6UMZWyNmSc8rZXWGIZN3lCzdd45lrCeq8ACDBMf0kFUIli8KbjDZtijkG6DTGGjjril0BNoL/
pNopBluWAdIRkRA6dYJF6FLvzWeKOZyVSZyWTp0mMuDxczBLSCeS/oFGtISTBo4vFJMEbUYyIvM0
WvADeXhOU1Ge4V5evEz4EvYjVZSBNjC4uFz2He9WOGl+HEDCOUeDkTOxw25OHYeXWV70JAaPPdWy
9UAHwgsy6iKno+aiNojvXcud1oKcYC4eEIu4HW9yB210DW1+abQSOV2hhQpBb8qCKyBbYMk2Jpm2
tfHpuLF548WeK9VM7Mj/aG7198KyKVFzDOFZ0Uq+vgXF+pRYGp7IDu5OOrB2pJlzZMrIDFd9WhUd
KV0rZCWXDwZUu0WvhGGaBSE/SRKGyTV4BhtjGoX3g1SLo1TD0CDsbHfU2orlDP93p7kzzPrOzbtG
fDolF+qjhhiUOyYBudig7mhUj48uagGOd5baUQfaE+jhJ2Vq27kfc7ZVZ2oWKHpBjopuioMLh1g9
UoUvTpfYxdjYer0oQn1mjR1+ubqthuXKoP8B2GGE5n6wxb4UCJ2FQMWuDvM+OKKSG3rk7RlKddAe
DuxUpMt2unOb/dnhVWq5kCv+StA/fkAswsGQ2vQ6mity3qHncOCPEsFH6lrHHtlHSDQeIXy/JiXz
8Cf/NMtvWwHgb5L6KicMbzCNS3X109be1Efl8U7zMyC3kcnpC4YQTQJjMwOFwvJawXhXCyuKy3e1
zVPvAZtOAlDhS5mki39s4MVcQJhmagnql751IEJm6UDNaUcygRDW9agIQ+aRLEoLhrznXjAjCwk1
FBDYECDGqXeBB569wSVevO61enfN9yECcUI8JoVqii8neVSjxnwWenAn+VlaZzMSue4u5eBQvIcm
8kV2GalYW7hS2kQEbSqvhpj/5tOHkb9UnW/4AhnSrBzXpV+dHRZr6zJ7L4NWLBNxEzlJoaOrWyJ0
ESmk09ANBfjpcXM6YK8NuiIWL7yBvBSJPIU6ddvEMnQAquM1I7z16zsK/yqnqeOFuzbFRD6g0+k0
I4jPdFhajwEf1H1nz3CPHFhbxIAWOpAf+V5EQ2q3BHtbI67IJvV2C05zYXxma/oZ467SaKTehZ1A
Dk1oCZM9UxKA0Oi/goQGYzb7rU6wYXz5rOKiFTmAY2a0CWsEpmAlP1QMb5bKojUI9A2kgJFgXePm
V6SCHDG+uu3nSGVhwUodRGMGAIrj36Sg+YIhEOn3Q5AhOB+PFWo7mQR1w/aGtVvcLbuIaOMGbjoh
D3CSEuErRXabeIYpsVN9aesaUD8KvMddtx/8i8xk1gr62NurWUWi6xU4IMC0k7e66o+QAE+liL9s
me9FeXedc/G/teioV91ucFbU81X/MIEjpLN+VBOVHAPXoMLQwhI804IPiTgGDqudSur9Bk8GaamG
rMJn1poj/OVKLdha7qLzFfaNoqq744Y849R+sV66SE3LN2upluR/GKGWJuzYMyiQxeVcSoy1KsVo
CXkPr1JpNgcUcs5GMpkO/ioZw1c+twE1eVNnSousVnom48W8+AHJKhj40fYNuIAIdE4vix2r21C1
cxrBEacmDZYAeZTVhQig90AVQ0Y73H/ClQHWtls+X3VuoICgx7RhPCzjsG5P+hdc3T+JKFwj5pcA
tMoSnt5HXPzrfJt1tC9u5BRdOekawg7VBJ6syUU7bekGSfYmfJ2dZrYsj+sYuM/sTP4IIsrAgLnt
druirJAJmfW1q7U2mI/TWcRqBstdE6evMYdo83OzCNkC8nUegc2Zf81V6zmwoihOLozC9H8s2euQ
hSwGUW6LyNqmPGjLPfVTy0AFbD/FGJqDWxRE9SzfRLClrC/cRrtL3iqEiYfR1lEjulESrS1u96/W
j8A0pp78SvYEr5Fy95BF7bI3fy5cXPG8uUGAW6WZuQtFqKg5do9KwMcaLTYGeMLvJSRnvhNy2uGd
DUh5CZAkD4tm+Ct6vwnEKJeyT9MP4J/ttH52rngAa3IYiNMOJUrNAghA16uMo++KuBzTuM9u1Gke
oEibCR2CElv9GSKhCBvRpIsvIIspTpLGLykyx9w8ikD21Y/vmf0Cx/90qwuFaooH3bgw41FdhOUY
mr46NE+WYkotKOfhfGp5+ajHXjJDrjpAPZ4kYIIWKH/PFgAKlCMznWUgg3bYmHUMpzwmr33BMS15
LGZEjxlfmxo7a+iWlLJBuZ63zQb+YryMe4DPGOmE/TF+WRy2sEkkq4pQBPsSpczGUNhY3sg58Bqc
BV0eeRN/pd6iB4H1HdwsCt9qi07+ep4OKy5+8qQgeZ+uW0Yja5tm8iEs9LJTWeTR/2raCZBiwPMG
eAAUXV+b34VfYspbvoU3SQaqVfbXnQNBaDh/ewM+GNYEjDsSBAemphxvcy9xjDUw6iu9G7bgwxD3
/0tsBVZ0G2oA84k0RiVuAL9qea4Pf8qCCIlXfSTRo2uqAYY8xwDkJE7U5FBg8jRAe2fIEc9ftQ45
tlZ4XtVBrFvPUm9RMZD1OS7zZOTTK5/o2yNOaO5MmCBzblSsmuMBPhcxxeCfpeKiU8oDLa4dcDtv
VfOG+O1MzFiSgUZR4d76LFJle18q4v6uvcVuG5CXSC6r24PUfKU6J0nTWlfAO/zN09XcbZDrfrgn
APHlCV39F/UkygLy8xzEE6ZGxQKdsFVBgkWmRDN6EtnIKRYwXN7Rwexs3FrHaTNrtfrhOuPAALwC
nDksT1e73pwt+86tb1Prza/gWX1chPoQqf/bqLpmAZtIpinld+nvRFRIbbhWZGf/U7TCI7wMZn18
NSWvd6OFv/4fG2g8S48tY0wAJQv6bXrL7DyY/dQqTNe1AXx2xS3R97ZlTqd9T/ElkNpevjTC+FTf
L0MfIrvArekGdZOp8c0WbnXEiAhU+ku80hpl7Ec9+bSPrZPBaNP4H1Vv9nPZoOKIr3t+bVe1Ewjs
MFi7X1ZXJJJF0aEPg0yJ+kvFMeA7O6l8VLSK+QkKc8tRcGFtymt6dTAH+E3MM627VBZZl/cliCik
O+WBhEudu7LNdl54PKcg4J0694+AmxVtM/NzyTcuOgKUk+NoKR9+bA3KWOKf9/Y7qN1GhiDNdlCd
wssNJTc5KOOQ5X15FpQIPZd6a45M/ZeeHzQZ7/UlldeBDxheDcbI0ezMt9y0BD0m276I4Avub6QT
nuTPMEvKkWx2Wq9E2vfLKcPc7Dt31b9Bv6wTSBtP/xkG/8+4pO24g762UFe7Utk0+8PF7fV58mKM
1B5omvb/9R/iFgOOxzGnOGK6sOOrVhEpoZKm9qOmX+I8ewX4xbykZog5hDGpK9uP3+cxp9VHaSAl
JU70IIbsDd3n+0JToQUrxYgUVstcuf2Nlb/oxf/ssHK8SYQVRnxnHVOY5OvnEcCs2gVC6MUtLx4D
Mq2x0Q1TjbtpD5HXvvLRJ3MY2rJ8E3m3T7VuiC0yQ6t6+sF3hQFcp8rVeJbEnM+fwC/almK1ZnQ4
E56que2FUi9tmxOt6TZJBwUuvwDMlMsGwETwzkLNQOlBRAQudHtyyIW9WZet9evCASgUrB4nMFtM
Qk+qGtdTlfd2JjJqEE+Ulqq2Yl5dqXkMjBd0uwUV4xgol5sZSXOZ8AlS2/SPLo0DUPNqwkEMZGa3
DPzxte3qqgu6KUwb6GPTdZhNjWIQFuICxm8Bi1IuobzNxAKMclXxe/ABFkemlBGAqAI9xzLmdITn
yZ7/R6nbp/v2/0qiWQhruWQ1x2nnwjud/OoFSn+hpY8cEbQ+XYFqxhVINlst1KMTpRcfRkt8ALwC
VM6kzrxBI2zIaKoyKEEx61zY99RXVfRMFUhqzo7gkmBjvxUYhgofo4TYPz3vNHkS0Ri9Cv29uhUq
FenfxqxbllkG3DInlOypDVL5NlyU87Nx7j8R7tQWSl3dH63mLNLYBrEK9FI3L+2fHynxSktEtEUT
WdHNYCpv1HtXaJnUyBVpUa077TaaGooLey/XBmkXboW1ta63cUD/lXz0H+wslinXsspeX9TmicUc
z4PhnYqPnUs/6dY8zQLUhwOOi/4U9JXF25f7xq3csmgIOmg33+97AL1R4oUZOpPsUEQRTsgpH1Qk
dAd37JiVGgbGXULNCqcawDeAYNs1hIT9gOyidAz0oWzGswiJnI4kYkptsFL5jMSH6o7HGu7H3SJo
3VH7AYNBB0b15ae7j2XpVreJJ5+Sgb5jaLcPMqgVF/UdRlrXq878HKdrLBxfw3gmjFX9cHEnwYCX
WeHdyRuPtdb4j16eWb+IIcNVHKnuBrlA83vv+xYPhysPSwWF7r5vUJfj6U0Y+0q5PDAMMQExvEXC
r7Qj9xkoylLpxYDcQUueVCOm/4OWz2ZUz9PHRxYxdC15Mv3ttPn237ulh3eI9MKJT7s9AdG+HT7E
dWqRzQTHUJe52LoY7S0UPVq6jkySH86mPNvWudi01mhIsbxgpN4JZ1QxoIwmmMiCxwp0hqCo76mS
vKIucYNN89kt4ZR9wyi46cMJgMLOfwklHqKprSZIjnD9pIXfMbRRLMdZ/ZbIb7N5jOTmW7i+eEMs
dV7Enz8GR6eoeecPj2k/swr/xmr39KgiFy3B+1Zoq9/7+Z3X69DQWem6TcFt43PS86aVdITRagqg
hGF4khD8Ta0Od08lOoHn5Y2ADGm2F9mGt7rO9Y+Kaetark9BfZOKX7fCzcWY4G6gqKCHLv2+vPvF
fRGfF0f5b2EaypwVkFB1UgPESm0B9+NFN1xsBotmSPHM5eIQQrK4ZgzLctlXssMPbievDTESwu11
eHIRnYxBlwSZa5nWpI3zM8tS/xyBlReJZDR9nhwZlshhX5N6vi+oKgIXJBOsdU8HMcpSby9ew45q
3BUKiGMCc+OvYxe99EKdwL5hiCUQmXwFF3ENJAQRdDR7vgWw8nb15gn/AHCPmfIUypY3o6bN3tmE
vy1gUXHBlnVOxbQDp+h+Q+8aLzYR6UXdpaGsLAvo1i+4k28kubtsHPJDOl18ZGMtgmgoV6GUK/tW
ynoE1+Q1D75OieXw/I6CuAaDBwUHhLfC7yL9K9i7oO8XT+Mk2VeYWDDpVB0IXH4pTTHdev9iZ+lH
0Egh/tAot3KsoXk8iETTlHW+QGJwe1cuO48nHh3YslReGkUKHFDL2vTJok7pJoPm+DMrLExHN7BA
rJGWPoP+fnKVJUjk4ahjPj+SV1eRUqvwJ7KIIpovMmMKZfiSR4FowglgW0Ipb8EJY0tFZUGb8fKn
6D1sIN9cIFIcShFldA/V9z7bNdv8YJN2e96iEhwoyGktPUKceIU2n3wB3xtnGGGjLBFlM+J8YkVU
fOfrDb84DtqJbTjOoRKv8ubKo2lFH0f/FkttC4AtMnBO6RVKulNmLQpRhUAoUyuFkKUF/J04/DGT
NxTstMf5g2TMn4YWtYzCS+XZkE3rTeO8xRVYbSd7mN9IRZ4vLAdpGG/Ja7MzorWaz3kBLpEXX/sw
FeqBhK9t/oXXw1wyhlBtUYpz1OeIrVpCGr3nfec462PuN9raGErwUeOV3Kt7xTK3DRoMj0yVYa0o
ZC5Vnod5pyhqZmMhujWO2VJWFbm+GE1JrhpInhzwHhVAnR64003VnHrxs01jEIGi808qWpDG+N0q
KX4UoAmOOgr1v6TKcWjFhNmX9DGFwq8XnEpkZbru3nLViIbTRnoxzPFufhLac1aBE+uVVvCvXd4P
phtpOCXJAqqpP2PF8yUGENXo9M11bdNPOzp2Ljz7awHCIdGn71TiC55zLVLoRgj7/STuPw3Odv4o
+TbJVe9120XMGv//e0uO0VByQSWrDoEA00El/yvMjfakgYdpOwW4G8IWIS+IVvU0u++ZCgHFCzFI
WjYUZrXVPARhJWDdyYdlwKyJqBfPSG6wRfjp0NmOzXk8E9TjmQHA1Rh2f7JRkYG6Bl9WJ26EfyPq
uvNNChzMW5CWTBQGFTIzQmJPot6nBWLo7qX3gbhRR1l4tI83Ah4Do4yGoOmoTmRYtMSKqvRFV/P/
sV9QbUZ3K2wIvPKCQ4pOQQzXmTrRORRMG14Yb91E6uJYe0C66BhTMK2Q681IEq3Di+NofkG3MNg7
UYlkfYVRWy31NzrSEhwEmp8uognHtHhsbGWDt7KOKwIQLu5jFlRWCN5hguHKLutgrlp7u2UQ+sn9
5ZKA9gYQr8BYMORDmimu+6zvFyZQNF662Q4PHTpsq6ZHV7K1W3cr+/d/Eh++pWbP/Vn8SoCZj7JS
F3QRJG8SxSLSkAGgdhrbqPjCHf6fHdFvhIOBF4Hspe4W+12765K001dfgjTQ7VGjLY3QSfKzRc3d
NajWoBiRMp5xKBElx72FnuCzoh+8bpkGK0LX+qaEoowAGdF/1I0NvH4Y0lbbslQs+DOg5hzwzTjK
m1tDSdrlh0Br/DUEExXvUMiZhe2d1nfD7jon/stb8DgszHKvYWJLiPgSoQ3kZEw91aGqXK7WihSB
mes+NgUoEp23N1QXGFr/n8z2gNSwbZ3mOgas53ZwnxcbEIXXFDUXX8uMEKtoaY+QNscFSJ0gBa3p
JsWaKpBABvQ35zNBMOcxUpjFH4NbjVlCXz35CuXU2Mi1xgDuRvzZU7eLI4VMyjk1crxMnmAjnbj7
8tQaV9qnpJ0rhHeQEC3u0xBwayo6e1gwkmCXCusRH2AFi2q3fDYq6Lb49TKl4Gsg0OYKyMLwndkH
6Hefj4m1kp5b/a6nOnQVJE2R1aUGZy9nL4utn6wD33B84lr2aXh0nmvJmiG92gMa4BTAjjCH9DGF
Y9Qk/s84Rx9S244Qy5V39CmA3efe1GjxaCUzqbHS2+CEFB+AeUT5lBfxbVpvwcMYb3QzC40Cb8rd
V3ZLxM6J6MD7VDbzDzGgJIxYQogeq4Gr58oq2cw5ljLdWjb8luTktJEtH2MjHEQ9YPoP5cMlSQ2n
pR1bPTGG3N007D4lpxOV4g1Jk3pcbEVWPOrPbLnEUKcbXAR7Hw1uAfmaQPhz2FUnkBK00EIc5h8e
dNc6pJIXbFKv0Xic1Bq3ZtFAOCU45pamqwe0axq/RsWcU+mNin1V+OBl2CV/ddAT9te4CWxmQ1NA
ECiJwQwYFOJeiEOcO6ALVe14qcN2fkr8hgn1+P1tuvzk2R8NXkR1RuDyewbK+0J7C2i8Yv5fws1h
yuEq78JaQwmf4yzVTpvLUmca5uuFhIcUd9CVXyrSMe+8y0rzuevNakCT576jSrBj7fdFF1pHVz/B
29ChVEmolvOiad1cbtBQ3L3/7ekSWrhSVeYQLsviX1FG/yZuoBKO5tEDOIfascm5iJQkbF+u9Xm9
dWdqkaOM0dUwYltqh1PxIjA99ryvpDyL5DP/6u4UyQ/4AURiXIHUPJa3t/Ox2XXrv7+MExX1LF4/
d2FVn98Qvt9rJMOz3WWKePvfU5dHQdODOQDxXees8fZvW3SIzFHW0fKiEz4afQU5+5vYgAg4Tjvc
Y/NPv17bZnefGO+g0h61nLKDgg4ZUKlKzL7ui6nZJuYncptKa/WO3NrYpgqEc/NTeiV8L3C7lqqj
L0cgeUJjfwfDYmuloF5tICmndIZHkE8P7Kp3w8tlTf5FMzSuyUQFKyuxqjGTzbEfbqGuaV9LGMok
m64QQg7x2wqG24zHYvaLgnNY2EDO5PUvwzp+sIObywOf4xXCoqqIbzQO7+NQSri9bUjtfDpH48j7
xOZJo1v3CE+3uOY2kkZqQX4YKkesY1brptFZAMZd0d1yaCJGaqgR51O1Mb30SEzoBOa6WTjoUqP7
H1rfS59F9WzdVMo+gc0li33gKOYOx2goQILbMsuBVf8PI1QNYT++Vww88L3rC9P7NyokQBwmLPU6
EfSSGmQ5IwCN+jYmKcJSf99RadItaNHjIBXV5hYEOWMIxUwVSnTbvGPLxTi3BQYtVzm+nwzUAApx
9xplwnsE0GUKW4SNUyMzVjsfSt8RA1czBRzN+gY8Ah57pTZKoL/x+x/XdfDPK0aUJhGlZ6xgJROg
zC144ilV9SuxCYsr1hS9CD9ovp4R8HO7iuJ4/EZ3C8/O/XKh1HVTpwf+uZWIlE13nNAT/ZfGFQTZ
9Gk4qfYdvR+4OPD8fqIqKqKQEM4jBxu33oaaNTbyfEC+/pLMTawDSma0tGALHUkZEz4KqmJ200Cz
WKlGHqbOtqsFhsy0GHPeRGKxL7csQ1F/GfzxPMtgsoAP7hnmF/qRW2In90CQgCgc7aX2w0QgcYnr
I/VTai6szuEZbMPMIEy9Yd0Ok/vJGNE79L35vWOWFIA4imyzDU5NYO/Fz1R26xb2z6P6UePLY+tL
4RFZfAHyfWM1p4kgWJ8yENYS74Msskiv2vJN3Q54oVdtjgUNtVGd3NpdiWzYuRrabqUj8cBub+3y
CAhpPDTh3lsMUDh6KIkzJDeHq5PpzWaDqVpqSSmpf0CH/jA/qw4B5C0oec7IjwlQT4bxdl+Nhkdz
67wHB14N0wcAMzIRtZrebHzh2biPVNpoqiy3FU5s0D2NwNtvOBrIAywCbSH9IAq5Rlr3yKrcvJqt
5UpohF9lH07QBW8aH+VR8s5lZk8641nuvdW59ABYOwjOWzbSnqfBGpDInjlDhCCLysp05S8UgHAg
AbCFkfkgxNpMxG7r40jhzFFYxHgNV3TvXXaWOOFLdazC6c4vst8AO5/49JdWjelDtGVhqVXKzc6m
wlIhcbtHRza0qG9Pnua4x8y/LlbFxb2yGdBB28iNqu3CClho99qHNlzpBLUD7qmqFSvoPpFoYIko
E1/9ixZNJOaJOHv2Z8wV9XrIF7ovc35h1xgXfY7euI+TQWjyf/8TU/od7gI179DvF6/ep3BQibvU
/uiSYJjNYj9W+BUiXiL1P4eMC23OTlac4h5WnynuziDhZmTe8JPmTWH1rckGZNkuvo62sL1uSlSI
ETZIm/s1FYYgoMErHyv2asObvgsvg0hj3dmPS/H5cFjaQ4VAGylah7K5mKCsIANbljc2RAMKY6WV
MXqLIQiQLpEiCZrH5CDVmWPluH5V/sV3R+6IDSwop8GRzAEjlWaEF/ermA3qtdoUBkKZtaMAc4Vw
xDmt2pM3IO2E/ZReoCqyZe1LK1KsRgbcXEa8arh9NKYbgQWCegyHuKH8Pb2NNWL0+FbrI1PjUJDA
GlBivUfDeUtuhzWL91WiYuu2AxvJpClo1g3gNQisWDA4gpwbDaGEUmWO+5DbOuBd1Rg6eBQ3RxTf
oDGyVpY9z4DHCYxK26LDxY5dUrksn+YKF7/YIn3dN7uvxga+4m90G73j2TYphi/gTMR12+CWIZrx
0tlPQHvrvEkYuNVnGExghLHPkt5hXnGAfc7/4DWvsVeEbiHtL+x/qq+736VFXBAJe5GkG/xNAteu
BMFz0F2DyF5EkN1UeA5eG/Z/UuVZssYPZjvCtQMUPdWqnoekH5wSQZPzV1OePiUNzhgPis57l4TJ
zU0f4K09ZCq0J5jbS9dWM5i22nqJPmE0R2F+e2wGYlzQKTGAR6SniTpG67498AxsH2tTn+r7jt1j
mVBkTWZ2YNaehp4LjfRkx00JhtiutT8WWkUNckumusJDGBKjPhGRXISDQ4YGVaphb7tPGwQUDkQ7
2TNi1LXEULwwNG8M1CeOPQtWcEdzp7Z9SWrXuQo4UtsPZntrS/8azuthxm6+GNljI6B+XhHwXBaf
BadHji3KOVC83v/new39q0s945VezIhNdiih9X8HP/Ovt2BOQ01XIU7EY9WP4nzUanx3mCSfy8mx
xPcUK/0WeTsCZz61rww17etzCItKLn3Ak0haNYNwzj9zEZHSxBo/aCVqdoElJa7lhhBtDfh4REy4
mCpFUyuuzwhIYQ7T2PxWC/iFMH3NiEXhOaSR0oKDNcBAGqpTHc7ZwX2T2DqKHZmIOHZb1C6gNLBO
D7rrbUeWr9q2UomqM8jrZyr1OCt6fzgJAUTvPYexQls0WX6rzPvDZfDJF5bBD4pb+vN6vXKtADl+
WIVIiQLIHK15GNjtf+WOprcu+oBKc3BDdyVyr6ZBCGl2hIYcXmjMzAkbHCjYWNxFu+7sTuQ7phJw
MICTVLylC4ovHunqtg7nZdBRzFcnH/AAg+mbJuv+T7mUlfbXS1nYwMHWN+bIZK9crPG82D8oiaOu
zwerHOof7SVoXn/yIcJOqYb2/MX8bUEQIcHS0uRkETJtjN4xCiVdFaqwcRYrkga/mAiqFKlHcvam
NumitSTJsXlAkUS8fBI9tJCMA/ca2O0M3EAABkHRuxCkEYBcX8y0di71vkr9t84Y1kBmxc3U6bJ7
eN1S02bgdHJGwz8E1RP1SOwiWNiNZFaOp7L+04RM+0sIbRfOEAuL/AqOUQ3R/yc1lVA0Upxb3aZF
blD7TKK/LnRzd0TPrtSyxsUxPfo3VLO0xkFFu62qzPMPjJ/EIZVThGIr4iKmyaUNBhVi4c4/GML4
9YUkn525v9i0BroHw8PPpI24J3Z0AjLyi8xMoikgELVmaSsv0Xrmz9B9FikPTQf91GIVoHtCWz2F
/cgBi5Ztz0HZEKf5LP0Kc0ubIOLEC4qK8GxhaKVxRJhCbqQE0vEmlzzjVYf0FQHs7TGSB5Kr+CEI
jrqPHNKrNCYJRijz3g1xR5iDMWpN48aM0mlc2dx3N0ClnelqzIWkfA3glcbx0ad3nsdobihCWVzF
KGUXfk5Of2T99utHhydRrr2e1uh6NceHD8Kf0Rf0yg779SPNtk97gl4SHMMSkTNaESB0UTHT5zpI
SqhB6FaDr0s/mCp3j5FbTNsNO3X7XVPPmVKZ282h12p4JYyUJWHPadj+70lX9XhOGCHFykpjOMPg
5OAAp7aVRHlS58nSW5zovhVAQfaAqmXMqdmH5QcX/s4yM2MQ3sW/swOEhOIlAgiYVugEsJUB349f
++ou7hqL+LK2H9N97BfiWe9UQ/c7uqhz89Oh6mN1CeDSr9cOrs2ndjsAHVBNRyoHR8JZvKHWH4c7
iNAIx89dEkXdYpKTF94cOkyap27dWUI8uvxHdC/hXXNQd1XogCQbqB356+neDxUlr+lcQV5p/THv
Wnz5QW4Ue0O/D1bYRP2eqxgZZ1WRDTVwaEXFpbaaS6ssRCxRDjGFOPfxT0SUHtxVW0LBnbXTR5Ef
n4GViXn04GsxNgtfuGYhxD/lRbAwXEBVgharbv73eRW0NL7z1nvTyg5+w9btR9VqXIjo3IExXQ5V
hOLPNppbcpD+X6zlEQuKXAihm2aBflvn4/OG3N1ZbwW/oKUs8oit/90/QLGIn+SKsV9q9od57EWe
oY1AZnVQvHE32SWkjgxYy/JqUaqSkgdhiMFaEobk9FbqRxLbm4bAMqFAT3Q/HpgVEQiBG+c5zns6
cnJkPbJFfn5cUOtgHgWJCVGJVsku2bIVOyczJga4IsgQuNdAgQGQtQKcJANL8kZj4W8MYmImWOC0
yenh1hJVFmIos6F8m4qk7w4fGwSo8aFZuLSTiReoZSr6koLxbKbb4XNh6v+tz0T6FT5V7Rf/5dqC
dWO/Vz2zy+o0lHVBlwtWMrKYk6IZt0C4HLjbOpXGNN5K1OkNzYxadczJVLXC5AzXUySJp95Mqj9P
XtBUTtSovbsgu4nbom4Zv08S+fZsNHwyZY6cRg65LIHAQzPaGrcRt3JsUB/mkkOVW/rIrDsxhNkw
0zR69e8Mza5IZNJ1OpcMvIAAr0u+RnUCXE69y9FogAKYR8UkaUV+OCJn2OlnuOFG+DAKLxYWqJr3
SXpmPp+xLbpNtMUFYXPeI7fxZdVxKFSzxQJnG1gz+tTcpI72w401/ahnrUOA7SEaaOlnF0Abi/mP
UomRzRrsT2h9NIKHcKI+QTApqQ0UAsjiemv2vqr+dPloGPNJnnvP0oE3uHsaw/nA/rrz1UW5lRtK
VLQD+J09SOUynqHY1T7SRuqCbUKNx84ObKRkHh6tA6fclyRC08etMQrheYFyZU5+fzRaOEzCSmLd
woBykAV1hUlHhzOyaTpoHfEJ/Ct7O897YNG8iHS1wL/aWmBfG6X/zHYhTRxZfZ4NPAZoVYwQDKZO
i8oCT4iJtcyTXLKeglpwRnGdVb2LKzri1tJfhBnmiAqHQn/gY248pH4W13tyOymy0N2w1JF1weez
snl/NsPJX1k7JCTUChSWn4e4p+ZhFmYY/pomId5jY16rthw3mYWfH6aNzr8+Idm1NwX4NVl2Z+r2
mJb7CV5+6opqIGYOH01UfT3BiWU0wMIaofDIlPX/Ej9OI96YdQsba96i6bIoIR5fzmfTvQGFS2SQ
3y8MhIFmWm1ZO3NpzPn0IUZz69z9CMRU2WMgNe2+feJsMzcpjiDi/Nlr2H3ZzgLx1FOB1uk8abEt
2hKq7w/NTsGa2CLxHR0C+hCgF6JqfbJzR4ZpFsrRoYL1wXXt9mF/0pgFSjTAB7Y5Mkf0pSx3Rv+G
uXGHLJ5QaLaV5NHYWTkOATjYPrsnML/QVkiJipLRMTXNXUkV8XSrCuEHadwykgXalKskF58m8Rfk
s4E5DzFQm51jTnBkg2l60nAqT6D2T2UFkRkzHmxJim/VF2EmjKjnTqkJ94f9sskb2OALcXTC0f6n
vmJ6O5WmR7HOjZufQjeUdTxXh8a4QN8XUliymYeJXbt4B6MIPkFgMT6wkAH5bYXSwvyB8QmGHoA+
mfLVHcMPt6XKI3PpOj7GwsJBUwXzO9QRrzSL3iqfDf/BQV4/0Y8N6+so4NYgevHE4Z0dvdeUtO7J
V6FlVqWylvlFNqZJyhCsa792cDwNAF4SxJZShSsiPuf3XOSEOWdx5Y27mkaBQ/UM8xPdvDoXN4cC
PIBpVB0DAQPwaehRPyeslAT8vq99zE2gu3mZmFwOX2RTfGtMUbXrhVVybi/92VNSUYa9tsJFYt8a
CFzX+SE9Qjo4qQX2w/3QhDDR8tgzzlJKKTOMRTALTmQpzbbyFgZ0duLfg0v9w6+PbxUt40PLCc1p
93kftC5+7nD10kDvo6T4EgVWQhbq7w0xCwXSk519rZvqCrfuR7A9pift4OhHOplCznNuRXPk2bjJ
R7mzwJqiktLsxiZLJCmLYwF9B1/RNeAypjwhuUZPwgXO+QRn4HH9vJLgoKYSaTdPSReaBB1bkwAB
9ik6sym4wzlYd8cfR2GucTuZMUN+WyQrJfif5Pya+924wIKCk2lOxaJ1K3W9kxw/x8IXybOkvdRP
4di3cImXLXsFZLVPc0epguj6xKgRNOs9QuAgugn9Bu2WGKm4afDXjt2TOV5YO2fpSF6lnQ4HqxWx
h9FloxPIsDyfHzQP+dkF2PuD45Fwhm43C0E5ktbwSSL3P59mdcsBfuTUuJojYNEOW5UO6K73Z3ep
gOIgW05emsm1Xhy7ZQlLAQALsSBbj5AOwmKRfBHRwxzxaRt1w9B2nN27OUlYsIPEniIBJofljIsQ
RqQAEVN4q9bzAfBFkbjC9Ecj/WllmWaao3hRE/hzTRdoD7vIQ+vzaaSamgTgTWJ38XMQ0wYL5CWC
Nit3BMPvqIxl6TfjbXi4eXkEoY2ltykthiM6aOQ2JGDTEnqgjMmR+SqZGzTNAppkkix4MB9iXhx/
zqvFxJX8bHYIYORHWULwkGwQfRBibxbUW+6tLjSItDM5VrWXuGu8n8qUD132hYqDvhbzASFZ+n1P
pJNOMazIO70v5Rn0XYS4MyUxYWhuv/QtEg7ldVoZ7iP5pNnVw5NyJ6YXaqKFT+sbniJwx3PjAXCV
Z6NdAQND3X5/0Un6ikF9nkeMcHEkKjgp4jaeU8jcxSkeWfKESH0/8504ZJ3DWg+VhchchoOqb0yO
BBtisnPQcQfVdI7sc2GqmTBA9BsiATfWzmd9JNrQg5lt0/C0u3Pa0hv8q97rpBKAJ5TBaZATTNWF
3P6nB59nKiXJZeImDxrwpMTgcIQo/+RGMTDYzoWMd7568uB9tneddddxcN7CH+jYcViWp61+K0qS
0CrEADhbPq9HPfHViK1S7rSRV3RDVQerNwJJpoGdTr6VuXa3A04P3hzShCzZoRlbWtsrl+gkqcs0
RWNwT6YnmfAFcVXA5tJZOtB19PkL/cSB4YeTqhQVX3qHkOeMo/JPEoU/jz3waO3YnjN3yWaXHeVV
+6BeBdHAAjpSznjnNFnsW8/EbSQL+/yE/KP5IcGuqiBAcdtqASoehzGcZRpjjjT+rqL1AozqkU8B
aNS8FGf4R+xaKjx7/Ta97GFnCM7u7YrrcTx9FX37SJIiLRQ+zM/hepN4X4m5IBZd6WIDIF3KRAk1
Q1SpeOUXy9M9G2ZFTksatGdqW+4QdjIxJLlgIm2iB4itmcxHNJkn9VAWY4Bw5BXBh6stDIKpEyC5
O513X/sPxlPK46/Qs6lEomSF00EJBH2ZsKfJe8DoQy/o8KUUbAqBJU3R5p5P1L+fSUYvNBK5+/qj
iyqxHWBKQ0rfVf/9llLIrflM1aRDh/2PqizbsyP2u2azSdDJORxO+uLOuLTmqgZG3LB1JnHH1F/Q
pwtokdMyM5GY1B6Q+4AgvMWCimK/0MzpxHUognIiVR11obVU3nYcKFlvYhnWw5KM6gmlQ5tlaHKo
01WmM7wUq7SVV193pkh/2C4v4L3ced9oSAVRoV3qhEGANjmE8io4pz/xl52+KGQVb4cOvW/6BooC
BCC70wn4gSadluMpA3YF/+DZb9+JW28nhk5izOuHRd/ChGYrfx9Dk7wyyiS3SnZt+XZZ5HuBQcXp
gDQM22MSTHZne3XhjJnIueV0k/f6r40OAZKEqZnEi+3phgsny7YdLWdYxn4tZyJFm+YkxL1XO7hd
v2IGnmpfbOJTpn3tkw6s80QJKKXFaM4JNm9DKBImkc3oTxNqSNP/kx+scxjIWBwHEEGqDh9e8VK2
hsTj1R/4AwaXSAgvWp1KzsnnP5bVBdQp5oUZ3mXZllf0wpSoa6PQZUiBPHGM/vi1dzeq7WZ/b4Af
jCNv8c+uPSVDoCRRhHaE4+HHPULQ3HiCZsCIsQNyZP7N19iFgoPO8ZRjldvmoPmZHtmelFjwlIuW
5VCMA8/ZQ9oElqnlGi01DP/e8jsO1VcX4GRMdx8IBUDEqXsCcyOSj60lQmJa0zrpkI7K/ZdDXVk1
VyHyOWNQQhavwOK2GMIftQKhKg2mtx/CBIl0pMeNrRoucntwUXuGotIARNFct/i8paQTQfDVmS62
CBt5u5AS+z0C8swZme4+K5y0yOI9JrWy/S9nZI5JtxM+2oykKUU/lnGqJyThfTRa8s+oQTNTC3im
u+v75U62bOSF/VA56waH/y2eny3/E/XMTQYVXna0PJzh8S+/oeqVIgyGSST2tBEw3rxn10U7rtIx
B09WWGZsWybYkoSb43FM7+reJfJc2ssYtdvWIIPztXVZwcuf44fWyHOwp1zPGMJCh4S3LlYBZX2a
IEDPWReOveBBZ9EO66AFJ7+9MojssGLAGZnSHS8ViUhkvHSYX5UHk1lyNACgqD8z82A0wwzcd9HH
F4GwTZTqhcBBpNf5PTQ7zW6kZZ0alwscaTABEIEkZYiGANcChjL3s7dZSGLIM+cv58+vpEzQYYUo
ITxiuIHFM23zTMemt5xYCsasbZOx7nuXOzbP2lAx8p19kJsdpGI1VWsW4aRaFE0mW866OotYVU5h
OqoeSB3KI0X5mEwwc+GnF0bX3PpxA3xe+G3GBTg8Oa5NqzC7pld6aOU9C3qBjpvXmZwmGMcrEIfR
RtvZi5Slmk2sSq8siBjAqQX5S7YytyOYG2j4aI6cQvTiKjUx3Mo3IKo9GwS6NsfzKxBJlIivOfrg
FaEctFxoBZcixInHZcDPB7lSuzKUVck6ciHIOa+Q/BuoR2l4YZ796c1Q+DaZ5STgQg8UbtuUXgNI
utvrsOmI92WTUqkX9ackT7tuzwIVq67D7TEn172DcrIhzh0yPnfGIRyov1WdvrsKRGsvroStVeYI
fKRRm+P7beOrNbZkKzTi9zAUmYkPdeGeaM2kIMkevDO333pdDKy0dMWfDOBXqnZuC84TQrbRMUXW
z2yU6Sh79G40FBxeZIVwIit9YYjnwWrSgghqf8ldTCA+V3pE3y6yKlOkSDCu6BimOgvWAua6rGll
IGasYTtnLfvtYf3pFvb/6tKsA3dkwzUGPsG+xbQeaioiZyjhZhjqJPuEYOT3YS83KIgcnU+BwziY
NYk0HivXQGCI/dcdc4LrvhaZEHagz/lhaL8yikprRTo6UkQejUr1Ig8/cayd/ERC7CP8TAzUMTAL
uWw1PQ4AcMWuxRtToInLvMOyjAM8F2jxWluaVLSEcaz86fRRjF70DkynagS22GOiQhr+kLVIMuJr
DDznlOi82UgedtuVh2k00gOAQZCdYZH/BNr3+RpKfeG5Ql6NjTMUJGfU6I8lK7/vSOPQcTSzW/ys
ubdIAxgCHo9/R0wjPCNnA/+LLiZt9c9muzj79KSma48VnNw76mN8ww4ND5YkaQ/hGWMoJkLZVjer
Ct7JcjsjIvT5AotRF6y7JG4PcqqP2lqrW3eW246POZle+2oZdZczBV+9494yy4LKm+3jc+qfuVTi
Ye3KxD/QODjNc5TQxLySaypHq5k2qAM9AqiVeG/tctp8Hq3JjqeglknVvZDN/0rxtwZF22pOBrFG
AN4ydOF1B37tML3b8bdD3PaiPJbqs8unuH0mf37S8m4f/l7YslfEPsDj6fQzWHUIdrjX2Wvf8kio
wydSKadJuKu0FAtCP/8LSrYwhZ+dpYIVlEYknCLfTqoY3iF/MfVuHNm5Vgl+K8WzOvH57grHA0UL
VQFICUKD0o1XnoXMcBsu+cwsijhtGU2+RfQEYYMzrGd971pxwXTwAFhyw8i6NHVX806Dx+zBScXR
p3nAHXt8dxFP20S2gU4ACo2o9oNl5hToPSIYjzlwJcRwEjLabN50488zuZ6jXD/nmIgoF0yi6+n6
O1Z0UD8p/y8TTWq0DZ4FQiBmLUVr86Kzjk+Pmx57yYbR0F/eXJdQGARDNuPzvMGMPLTFNT8uCxfu
l4Qk9a1/GwduCFl+04HwPnidASVlP6fzDORM0P5wXovEvoHHW0Nwd3NWJ6GscGXiFjn1seIn1mvZ
/ZbkVpkejuqCwiSzdXMZ8YxRez+sVXgBRW5pJmdz36rv548D6xoxoWtB7fhGjYoZJxmvHbFS6Lo7
CCDZbB3GwPKJ350rtHfxO0ii7wz1ZFcpTvn8jTWsG8NzWX5fxt4ir4JJC4J+Oa6yr2dpYZTpVNfm
aC6MCTF6LVazwpoIdkRsIuC/Gq7QuvoCiyb2MEnO2sM1BvTvuxZNziO6v4gYpIz+X3UTO+BmmEc2
vI8ysISe8gblMsdfEd64Od+EAJc90NIMBBSgf51YgbgyXjBbkHD59KwGZGGmj5lMVh45w5X9LkOW
qWn8P/K0d4GzOr5VB+vQqQ8FmpXjpHX+FP0j1h3F7haaR4ziO7ikscAaYE+4bvpM57cFedzkeBb4
oTv4h+UJ3r6RYrYhfIX8ofJhQwZChAv94qkwFjz92lhOybM69YZnGuUuDM2oNWrZa7VC5BudoMVV
5q09xC0lUfH6SYKVZrc7Hr7AYwRlRFQSDBChy1o6B3L9NTchOVHGV8bmI/9sNuWtzuxBrTmBs/N2
vkYMgmmRsi85om/m7GjALXmXfzJSJaAui6mCmRWNlTRs2KH4jsdIxvKSzOP9beJ2XhEuilt4fIWc
g8cqB+RCtTiDPbXEL+kLFd11sQ0GRRSaBZdzfFcxs2NwTyLWt7k6lb9BFCb0hb6mJ8itPhpwCgaD
fb6YHj2MqrodqIj39pAZuGvhyrLYtwKEmxJzqU3wK4K6rKQIgAOQZlGpapXry+6ibpStf4TeY5ou
J8JMc82MpjaUB39IXshHzQdOyv0lLoY7uGCACrh/RWzl3H58qMXXkSdhm7UiBlqqxDdMmajkxAA7
KQ3Q0SsT38UqsXRCAje0nIJwsDkZKwD59sqIXw0yzAO+ZT1b4F7UyPOnr0Xih6J9Bb+aHks+IWeX
1xpiJWCy9NTa10QudaVDO7L5BjEskDsfvvUcyi8Fgpqlj4RSHk0uKCeHD3f4ZdqpwBNw4FrnhcYW
tFblroCxx4zSF1npy6s8bDK62UEzb1FtcgG1I6NU4Y3Y8kaW3REyQo5ZMryJoebF7nILkZf9S0lt
YS13WFoYsOI8S6poSz7ISAoydiTiSm0mpNQ7a+/5hsgsZZaIQC8jSyEA1Lsho7KyQ79L1iIC5O4u
YAs93f/TJ9Eb/r4L6YKrjHeh4S7h5x14+ttmCT1kGxWgejCylyr33gxpgRL5yATNqx1GMllU3q0P
ZszPEPRrg/Jbhy7zKQPcMP1f6dI2DM5Hj/o2vyqwHUu6MNOgvLtZ9EUNoZkclNxMhaawRg0iuJhg
jTAd3rwvgiLhPexjtU9NzsEJarHu5+RWMVwY6TT6Mfwej18CvQpmYtoqb1ghPXCdVIN9GnXmLG/9
3hdLWl62oSs/zmNzGj+1TWzVP90dIWqigHzl5GdEchu5m6/le77vin2P03+0hlzwdMkl1eXY7YlN
h+mvHLVjle4Po1rujKLgZBBPXVzyccpoRFFw/RAO8d5Xu/ApEvcEGl17f+317wD79LWopS6wNAbD
o/cr5/XvyJE2GL6Ph5LWfhw64hS77s/JftTTU5afl+vcKG2JPD25n0VkViIUjR98zg8gu5jUKA36
RGuLzugIpQsuI2tGDinpLzy/tlaJrKRUHlFW5/gXwfxR4td7GTw+GNzmXTutee0Ffaf1CSgUrwQV
Bt4gzxVMVfqEPUOyWY4hVuDtTrw0Z5chocOgfn6xlUAtVYe63LGoy9QEpG5SdQ98HCK+mUV3oHRD
gqp/5d6Cd+Q7LNe6dMxsAY/uEUGAwmws+CHS4fOE+06oX95koAZFUWHsTxqneU2GUqJOHfBUQUAs
ZoB9yYFXIkfw9Lh/kj1yikimIqC84S/OeTnmWIGnEPCmNsC6St0/WaFeqf4TCD96Ly3e0VgZWO2o
hzJXQxM1pBQPeMaVKlygY0LyfgUHq+vz5h9I4x/WFcwPvKzG/rDxG6BLL5RCKM5w4SD+42GoJ5G9
1hykuw/n3uzqRZgM1Q83nMSfogL4XtrnS/JsnHGgsRsWaYYi0Q1jYRmx2GRw1J6Bh9EKTug4QRlJ
MxUXJS/WYJq7g+FEs/GSghn8yOu4hyQVWb2RN720a1Gy1EmINZ8GusdvwU23dl+/UvIUAjb82gsE
ibm1MLqLLI2oBK+Mk3xrkxEuzzynmwBlf4g6KWkG8HcFJN3xhzwzLIr6fFGTpJlOVYIC2BIMg+n3
43KTesaPrgPNzDEceOeQTHP5HigicyaF4YjLJhuySCiaPjke4lxSHODXszppvLiv1oBkeJ2EEvTj
+Jb4y9yOVxDKm2e5k2PiTFXk9iYvHUC4m0CHMNk8Ge6sKWyi4G21ji/xQl8vu647NcELx/VWi+ti
3v7Nh+do6HNDdKy0itkU4c8DGkba7SARteqsWfJMljcpKsmL3k0o2jzsJhBMnQWJ6lmEJZ9xMsZu
WzdeFt+V9TsqrM+6uuATmXK60j0Nm5AL33cfjjkbtZMOY5O4u77tICofBtxaogsaiDC/Sv6BFPoc
hGAGABHiZUiBcNK3c9QrFxh2otoIiyBUv2waumPKpoN3XuiCkyhCxwl4yznZh2rqEH9U0pJQ+O0d
AaKPLHm+9G/5kAZtZQ+ceAMJ++BQEqM6oBxrK6uEx/ilvqDACs3gaQ7w1XVou0QCj5PK+m6OULO/
5o7ETtSDYcgy2hTiTSUyAdeO5405M97ne7hNzFIFnGhUPT8Wsq6JCtJOhcpPYXbMa7Eip2Ol76Lk
2GMdgtqcsMw02ONRkeEQNAsaQ/yj01UhkjipE55OS2030zwKWQ1d3UjSJyQIBC5cGsMEicAuaHqV
ZdBQ2bgAUfrYRKf3oBQFBz2u7NKJE2xfc2Nf8cL2YghMuwCyFpyI0OHsf+MQgs7exiz0pCZNl4pr
UhCFffB5V6Fo7EI6mvS9soVQBtxqlQGqCXjxHZUEoRExz+MB235iUi5d3GaowEkIR7gHCUpOMfHr
58aDNX5vmOMNOH5vtNf4O5YgamGXxhJBQq9oQK4ryttAtHwksFHAYT1coRcgOnM+SwsxQ04KgJgK
bk/XcyAhlpGkz1lYJQIEGkmMi7A9twNBG7F/OPSCnGLRQyzKDtbECMLtIC4mfLiuCZpJpqcTS0KJ
Hjf5J8J7cnBxMA9t0tGh0bmf8e2JGeimVoHl37qfer0WAiALdbOWO2RQQFWA2HWx2pHdGMHgCGFL
zkqs6ejszqxLRDptVCl1/i1Q45ekWXjkq/gmhxsbdWEmQod1uJf2F05wkvkoEZQTQpxlwTDyWsDv
e0XevBCtWOHlpBBw5OW8GSSEOAStd+SzbxTCopCsnm0/RDCZ1Q6qHA5PF2tX3VEMgaPzAs9u6upz
6yxEp+XQlURwTcC3SXqa1yXkbdnFTTu2EvDTlvQe7hI7K+hTYuB8IJq9S6lsyzMct0/Wg8AjOCnb
Oh37FA9xxjPTAVc43h4Izls0oM3GjdgVwloJR6AsQ5WMiOPMk+jupNHFHiOVmEJlU6S6RdfKVUIO
1EJDznMz6inZN1aAaQrSkbTWTIP9eo4CTs6z08VEd17UksMK2PSFfsMco0WFS/CP1splSklxNnEs
3bnApNbNryDafSUiq3EKoDKrhE0qSB6uww4PNcM8V4dhVPz5oOQzXq1+8XTc+xogcra5h0E4PL60
pO0XUNu0rKCSUeoYJf4NPhNLbl2oFkuNZ4p/0UvPOSbUcTrLcDCPs0Qtl0VbddpNY68bU1d8pqxH
0yZmdvZcVkWDBTSelp2okXgZ/fEc0x5tMG7gS2KeFNoB6isFy7r9ojPKqf33WigBlZSk8kZyWiPe
WKgpIW321EH5JydoT/Nn/PGdrmqJ4UdaJwRjMA74Lg0GEdhS00NKi++rrBpJ2MT74Nfb/+wNgoUK
FrylPS3/ruA5+maPMcU8+ax2Kp9CNQRTwq/NX6ze1RTxBvkdHO3I9yIatlTovqUhGdVKtAADrmDX
Pct6tt7W+VHU0ZVckyiYD+ASdYgFjOuHasmAM3wtsHK3V6R2fJV0ZGuE2SlI48D+MjSTKhmY6GkK
3oXmceUAada03PQnAIk+DB2TahgLgZ4mC+JdhbhP3s/CDfoK6NGe5Ur42YowgGGOBywlgbFv0I3U
doAlpInovfXCyW4Qz2se8mm4p96DiPzs2gNPVk1gOMkL3J9JTPERbQnEYG8z1XO7az2EForw6lJS
9UDJv14a0NG4VwVT7EySMartY/N8O78FZldcMSPLTcN0uAIsIWDcg/tdGmNBPGT9og+UGqMKNuBd
lshzk/wJThjpY88YDKuSXPQBpDoUNW257sOC38GF/NUBKKau9G79BE5FwN1SB+3iiIn8BC3uMUEs
P1QddA3vNJ/Qjau70+/2rc/gUSRV8fvQVktBQysFY8EG02QNKd/pWCZGZD61UrLSy01tIb9b1iEf
kxBdS4BndVX7LuTEW5voq3VOGqhVV0Wn8EIbmucslg3UjN8iCX46O/NPdmmrqXrlT+EBo4cETF7Y
PIOhTKCsWHgAjH3vCks0KQNi3ReyJ+wCFzqbDRXOU+tQxINKpcQX/tKB2Tgn/AFigqHX32W9PhS6
AkEuS5dGYZyeXaP/lMWIGj8DWsqNCcrF62Hkui1Na3RjlCx/Y9C641xlkPmnOQcAe1UIOGRFej7A
msm6f9ykPgPq1Jyr4wvyV99X3wbGG03vnqLb31MaPb/cSL93pCn8EZJ8ybuYiQUno/dTbbCJ2qrq
Dsi8JFbmbdNH0NNQo8Lsfoes01Bvr0+wHO5J8cvaUTy+ulhC4arBmHh0LiwjxbPbmgSvZQDR1oGV
wUkG7H1fPTvJd5+1W5M/4zLq+5/6OW3EkTpM3ht+TQxB2etH1Oc66gBf4JQHJXE6LqwzyQUBNCg2
j+wbqo8LNN5XEuqpHppGWGvqGJWN7Ea4gAfPCuwu+wH9fyTeVGITT5mZS9iCGbdZ7BVm72Dc6wKl
LojGQe8lNCKwCKT+582Blh10/De545WZTVuaReisVA2hIU8L6JqXQ4w5q9uIeneVx7DsZZYdhzR7
NIR2GFuvGKT8WN0imV7/svycuRgZNIxvG5DJKhlwa/R7lkCym+sVCbukU7GqwsMATHFXUyDK1kIQ
14oMkBZHFtM7tiijyHNVr3zgchAPlqC08v7Jbf/baay2xwZ/Df3VVmHgZNqOzTUhifq0cH19AWeU
4xEpS5VETnrfsaogWNH5DEhWRubPQ99O0gmtx/n4DOE2laTTzyIMEt0RCyT/6KAsfbp1kmIpD+sB
yT9JRZdY0E6sBU/n2FlRud9empLWjueGw5otnDVwCLxxWp7SUgNFx7HuDxuyl8fvKF1j7pAKjn/f
CIJ73pjd8CKme7uFFdjFS45KT3MIYZAv0ZGVDEvuIP6GV4ceqBS4RD/ujszRvJ5Wy7H62JKm6JnI
54JGP9Ly9mCmZtLDc1VjPJ5t5sj8NX57oBhUZE54RtvUf+iJAzflJQFLJ6brlGbC1PBEIFAZ1dS1
czyWa9XuiOmiA0p/JCk0i/Ta7gNsyb0ZN8z8fwp36VwG/+aR+3YuGuMKsDzpZMSB2aesB2BD46fe
FbD3gYcdxwMI02X8d7xUFAXdCUzePP6cX9qS81Mo0KNS9kZ0rMZhvcS+IMLDmh6U7f3MlUyTyl8K
O7Ny79kB0FcHfxvLN/rATyIjf7662CwiCOmhIxps6b1omjMf49MTV1R+Epp2N9tpbNDapBRw4wou
tnqvU54CsrfvgEX7GwzXHOQMn3EpTrz5Ctd2NtkWztL9ZPszYXCYF60drcOM+0CTyaSZ09HkiPF1
YiLgdbeN+atTS3DSQyvNoVt2pUBA0ZtUiDgeIaKrwFIZMxEqkym5IH77mzXkOqqZwFGbzT/Y8Rq5
WLYWZ6gZlxOb+alUrPePyciGRmb17HcbS2ngo+qIjUOK9GZZKbijBuW/9osfJOEza4Vnp38LuV/L
cPtakDsYIAtskh+AOueZxqlTy++FwJMb6Ye1dv41nHX5RkgHxgNVo216otDuiI6KoILOmvJ/GUHl
EK1hK5zX5Ll5SkQwR/pxhlWKsGJcxKE1//aIkFFbjaTOO4EUARA96jOmLttBvR2eso4Z46R+T19q
hdcqMAvr0FKthoRSl/9t/oxBoMJ96V7XGqkyQTMDwOz9qchgY/qiaV7UeR2NG2vqnLYRhQQq2Nxy
I8BVoUyaJYWkeeGSy1J76HzKqj4+SNVhzd2Wwl/5nMc6CkPwxxGpzqaxDrpeuov5kx4e2sVvdJNS
KHeBFZeWyklLDd/a0Z0/Ux6LlGK1AaetGRmCIqfd6XiZe2zXAKKCNwz1Al5ueVgG7EMN+A/82hVg
f6hbSbPtCXNFTYnZhGTPQx5yqCXay/lRP/IVsLZhuwgzUpstG0E6iw4oMpqVNthf9UFWj3RkJtNz
3yvIexxGJ5lL1ppzvflB8j9BCoFctoBrJRsJmRnaR5d5v8Z4xSawqJVruv693U0RvklWUbdsWV/z
NoOVOHZC21v95dMg6B9ddAUvHj47NWWkq1QrbHEuBjvh0MP+fuFo6u6xQVrrpIl8SinOBxQ+NWpb
Smn945S6MQNEm+ZgYCGnvMvUAGQvWmMUkXQR14+9norwnt9At/SQIME/Uy9lvQbU2RVV5IyWCPHc
ogqIzWm9DyCiBJficve5DFHltOLPAudXJ+eJqCCJnH5t++fv6Ipd49jfymVVZJZrahckosaX8u39
dn1FzroSDaPHEnWLpw6k5TIqrDfn+YThwq2U4KypQRZhhJ44OGwZHLw6WptuesBB79OP81R6paQH
Hlr3umgBXcILpvkHbwiTt+8e1g4CNEpVwKSBI0WlhERrslLAzKvhK67L6ROjn72hS127ZLpnOHf4
EU2p3CKMdxyT+HT3sEZV+3mR4Pa1YDACld9z+m/mMFOWWbtw5j42nuo1HwDSwzwAyxhiL/6FM+tf
pRjTcz8f+U4JtyJYUjTFqBZe6DKwS4yxbE4nJq3GFrusjUj9mYNrEaia4JSgcP7aQY4unv0UXCwF
a28KHEibIchH/LmUzxrBJUC+YGL00FPqemdwyqd0vvl1YLa7j3R8pqtTMFCWYlikMqCcrWegx1sH
OkIWyRqTSj19dZMOb5gYOWNSt+QCXd5euLd14qWrRUfxg0HYTxjt2H14XgnTIZZzid4/6ltpDdjc
chOIiNnoCngy3t2xtC9PhQDDTlu5Thd8RRrYmAXlXg1ZNG11FBrmBLf3O5+uxVThfRHsnW9934o4
Lhv/NfxNyL5HYa/nk3OBcoMY9HvzdDI5dnNutGx4RCAfmTuNm42sdORW6VmQt1JgLSXL2gWEpexb
9t7Fj8Dq3zQFmYmqVxODhevP/77fPfOq4QqiA0NPU5jdhD0X4wqBEbbxXsjmemZ6bPT5ugVKnzOl
R9+S3DAPednUDh0qwz3MQPxFLE2atWm9q+Dog/SACL7nNMe2VFng/uJt+jxhWP1KQmMtncX20FoO
Yya8wH6Ka57My3o5GJkMMOSHkQT8QD+ogDhBR4d010xu5FCHvEvFUBLdEitPIgSduP3TrnsFN9i6
Ssq4jy9Qkn4aGeP7rt6cj9XxtKbYeHE9TBXrlCeFfQQpkFww4JOguq4fkZK6912IuKZAuGM0DUsd
dFj+142XpGiopON/ERawNecvfYpBrA4J9obeTcKWBAB9uwokObV7ulRjZ2YLtdJNwuVSurmS0Wok
jtBB9LlWDY/Wv1e1z5JdVl+xsWYcJA74eSj6FDiVtCDGJZIPbkD98rmfm7WsH7EIeki8GdaYk07R
wIfHwwEfuE+f+98qpkLebolHwClYsxfpT8BV346+hlyEpujVsOYSfCKjYkSvswlZ7CBvOK67Z9hC
/zhGPcaWxslyqJf7FklZ6aAEWH2jGlYRdLFW1AUIxLb+mTwVjH3tdWd/X7lpRAr+HFVXtWXdXa5f
g9HM02b5V6Ya6Bx131kUDVeRJU0eDjx+eYH7P4adYks9byZO/TuSSbbPYgqpfOLmbDGeu+pZgXX0
2OUzgpxyM5BwqiJqzI76URuHnN5i78O/eM34Vi0ywkr7/WlQe/nAFDEIxwO9MpcyGNxf8a/F8vxU
7QLljFQ6MIehx9aGF/R9e/u6U44G/UnCQlVd055gBwNiUbx63mdE960PA+MM9OiPJ9/EtMOZAptG
5Nf9jZNaBiynE+xYXGs3te3q4v5ixQa/IVA6Qpk+y+rbhR0mWYsgj6KCfNGvxVuMMXItei9mF2mz
08oIeQTgc1mR4UlRB0YftAzeuyC7/arX3iYlLajnQEtY9kr7j0h8+4pHJccs332oiuNgL7wUc11i
qHHd/kzDuVng4A9ID7kg+UqCBW/Dg91LUANbMQx9dAio94fPnjWYlycmo/aEleIDB3InKGE/lKD1
XXlbiNgidbUc4Rl1c2mg0JDR797x0sBGDINnAfCUBbTjM8SgsC4irY/m8qbJXcrZSg4I0B8msIUa
DEwyyO0rZMRBl9qU9MG+uwAHQ6sbbGHJuvTnNPd3OQkT+aRfv1tE0Ub9ZUt6ZXgqWJifCkhJpFu/
LLQ5nD9tVMjsiUmOQqIm9cD2n42xJ6ZHmMjqulPiehc70num2OBt9QOGLo9UxJn/YS3njvC0KixA
g6U3DyVB05fTK5OFVfaVKl0ZcOvf0sohX+3lvcz1WeBtnMu6+uJTvUdBapdAwb1/rSftiuPgBPTr
j85/v8sHJWKJfGDhGBRQYUWg9l1yBeDSGQRk4L10nfKKN/VPtm67R4wot4c+usTo+Pp4B/CcoiB6
+lgcy23/bDbOZJCIagxRIyNN9hU40wzQz5tZXMyKkp4VJDmDlOteKA526QyB7lm+C1C706i9Wfwb
GW0DZ2WDBZBLV7RwyZcnzlBioHTc7PMinAmmLZNLV52bJRHf9bnv4A0YdVmkLo7001RWpXVnhFIB
YdXQnuIE4Qo9nA4DiRVNHORO1kV17yeYPVlaFnbdSTEAPjO1Twv9oSgzbRCKCJKgOCdint6+wbqj
yH3Xlxj6y0ylvNIWDc8th8F0HZpJi2iG5T1vSoIsX0UiBF60Gu0tOrMAbDh0d7VadaCPMK6yEHqx
wbblCMtV5hlKc7DXKeBRcMlxtqRbCj8RBEjypIL1ROWIVI2sFzBc9Nq3r7JJ7teCOy+IxzD+kmZN
QgunUKs7NITGYGZGJsAqUMKBbzNbPy2jXLsYSEYCMMwIKTrN1+ANrxZ250Tn/IcwRGt2dvVqWbGU
oiaS7LdKNIoirHkGoVvnEzHfyt7tFYgV0cULv/N30+t5CMd9k9wxVS3I8Esv12WWUn+5C3raWWFH
dfb0Mgl+zfKVCl5x9aJ1XAuAA1byWuwjciORaLb+VngKIUBP5eBzVdh7eYRiPzZvi+t5o/L/ptvQ
TuWJ+RxJBD5Kyrf9iHWrRAlcj5IdlDaxC5ikCU5wbPeCZL7D2xbVtZ2q4dIeGMz8/Ge3pp8qQpNn
lFNmPb4shhX+08HQU5oYQ1NAqimI9rHsZlac0vEGPNT20hapRtiJQbfejsc8H6HZeiR7ubinrWsi
3VCYrWnU4DxHZc/OoMhTTKAJ1lCIRZPd8r8a/VdQ3maIVOXAMYQl0Ply+CFbW/mWVrHJE0V0McEs
4DVMjE+WukkJc72E0eD1XGrceuJTycjgwQ3SRMSSlQ8iT3S3LEK+8f8rmhvTxU0x47yOHTMD5pLb
zJuPPhTJ9jASackIVrndexdax7S2v+X+tEaXyRpxUrOhlcsLX5gs7I9Ugz4RwRqywCI22v8eMwxk
7pgS0dvWE/hR5qFlUC8+N3lY4pgCaI2NYZGgzAamvgOFxqNBjy6lzR+ccV5liyaNZF9hjkbbtLuM
ePxMpU1dKhdGavPxypITjw3EcH114bw0qZL+XkIKRL8t78WLUO07VPcGGvtwkOYmW6i9wOex481L
8M8NxoBSlkiUycSG3GQ8yLhbWdQ9NIpv2aUCurho+mlEvpbYcy6htwjwFnLr5ok7lfj+9Via69QS
uN9Ly4FYuLeadiEmn37YQpstQkdGNU813NinOdd6hGhjmmdO2qvpIEjxRt5Vyuwx1f4npUxdljoU
Xe+its+4Q3Wxm7SCJBKslxQbAwkqfoVAIksGWIV8G0czqEazUs1QbxgQ7bjSYQgolB+eyzA9ZqWn
v/NZdtGRqF+xE1AwtpaGd82wK4dU4P0v1sYaDA00XNNYXLfZb+KF/MrvdmR6tgPs1RI/e9p/5ylH
gIKvfIFUSRrhFYQIMlKY2Rn4OrY2620O1jaQ4VtlUlo+joSX62GS0q6H3BgUJP0oMFrMIngcIn+J
n5EoBDgwJll7eQC557Xm4ETpT86LfVPPTkAnHk5sDqXBhmLZ8oSaelCiHmhr+7IpWmJDM8V0NewB
Wmni3XDbipuVv0/CihHvRSoWzjoDpvCD8HOTnEq9EaZ0jBT/PGPAipZ/CRETs9CFd+0jUjd4GZ7W
TwKBRlXKxHnuwk9A8uXkw2JoGL73FLQy2UWZf/83jZPSH6brkW2mGSMQzIn/dniPcJfePG9MCQqy
tqaQDNIdjDIG1+70wn8hswpt5iNxtNwhl1ndyR0shgpJ/FhmkEpL7JtK3R23uh8Y/T/k5TXHXXSV
ASVraI2pn3sJvsMiHXbCJGBbpO/N/izsIWdT+VHt400CcX83+qpH4eGs7Lo9SvhxemBlsaNWFNpD
qcBeNBqan1D43qXDlYQqfgPGk/S+TIZOB1g6WNaZ5L5NbbB2xidioF+MerflG4WYC7y9oD74zkrO
Rbbli/Jc5Xpn45WBY0Z6QRLe5/DSjhFxmI1N9P7Gh+QmEatv1Zubms3/XVq219VEGYnLICYSh8f3
asJeQJClVqH1bbp2yxQRJjpyZY7MNCVRsR/CPXfPjlosp9YzZIBxgv/Zw9ZUgPTqT/elrHDEom+N
1eich49GjoJl9teTiMNIX1L3gwpeZC1fJBu9FaLQI2QFyJkja3J7+m1s5qnXc722EiuVz6FRM+5Y
ZVWhJJJ14mZhU+iqJ3g4LyuVfJVH76m9ZgxPFE2KlKYzVgg/wpQprViS6IGehFAhmmFlEsg97qd5
C/gWuRhg9LkOT7nxH+B+nf6FjVHF3MdfW+3JG7NhEzuoUlnrazhBU7eeUELaUw1O8Fk3YC18OS1+
1eFPNF2C7dPyNr2LfhW62yB+kURdrWVRIX3ofIIoRk0pnUtidRyRADC+vED1lODl21V08/gpihXf
hFpqb4+dP/DjDojGgex06p9tft2G5Ij5flh1UgS5FLTpZbJiRECq/DbTPe2qNa1/xeUAggM1A0Wt
pGjeqU8ExO6NWuh7HMd6MniW+HT8XJYkCKYr6x0Zt3XbxNKQ2G25nHWdxdy66ysZm3b0jqswgyIb
NjCXkl2I3TyywKwQTaCB8y3hHfgm6oqUk/s+Q7kF6tZkdpIiPDag4TKV98gj06vQA+G6QvO97DW5
W3UvUm4rSDEVRPpg6+iWCvaeSVF7ItDKIHTF1Lv5tAisu5hou3uS3+0R+mMvVLUye3pavtC/s3Y2
QzgmsWUXANXOd1dm4/qrpC7qC54LeQGSKw5rtY112T8spZtvHmJ+Xdig/y4KqD54ipYJCusfuMDF
JElgRzqFzhUMMdMYd6qSk/li2fpr2lCoaHOIVNu4STtds8ygKfTcqtArMjyvCBVcxY09JG6lXb/C
SfAxr+Q9EExoqoPPUETLivlLLamozSe6rV9AzDsJGw6uDtV0N4SxvX5UqVyRvqxOjLq3VYodHaYQ
ne8U2NPF/kzotdibHrwMGsyDg1NFUSkAr+VVGu2Fcnn8i3AngvnZcJ0Z3N+VaKAVMWCu0hxCQxva
WnOwj15qqfBnkjlqbXGYz8hpVHwSni592zljvnJuMJrhUTZZZ2+hBu4kUS7oVHtrsT9hu9z41XUD
pgTGfo30sWXgSW/zHG/RpLRZCLYGFsE48mCd6/at1OMGt4V4WZua/MQ2BksvmwDAURkKvhxF2XTI
Hpje+kGRWW1Hvgc6UQOzbnTieNA+7t6lKGT79R45E8rh0t2YCcX3a243vjci/bIhRe4stOLL1pTe
LtXliqEH3jJvhmxQC7AtkmXdot7gXmi6OAauVIVhb45z9E21J75eKUBBahlmnVR4NgErdiv1JQtB
q90RGBNHC0rq7fGiHM5uq6z5wpkcKzsbtKMsWv0COj3fBbGSsrqFAEyUEBXxGOEmyrFl/KMenzVv
pIkAeX/Ms0XEjllooaBYgZCgxLuQ8dnZSpTX7pN1FDwEmQEiPWs7pkDvCDpwzAlQE+jNCDIeCa1G
KD3IvnV1/6vr7315Rm/nR7mAsRsTURUQYkfQEdZwvNTOCHUIhWq7VlTgsKkk0s9GiNadFX8+ENSz
9xkNEUwBBL37Wm7opsA0kHLgE2Y5ZUQjDGUKDhhev8hyAmRidEccTl+fVf771xMEJ0LSNt7nvNjV
2RcmoVSncJbvvNTfracRGy844iXu86btAPKTT2xtKhQoJCWHi8jmofUGSjdDuAuo8F9r/jAJQlU6
lqkxmlHvLsScwJjP7869BrEU5aTMiqshsadMkfvp69xgs9ybDZU2hznFwc2u/a88vJzKX2/MdHtF
vZ+j9saxdHQRmi1unfM4eEb/LNeonPg5kVitU96S6YZqOhUgSgCeyJsN54ihdtleK99VrfY7lFvG
PqGvyEI8wITny1n1hDW/aie2J9TNulZF0Tm4p+jr0+EXEesO8ekJCrRRQnOjuAamvUa6CA9elBBk
h7Fo+LXDhAHw1IAoJgBYQNqvy6sTp36C0oaY283vBz3xxrc4adCD5RGtSAruAyChvfDfdcu6Rbqj
fexAGV1FkqxSpSxvstneLUF4MGl6yGaBo11OecfMTwSIVe+mkNBY28ElNONZhpgdXgo8N23m+rdW
yxq+gkesuVJdGZ1OW2lpruEaBR3Pk95HF9Gk/dYZBKeKQWAjUQsmWTX4GVQLb/luMLms1KIjcY8T
tTPY77P+PVWSg6yscMP8wi7UQ/bAetLoZL4bqjLgdGQaMtzlVFRqvdhVvhZbt/pYkNw3o5fdxTjj
gpzRhosXfZ1G7meZS4OZq1+H24qre1MrZ45NWpKSIvD7c/+vivjU5wDvE0tI38weMsnBK9vGWLFl
lnnyDn7LhR8blgR8R9z6STRc4DA2zkO57oHCfsUKEd7YKU1iLGLLUr+R4Yj/F25Fnkr6MUgmF7Uz
BpindpxetaUvJ1Q+U9DGN0m7Tn+BHwuPi9lK0MeoTUKYFTD73wrQ63hNK9y6S2jjnT62GD792rL4
rSkQ2kUpdTW7LyxnFsjcGJ/y1/Io/Ezqpie5v3GO8xcMmmUjnOraQmwLNrsgXKxzr5xcy15kEFNF
9bq20yISZPRAZ6xI8twXFd3Z5fo6DkJLrYtTBu2F2ZjgRNUyCzoYVbPzeF69MnrPQYgB+Nke52fF
QI86kCcZwFRfmXNac6Iy6rMEWZUBXKiXBjv2Sk1UiPBpiiq2BrVTLZY9AWTax3LsJqpRNsYrAGA1
hSHizAlHGLk9pyWYjVCmna3WVJol4tO4NKS4eE+V2QWC5rkFhEaBmRUdfQDf3f2eFiIxzSbvAwBX
ugIU5LchXLwwx/lfGQ+HEUxNesUSHfbePECBtTOgkZrBoCehLUNGmV15hC7lUWrPjIoOlm0Y1YJ7
AvoHcmnp310gWl7pBrLn16qrLafZ3hPJSr5/AIuP/e1jsRB1O6RGEGW/ZVmsV45FUCpz7Fa62RRe
QVU0mSAan1y29UfMwCDXpo+HzmE3I7/1/RnwvChaN9ATn4dmCN7GJ8pl+nIDaT2CR7w6Cjvzm1oS
R5A818moMBnocplaVbyeODq2WtHJGIiPFIWoxJzqVNopHHUeRJX+5OlpAELw7iC2Phjg24SriY3b
6IdpyNplux5mW5cr/fJRkXoq3vinUO1mSUR+cAvH436ZAsGB/ID6SloMkYIv1K2y+tR0CTplgwGq
ivQAhSMSlIPZ6V7s8soel0dUmG9XHkHUozhLKWP4BJGlV2t/CRch3VRMXtzVGjFkRIp3qexxLUGN
vijuPBi3EfZeacRgn4hpxBtl9VG7kLFnhUseJBkjE5z7oVPfVYxwLI2HYeJmYd3bQAXoUnO7d3m2
8pVwHTaqYwwWcAVNZkZ6KstiUWPEadqcmow7PB66XOtAfAJTSzSNHw6HjeGoC//OK7oM96tiBXK1
RjsxC7e0aW8oADFCbc3vAarRGxhgZKJtacrP/0Dnlw6COL2NJ592bWsHQeeF/L/qLC32Rkj4Xur2
YFXDvQaUKop5+0Nyc6iBjMWegjYWJJl5LK/dgw/fJ0KnYrUDXk/mrIctzhiCtgUrdJ6SIbU/QOMM
bFUQdEhjHXkQDyHGBzPx0kIpmINDaHa2pRAPb/0M0hlU8Wxv46qR0WjbGTGMdxNdnRlRsbVsVkMV
58aTra4sFiIzlrKcte88ha+LXdb1UvgnQVHi5moae8WrSLXw/+R5XZmEUOaNq6bckHpzjOAecg0S
J1gzOwHBQ+dlvK64KmQxl/KaPyj0bOpGrR2DeB4jdEKpRMAOiTk+QcRRuEv1tz0hH0AqFkGfQh6f
e3qhTNKHsyhIzoLHeKn0/cfXIdJi81OxKL3qJqCaGGLBkyQIfF5gVeTrEu2jsHPtt+sx6f2m3wAL
VFut9XOjDDSfpn7zJOLbV8rc3UHTIqW50gnH7/Vh5SZbhWlgkoU+aXRc3Sb2pPxUBBp+qtTqqwmZ
SohuHBquoVH/J5yw+M8nHVrm5cZZ/JOmDo0Yw1sX3xZ65f3VzzH78+/lJKLndBW7E1smVxyr0j5t
gFD8EApqsu9YzgMWBQOluAw3uRpgzqtQ+EmDET9nwL106CzEGaPr2DJmc9OVCUpAXGjgIGPNayya
hoVhzShmmF89plsjymmpf6bz1x5ogWdxYv+pKAsyDoYpOozqgiIoRe8fvUmW2AJuvtLMJjRL5hq3
1Iw7mftowaQYnPwZ2zZPfKDxH9uaXqUWGPMxRx11ufl1ntIJnOY2sAZ5A57JW0+clh5xBX1AYdid
2XgUSJhmybz7zaYs3E/OMGTDrEQdnYW7pMgT/yn14fvy+tKaC8lJd2WDVoSKKzRdJYZpKQOCcoEH
MgsdekI/nnfVBAyI+2+5ONi7Nd0M1jBVUbcfc4x26RhARhBAuLKK+UaJ8RjOwCxA3KHrfbZTaHMm
Bm2giWNUKfK+cEmfTF6r8kFTlTYcsMIhqgNA37zcjiWWYTx8Jq5K94JdNEfInlVTT/uXbDx6ffOa
Y88c7wP2HRNTEGFZTZBhqMZq9r8/kHbKmX5F0RZCom0cvT6hRngrUHCQ9H4wVFtFSB5jNoOdFqBy
vUoPsYXNYn+g5XvdQqkFdH50S35a5Toty1j3985eOseZYFLlWHfi10UbC7dkcYezT06UZ6HfTE9k
MA8aIsoU5ivgsoBTrm42W2qpgGq+dg7M53r1uWLGmI750fktyX3OcuHUhNhJOO+Zlym/z8vsJk3V
dwof3aj0Tgw9PlwUO84mS4gq0t+2FOJNcqtpyJhy1ZLO94qNpQIC7sxMF7yF2NcLzjrb6Beayjx3
tUD2HSumP80MYSTvoiN4XGxP1v+fiRbWibUqARpD7q5a0R26YoYc2P56fvPsmApraWgq9L47tfpL
zzjgsBrkAntx4RSMZeNiI78JukTfxvhHNpvUEy2JLxttSERsg4loqNQbLGtr2V6RMjZQxK0xUnB3
fJ2C41Eg1mEYoHe5WtIgp8MHBzy/z8nSZ+GbNA8sAM1MKrGM/UozepZ8YtS2VHLSfBft2gPAchUZ
u6eQ7l/6U8LMQqVDynfY0xN7K7n0w2G+RVAQyrLOq9nvV3r76GoOg92sxmXL3ScZd6k6P2k4DpNr
kXMOWsgev2xkOWFHe0X/Ezi4SiqmJtCuya3LwcWyl6QbFQC6sNlksoaqxq8JKjamgmTF+vCujMjQ
jPkeXVQ8IW92KxwVlqEiN5sqDaIEYoFpAg0IAJkUmYEeswcRLX1wL4pt9HZsibzeNGFOXE1tzxqP
l6G5b2MLB4QAB8pZmbf2Bx+71jmsuRLBN5AWAEN0NPTj7fbmhBB/wccqun+xlIMlC8lATjDVdwR7
2nhKZiOtvaTQ23g6x2FLAT5ojFCFgJUQsQOx7LjYYoFcFeFphZ7LDduS/5A5xs2lxozBysuQ4FkD
1Yqf8vpo5wYDkDfNURPKb4uZB7FCldVramEdzG/cDsluPYzRrPEwKyPROItv5zfMsiEH3FJJL8fG
a6Z23ZNLanCa3o+58wWGlcyeptEvKmZ4g0L2yOfHpLw7fPWu+Pkk809pLsfCHA4A1cWQOunnQmV7
5SX08lR8pxLeycnFT0ygEFrrrYwdTFd20N0y/Psd5cW7mC5KLemKTwk3wjzHz4vYObkL3dqbVOfD
+OpoS/WofwQ9/D45/MIlkXEoYW5qRbtEdL30C0+zBS9IotdBxNjvYokSRxI7/S1VvCchSVyZoFjs
3rCsK1SzER/Yj/Y8qTv6oEN3mMkfyeDh43tylBzwhjQr1UQmeBVMT5VAJv+uEGRae7LfQsHXfyqG
rlIkso6lRsmeLFErmiB+TbN6cNCeK+nTSFf62XEMn6B+3mKsigWTMsgiXfhqRaOv0MCQSwKGn6Ri
Ck51BwqwWKKrC1qGG4nGdZxBeey/8ChamaFAdjiyeav+FoDcRXPRp438avXJTnHV9jGr9hlfck04
ZTagM0uBV824ZEpfw0uCal3I1X9ocdQfveZRIr6vCofpWXYHa9019xyqsI1XcmC1F5/xMxA4Hybw
XJ8xG4NRnU9reCm1ZHGcIofgm+QFq8qhtmaghxFm3H3f7tHYePBZqbc5yp1359s6Um2f7oWmS0db
Ifw37xK3vfaw33fHgYKCju1y9AerI8PZNcSxRdrOHYAxfJyRMztR2gBl31cIK1spMM7yDc3VD4MJ
hrXP2v437Xfs1J1MkG6tpqZD03D04Bt+NK1jfXlg3AM95TF9PTq2A6slWzwCv0hBqGArGht51LDU
xFR3pbgPlTgu6HgMS357na45XtZZ7kNge6H+TrIEFwlASfLZy79ntClWt/DSmoLu2ilwgbqbuZNI
Ekr5GrfDqm3XKtfipprT9N1bGJPZxu2FHqg9CTRdUwAG/UUXIIbVGmcR0QY3nnfB6p9nmC77I4+N
ZuTFmdpnBwM2WwzfAoFF8HqLNJZWTltm83Z6C+dJ67oQ4cl1iNP0eyuY2rZHi+AK36LD7/jjxFMc
6AVd7cXoM/i8/bugYFg8+J83VdvJb+lCuQ35eogFjy/5iuk6sU/aZjvrdvFFaUtXd5VmQcXjMFjG
VdoIrft9Xfm2BkgD/96FueyaDyChlIk+auOubflO1rnkOupV/V3IE0u/qD4k2Sq52Qr2QIMagRXs
zqJsfZLsQMpGyqpDVLS0FvMEPF15RCKuNM3EBiDtPuf3qzLn5i161jLuF8ErgK/Jgih+TyhDidkD
V43UEj/ItB9lU2SB/Ujn/OEV/EF69cxEe4QFp+Au81/rYpMsTqNncN0NLJnsaTJTPvpcu0Vm01V+
LcJupzq+8MBlWl9VI5i/fmLxijfu2gIASfKuwrV3cWJVJCISO49pYHNAwHGVzBKj6R8ZVtN8JvYR
lyrBZTxxfAsRfuHej0Ta2T43ZVE5Amw0joclvaUq1bjkV0JmaGo58Fx4NSxIjwsXwN8WyGkW6Ts3
g8npmG8JOh4VtsLr0c8JB2L+30i6g+kEukZcURA1fq3Boux+7a74zJGarmJ7BJ4exGdWCcvDNU+5
uoit0uXQQhebZOZ8JygiyCT8TINf6LQT//xotAX/dekfU4AOwmKoCifZ7m4bLWPKOuHdveAS4rrM
sBVFuN20yQzliIPtvmSsrhxPhUSYyTlkKJvTvGb4UXV21xDzqga+TzjY8vdCtOh610BIWXZqbKKR
oS9TmZQKX+7T7XBSVRXafjk+SW9K18zbpT5ul4YG3VCsFnfMhIEzmCRLmhJghCW/GII7ya133loc
czXbig+dnpBr1ZXguMYe3t2KyCYhlCOcUDZD3euXgg4EYnlMpQhFvI4sw3Xjcz3TrPObomBpfVhm
IipsZ5X3Yc2fTZtCJllI0opy2yW9m/KJsGqULslklR+ApdI4uWeuRHtqu1pQkfDtN9Dtt5qKIXuV
JNega7QZLuClBmYwie1hA0evYNzuup6GHJiDSq3SvOP7/v3Ol8U5X/hamBQzEpO2UvWmpqgvReKr
BaBE3u5lgcxftgz491qFgWnClfQxy6yj0Hn/6mle2WuwJZKqSu89Zf4KF3oOBoTiqAoqrW+sX4Hu
vjN4PL88z9A6BmwUbKJgYCJ2S2mE89m0TDhV53pDP50cz6CD/NMYQ8CXbYBajOCem+xg7bKoPp57
y6z9hmBhtRGjK6Ac4Yvm+2c9nNJ4cGLKFr0bRsyzHWqmZKaaHt6yTAOaZOxdRRJRpafNliEFZovm
UVPTT41mgX6+mue0LiMXYAln9HaU89hBRubcSj0sYLAdDjVxQQ2HgZcS/nb7AjDanYX4Q3GpbJgl
i1RSklC/0WUcWZenEu2Mr5v0laZrEQcZok0KOc2J+DLjsMoouCrJJ0hJHlEo541UfHILUNgqClLj
TN4+JANGyX0YKtAV4JO2vFn/F9TzjFJC6sWIUUAUNKMi3aMTwSy66lLbE+WcvmJqps4VNMLDPioi
yZvrHnuu6oM0dUKqfZ+oe1rnEL8ecDZkXRpWSBkIFmk/M21TDOeRfojXRbetEW18xj9mA03ar36s
SO+YjkjFIG1PcBqbUhL70U1gfPS5yZ1Y7Z+rFtZxCXVTXJx5OGmG6tAtDkkDu07xbVe3sOSEsVmt
yqhODGxQA0iy+WBQcZfsvkPkFvj6mzqSr4iSyNevtO2eaH8uBxOmhwYHXPEKmYqQKzRnmeT0RpcS
XR5+8mr7Za24loZoQmNaPjQksoeJC2ZJR/GuBDrwOvVvosu3/fbkIDx1XEMQXVAH3noyA9jj/e98
1H+EWEqs20zBts3MJHFT4ROWfBKewtNfGgzDLNGKB7azQ7gbWhgM1zD5XKAjXdAmUT5Ne5+X9eTg
nruXY53hVmRuXDpGToH7X2zl5mhGkbHTUarKklsXne1wH9CtspTVVoxa2ceNYT4BZ4aYqQorAaqM
aDlbt1L9hvv6rIQ9pcSNcqoi8guea5k7g5MM1MqYfo7PP7v4cmN8Pg2A88dnxbPJVrJpTloeiBj9
iuo0lhO2/EQY57zMFe/j0il0juc1dhvLqPu0qhAYPV2Y5YLuLE0Mm21uxoNdOdWzzHCQMDawTLy9
aqG7HNuw0o/dsjkRMiuGDBGmpNCjt+EYqhYVZvk3aucCjNmbPJoeFnJTtq0YFr23UHwsXyTeWkU8
DtWVO49AN4U/VFx3imKZfh/Zlpp9LFv3bR6rmMcLVHX5o9Tx+FF2EFex/yrRWfUmYcJSs/4wijss
Rr4Y7+lAISH2sg2ma2rr5hZsdl7d1OLfGwO41nZxlb/6eTMKbrckU2l8peYtfOn0uzCUvxnvceQe
KmQaUecUUqdMh6UcfWTKn/JgNlsjO0hWRMTxZnKtP+KQCOYIWLWx5glUN14gq0wq27AxTBdONtBX
tvYDano3G8vh8WJqvGnJzUPfmWfYT9NCdwWeKdCJDjykq5Lz1D68OPh0yKJ97y9bMrCnuf5ObiKn
VhY7knFSdB4YOxX0Z3xSJ779bboDVLorQ0ajn/xAQQBYMXnwxtiKgDaYag/6QYVLp+zYxPDmsJQJ
uQQlk2RBgVUI3+s8+UHh4DxSosxJklZRL9wyh4cIRGhKIu3WlBygNtuInFc3EAQ54SuFIhdwrfr7
zQ1bZOrdjxpTvDKlHppHg1qwNbLZisF89CbVJdTh6jLhF5WxU1+agsWUuiLuN2D8e6RnW7KJ0kCa
1Ant6z+CLhbOgrHGh3vYkkcyF9OGHexO3VMRexhMsvG26lciQHb1L0mkujZtqz+arOjHTLrDtgkV
ItMDp2qTac4gI36DUXC7gTYbPP6UBPm+PsH6d+TKMFDoe0FeqStl/vOl3QKtmfM5Gc1V8lDkUUBf
rDzD5NJBUyjABWW92qDw7KV5RBWdlX4W0wmAtckD4niJrFjKRxjShja8lYPtDfSTS9n1DJlMcaPG
tftu/I5atyanlvbjeBqppq0F3uOxpqEizcwcmFZWpESLDEgCgf0hRV1519oZrTc7FEqwTiEa1kb2
9RQR+aPb+Ev9Ug/WPwjv0ghwAaPi3XDHapzF7XFqXrPjKeY9IfkGdEDzO78/+laBAMjL7DAgBB4l
b8CC1WrrA6Q1InlcBwtIJ950JgUSruBhUhiSAK3OV4DmpXtMRZWdoRyqPbqPwEAwz9xV9n1ZBGRF
FM5EemsSgP6aZetOPloiy0J/m+0n0I/iupL6Uz/CLp6F+LbEzwA7EqVvXiytDzWRc64exPbiIu4d
ah5lSXt8nO65yYrD0pIrb+e0SRjdraAu+Q8U1MQcwmdnd6pdFYrq3qyAOEewRup2fXwu5WZ98Z5Y
Vmkx3arxa8LgnI7+NGppIIEznzTWdimt4gqdf4mPu/79MaCSQvMR9t9XkpMzMhGe7+Gz7cjDFhJ7
614RaPdSiL2UuFd6NnLH14baaRpRwW6xBEmd4QpcU56ITvEiFuH6lHxol1swBN2BiAw7sSnJXJFV
x9qJK1tWR4HL1TzU1+Ik64/xBAJ/PK92F3umWf6Vfw1qLj+F4gGMGRo941WADkjF4N9uSrSqG2Zd
22QXh/aNJxXPBsMrYDQhrrG5F9u4X/zcf+oVjVOym0cjFXx134mSDTFEIBkTpuQE5H3FMygduruP
xyP53CdfE29wyCL93fb0uWurLCeIBjiWA0Ak0I5I2dm60rdlF7p24LnfjlUzejvJAym8SUuZH0tn
6+r8tYQBFpBjVzsP4p+8Nfj57AjPf8Y314Nv7H2TOPtiR93Hh+0HQ3dAOS9sXmXI3rd86Zw++ot5
a2QWV/HuYKf0Ma8GfBTQcewk6YsqpGHK6i7fQMWVMkZFUH8I3nDReJZZUJeURBpYeeIv/vmKhZbG
yR15CHAqFvM9lk4NGMHBYR0rKfe/9FomsZkgKOfXh7N//U7IYWpUO6rwLuWGJtwlokAKaKxN/Y/A
0G2zPufo10danCk2raD9Z9nkuBY7J0K/lD+YHNiqsR/whlCWIfUu1UvD8g8tYVMzjYfJd+86008B
FxWmGXMCFvDjzk+h9abPKhr+j8QQsDLl4+UPB/5pUVJkYwC39kLoZUir+1oJyF78gSSSwDcwXKtw
c8LlSKzji/MNzXwr9Txpusyr/Qai7kaAF5d0r5Mdp6j7EzWLjeFnjYu755rntf95O0j8OeVxiYaL
/YszXA9PiHxx46WT1g1dc12HB5Q10j7v0cPbI2zaTtfSCjJxvbAXuYMnF3aWS/Of2/pJosUbceV3
4d8JbZYHj4gbjzVb6j2CP5FhAZTXQ9XpafC2Jeicrcay6kiCw8hE9NMHv9Kkp3014AqcePKSvUjj
We7MO/Yw59gIvFeUWG34HRqhlDZMqkuHG5VqhyL5YobdB1ttGaEJiupCsdT0HdXb9zKWiV3Pem7r
aIamPR//oVb1jDMCaNQsDRuOIbjB/RXt2oX771z9p99Blz5q613oJ4aVhnGBiy+xnvhqeBHtWMug
/1lIXsnisQLiRqGnXOE21+LM2DP08LKFU5n9r+rRzI26wgm2hZzrUUMjV7gu2MNQ57gPpbYELfi4
ISPIMaPmlwlhrV8ccsVI89vZhH9NFMySY0qZNwgqm8wsBKYv2aWKl5H4wPFovHjfemmhq1uzTVjp
yJ/DgR035f1jfxnhlTpXAOMMbzql8b2izAJz9ne1Tzahj8CZhFFlgYVen8i2IfNX062ZO8dmWVU5
XyySrlbH1U6dOSIIWXP95u4OA2Yl+kKN99gdQuPWMfC6u42+gd4/7zFL++fMdK4oDDQgQ/poLqCv
gQF8IWem2zz2uOV0bQjQrvR0eQYvfFNPf/U7lNSbhmpM5+m2BfAMCq9bfvdMsRkkPZD2QwcJowOW
RiPQdvtr4MwZMe0y1UKVpFuSGoZbrrg8el0sLODgQp3JfBttwPHHFBAFipqT6yHeSJZTWcw2gi1D
J25P8cSYjYLpS5k+H83Ya9KuLTaJCHWNmcK6ruBGe2K0yEnVEEOEX3rDXoOdkrH5znWUkrz3UpMt
mdB1cHSIHOFP//GEIl3VBtqZX205wfRObDUu8ydLx2LicKJC1OACBmGwG0nHI1NRzXkrDfoIUMd2
57mnjGZN2dceg5rQdfj9x4XENs7ppGR6q/BYnMH9NZ875oJ2EfawttdOFI0U1Ty+0VneVIc1oRYM
f+QePd2Z3jzb+/uNOwDPqQmiUQQYneV9fFPrGu3grRd6CXmimYfRMhX6kqkJLAbeYd4gVyCrcx3J
LJxPikPdz0sUiFKBggy1NdiCYInZFnUKMM53p+IO/XJzBBwzl/eOaaXvWu63iXR0OjtRKE69+l59
+oYJmnOgpwigm5115b9HedByNHC4FrB0iN3S4YIi+07ccUMFMLmMnNvTlDLR0EG+cKfIBLUKj+ne
gBJC7sgRaIupnhMtNOwOUoX2Nhj7Lkz3sP4RfIQt6jJ1TPmNr0WTcGTsYpKxcB0x0RcMaf5TTF3T
OZlpJLHp5CF9MQsKU4bryqOU9PGrbzwtwbXCH4L5+AHXA12DUGMK16va7cu21IiQLd6tPcD/WTzF
4VXuPrAfwN3dbKUiuxPNCDuQs5wcjVkH36rJ6mx291nnCtwEFPoZmgp0NZEeU0uDwJDNUehdMxhw
h7Ys8lbEn7fRPGVriwXIKEFMzh2j5hR7Ou0RQOO9Gbj/PWPQIe4v6iUGME1ESS6US7UJHzp0sOn3
TgMjhg/mblGFLQWFmMQfalLFiz4iVnPrdxipPW3IE1CVG3ShNLlWvmSKGXyYy78FbncBAebKTLXO
k/X493F05Gyn9/OITxBvY/Q6cRZCcqQ5390QlIuReCZiPh9VTmej0/wPC6otOy/jpMtwoTABBMGP
7uh68lU7CXwIs/oUKXylDaml10u86BbEhpFQxVYRzfdSiVpj9wopUS0AsbZnG4WXSMPFI3LyFmHZ
1CrER2HFU62eWxm+r1FoO5AgU0r7mvGUl87XFUDzadMthwdCaZQD+sK1vCjolZMtZHqjvQHFHczu
nHsEaE+Aa+AS9RjiYhjqKImZMxX+5HEwQBzf7PK3zxilYuiC6ENeF7xtmj/UY6oyTFYJPzRaT6C2
FCVeGlP4M6WN97GNdTUbXVKLP4mB4aOQai/fmgLsNC+j92kuWmdQN/rrQECd6DAOLXSvPXXmrZZm
wSzhHC7hFAP8FwYhzcmVUcIdRZokt75Q2t/9qZOzYZBu7spUQZnTcgUJrf0nx27YY8rysPo0Yq0D
oG+jMvu4Ic4pRHtTF0jvdxkAwJm9B/uSJHL6oVOIuNHIKwKrmnpMd5RZ6QifW8iruYjblBXqSP76
6AfwYypK5CAD04WAUvgKmHS9bI7siMVHZEjosCqc2PP30bF0V6AQjYXP9+kTYd49wd17sUzKTv/W
QmzK71vY2QU9xsJepGQd8wyHSgKdcHz89WSN7hdbuazkSHISelng0FNxhTOPAjpvxP2rc//NPJWW
iVFdNRudHpces7BW7I7tEISYo9lYWvXKo/r0sHKCDN8edABRq9SRKx03Qj3OJOfSJ2fR7H1IO6gK
K+rVnnNOHIr52G8FhhCUtJI4dXBxwy3gbiRj9ovHYwNbxePVSyh3rIAJupQ17WK1ZGAegLHdFoCh
Ic7/XNI2tbghgWpGd6AqxMTme8wxwV9u075fjKRuUY4qIsIKFh8NFilTZ6tHoOEUa38hwQXDyo32
5hqQ8jRIuJNHbgHVvvXLmU3d8bXP/vTL/m/ssvuBIafzcgWfUa97LteQheP1kU8p/gG6+rcZhbpr
b/sUoDO13kL1y6sJgXv7HHCMdLvq2551UfbzQKlXjuXGMNMQu4saCeWAxenp13GDsINh9YtCJ4zB
1b1iyIDDIYpnIaMkH0suXe/Y+KGJFCf6RNiXbZiU7Mc8nrEH9BlRXPIogxzxhQvUauI/mjmMk8KS
iBD0sffL1Gx6uYSDhEoNSj2234Pi2dZTZcFn9j2aPeDiHgRwwJywinq3BDlvGRS3l9Wwzu7QDyCH
jg2I6t/GHVkHUrJOaV+wxBl/Wccgc/2DR4MSXzgKM99d+oGIzJi/K9e7Hm5rK13QtE16Vkd+xHzR
isaievhPTrE6yRoHAHZMlktP+fUZDRmT0BzUrCxCFX+10YPcqqoGB/8fn7xOHjAGoMxsN7w4OPb9
5diRIK3+N7UHOxAiIUV7woiwSXJuTgSEfJwFi74DfMVHby8+NP7I6zyGIRwcXEmoyW/nzMZsa+1M
WZzLCfsaZWKkuYFE7V8yyocKovNylIKT4wNw2vktxh4FnL1AdjMa2MZiA8G69vK3WdFm7ripTabG
lc7ByMCbtck8mNyLH84fPcB6L5DoDSbIg7MZp8057mBmTxkhnhdBR8x2VZm1m1XIUfCoYpa8tL//
Hc366+8nxClOXkSAWlpZmwG4Vo3TQlExRHICLcYPzSDJ/a7945iMgvqqIRI3/W+LXwafT6NBuvAY
eFRqEVcVQy9nTLLVCJfI8k5QzIQakbtAkOu7wMCYJSvdK47nynkK/iDG6mtjN4RTVDJWTDcfShSZ
rii5mhAbq/syRINvdL1W0bUgdQ/LYw4CeO1Qy+qNj8u+nWdUZ3yBPpz9SH7HTcYexl8iZfAPrpYk
Ub4WNtngrH+fuKnpL8F+SoOnyCn6EN1hccq3DfOl4rqYoC2u16gpYno2LYJY64BoL3iDFCGP4mF1
S89uT/HyOyFCGwL2+MJLLYYlDC0Sy7S02Y7x+9/MV8VgzLIgL5e6pge7zh7VWw2Ebew8CBGNI3Vq
wac0bCWGlPWv7Sdjji7qlb+CVqujJ+lLb/K+ILzz7IP2rIiQrNR994SviV/03u+JFsUeHqJNY4SS
0svmHKaJJPmkftMQ7pmMyJT5CR5KXetw73f0pnhxwoXBzqqXX8snyAOUDVvyz1irVrpLoXVULly+
UJjG2wijzd24cLf0+T1wxlEEWJNa8kAh0ajZ/6a6r7GF0zDMG61vTNOZnULhiVCv2Bprjt/trwoL
8Pj9SNaJ4WerjCVYklMB7kR8JxpWgoSQmu0EgszB+BuHckEuU877qpXEH0tojlV7pgDVU/vvtZZu
vdcVYMicq9U4Gsi0vZQZAhm/nnbe5oCJLLOLKOsXmBEByWNVpRgyY1l3t+ekhG81KVtMt+jL7U+h
/FeV2gUIwN7F0lXnAPZ+/mJiuNd7PEbE0UHpt6EyrpA0WSjRm6jj4WvPA99qWMgMbuJTAZ41p9WK
zrqifiufj9wWTDoBPEZWH4C9B4BrMS0qBWwu+0UDhFGJGGiZRsz1UqNoNvs2K4PANDJgYyKRshAC
HUyFcz29RH9dv1KEqh14oKRr+U77YH0sJBX8JTs8kerKpBk4D3hQ7UGaas4qF/yibGX8YFGt6sqa
PU0ddoz/07rcPnaT+VR8Cvcvi9BH1Jj2lCApNPWRTTl1k1D2HgRpbktzCsSDYV3lG3HODIdFaYFF
GHSmqvDIacL4IXuTkznJ7eUcbS2c+UKVsAvzmRiKRv1Zb2ZomJSetj+o8xjMIzuhJVS1TXDbRARJ
LW0fL84Uivoe/7x+Bs13geOX+FDUvJ80bOhXqxwJF4nkUKix1xaPbPBvDaulxeUkKg1QM6kVurgz
akDaUj3Vpqfl65AEEeE5b0Bgdogd/wG7YyC3wDJ0AQI5KWdUoxU40302MWQLoxJxvDw5EXQabf2u
EfAAEbE9K0eHL0qT9xlALzVOaZWDQPfmX1MIuJ49pw9WTjcqNUfAsG4T1+eOa/gr0dI3yKLB14sM
0sCMQI6yvJYpieZU71iY1sUw3PBgmtO9gXkf/YXvR3uhRx84aPM27LiYqgJAosQf0Exey6GUmOm4
TkNoSZCC99VM2nAq8pfhobmaruzsXyRzulfwWy4+9u7qF2jNMQSKnVo5fNJC2Gg5HvGA/1kdOAAx
+f1KLrf7rHvWde+0YoJmMI6e+pmpxwvacI2OwRxOEq5zwo9J/PITPsVKl0zojj3iiK6XW0pxn4PO
hF4Uw0mndnve9Y6uO3fjM+ZqbpNW3dzI6L70h6V6qlj0Lk6qKKhsCOiiOXVRj8p+/ORfrAiThVjz
3FWnRbV5lwUdPDgWRNCHPP1BRtfs3Y3QnEaqPqSsp4+y6kgzVxhZpQFY3+Zlfxq5u21XgeWuVUqf
T61AmWMzGBcmv817chQjoiRsaDB/HuRSi5m6DRnaJIWr2f3YoDblIvY3sDwa359ApAajnEnhWh9+
zzuW2dBMavtFoaiU2ut7oXh/XbZ2UZ7AOGpFZ+xGK/xlefbp/oLr8Ug6u9cPOIBEjE7kOskSl49u
ZUrEs8WX0OSgOwkzfDHkXhkAOQGVq3XEwFfWTj4H+Pnqprs7rIp0xDzPYASiFYCbiRnU28e4/Roo
7svH+HJCxKv1Kr9PO7dzGH9cyf5RmcfP+iRt7QsFw2o1OwlP+I04wQVPAbhO6/sdOLIy/ba2Nhe0
KFij5aWCpLJjXyQAzb5fE3WN4UW8lcZRlZMNatcyPbb6MkTb1FAINCMZwspxoK1YEKrwbkxao9/8
P1PQ7Fwb0yCdVfiZYXc3FCcDJZ7RrPSwUBJZFGLVwHhJ7KDwU9Mk35nkBwWg6PF2lOI4fdAeUoj2
kruEm/cH94ZX+NM+uK77C49MGAYb3NuGTqEPPln7q5IwGFTAQHkay9tpNlC1jc9EVns5GwEz85so
RnzI4n04sxbTb8sMaRd0UJivIhg4EwSS5SsZwRU30pKIvlGGli9SFnOkeuhzVMrEjEiElmJhgPIl
qAmIb5Z5KLqqakOmUYWA+4iv/8QCe6sMc2Xl+JWPmlaV1Ep7+kv/eJ1NIjHz/lgGitfICNg+xQq7
CFrNrVBuLT4C+bDAW8UWS1yKpbm5o/grkqpEYLhKQV564QyvLB4ME/eybr0yPOOCkRqARsc9MQnn
crN8psl9RHXUInUV1gP8arBrDrOBkpEU8ZM66W8gYoyOW+H/y5JYdMhuJE0yC9pwEiqewcqTDJPX
lLbMOWRiT9O97KrC1H2Suq/NIHVdtZ1v59sKHwvnqrqklKZYDiN4VIOCoPAu++kow/YH068s60AR
YTDSZJBWwJRBCjoK3eBN2jBwamRYq74quS356XMR7/ryBFKFhj88Jfkh7YECz7FEsbNx7dDvaU/y
ecklkYAggH2ygK4Uubusa5Po6lv/zW2yATggCcV8I8iCndokDtPFnOWVmuAQvle/j2LNDiWIDi/o
7ScXMwxCW+YNiw2fqjZgTf8V3xagMfQjTOPGMcKGzNIOT9ZEcrZmfI6Ga+x+cD10j1EjIjcXtPlj
Mt6+95tfeno5xzm3qNmLlQjz7z3N3G2tw+NbKEDFxHdp1uFi1cwOS75jQWqAmE2N3/mb17AU5KaZ
Zq+pRivfvMEOBMOzQJ5KU5XLBloUR1p737tohE24i6D0sTS62EKcG4Fa+dRitodOAo4MKDCa/Kvr
VWkX2XL2nQGX7XUf+tzlGid+vzO9KhV6ML1uuKo5RO+CeLt3mwZc8WsBacm2UtPIwem402EoVIbz
fbq13i5bP//duvP8BEEQDboPKRm35ksEXYB5KxiQT1E5EMHW/bFXRMV1LUqBDomKoHFG7qtRh4xR
wVQnkDX6Au0YPAxkrmtM2uky+6ocvG0xkj4nsDsyX29MNyyEGDVRUnTZTHjMpcunHc2IA/4fpnIn
rGLIvXmquk4PpFtSnSoCed2MfuQLspjkl9anZCKOMu7oMC+msAEj+3Sug7TRq2eECO7/NfDzlMah
nEaFiriUG8khnw5fSixzQeZorG2oiyBNeyZAu0aaZwDIz5mr72gV/IwUeYKdA1GtXbrd3z2N3Wkz
2edUdTCWT4qQI9VcV6qZOsG6FdVpPFzMzgqF/jUf10iJr+394PY/y/zJgraNZCR0p9Q706pQKb1g
wtBQ5MeAoQ8AAPzI/qk1uBSFB3tNkY3XJ54GaXsNGePiGW0urZyLxQSXlFjf9tzdqVL9Ktq6Y/wx
P/EFR0tuNWuWHfOGrNehyom0k10p+6wybZ8md9UPcmh+/RSt7QQ4jaJ+vYsPRyS5rPnIEFz/S6uI
pH6xQYOE2v/TitaVRNzVDNT1BH4rt2BfgujeY1MmzarOoU4i6OwSxD6yrS6vXi8Vndk0GssRR4yV
FWbJStY2YE93ucv19yvat30CPvkDDbunTmQ154zKgQaYYnm862QUgCcGXn/yjtzKxxTOrMZtrp+I
3/OlQW4Jf0uvSXuxEyOzM/Qe8vmsuF5px6AVzAOgi0WWI/iXHZoZSRqCtyuxC5F4W1J3ItiBF8hI
0OD1FmM/7kJLgPjMkM0muisml0OcPfW0DfZ3+UcU/MGmdHkCkw0dz+onsAFqRtI+lZGrUw2RkqQw
KH89oBHW0YcKEc3eikGYdBShs2aw5t4kd/z5X/l22jFqFGjEdScdoetO2DMaekGF50q/KVlr3dDr
uA0n4C3jwLgs/R+NM37ZHWqYrZwBiZCQ+3VPDNUk/TVPOOfXAaNiFd40NPeX3bAdEaAHXkdHxdwZ
HIKTHI8Q9vP6e0oLv6wLWSNPUWXPOfdkwOCPjY08KEfoGcLmn+ONLE78Ep0habIndPdGyS4CVP0O
evB+EXzEzdhN9xpIpcMaM4owqNg4dwbFPegF3t2fFLAHHL2ZQu6nhKFxWRz3uj3IQKcvWhfLQ5aq
QnLlFvN8NHfoGa/lRdgUG36xpPcAFq1Tm4iXYfR/F+1y9j9vFXYjwDCsv3S88O7d7M0XuFhhRlbd
mMly6Z+WRoaJLrMd4cvFu3zKWTaApEHH0Jv7JmLQXm/TvFE1+kjtD0YakmZO9Utf1VCU0NX5qFnY
t4CLxMU8KzIKmHaQVU03YAGuxPZUTtKoVvt7gC1msOyeAmjyV9/SzbbdshUkf20VlPZXGhEV69Gg
hcs3eq6QYwroH/rYa3UPL4OBY/ooBYSawaL8gSaAva0x1SbLQSsmb/5ZuE1DVMMjcpmXkv44PfTP
H2hOenZ5ugaXXZZB2AMhyIKArjwO44iH1ClS6/Tw/T4c7w/nS7QxW4aAnMQhYfQo5sUkS3dU8rDM
J7XkebSAegkmcc3woStLUNKgqINfPg9DuFXzf75SLG91GbaMeh4C8QgpraE7wEd7lW2Am7LHo8yG
BbkNe/gDdycUcbBLuA58YZLZvOqjcsox33thAtmsIH1k6dYh6FHwvvqcacDgshNufc5Mm9zROIJf
Gm/KvQxALUhsutZSl1irBK8DDbz6qfsiLEpJcK8tgXJVhhTt6xnoV3QfeyBdgItQclw+QRfo21A6
SyAYg3kc9QveRrzRg7QXH42v1r0nTImCP0ZIRanMnMo7KfO06zJgCgk63xqThiAVm+4RKBY9mH8X
SxOO+N3iMKd1hqeWU+6gnhIsi2Kfcx33o2DKTrr4qcM6czjeMvvmjk4iitDELEjS5aSg3ObkAPc3
CXlw05ILKEzOsFaGevFqZ6eIQzrz00uw/7KBS+e1B7oumyURHhS7D0iesX2IdZc8PHwm6Q5OeHJp
v1AoY1ud0n+U6rsazV95fm5klNvjFOFzxcgRvlczEeDJlpltjU91Y4M6MFqQk5gbS5h3NvpDbvA6
yPvrLp0jBjKc0Bhy5TfQllBBzTI4lrOpi7LTysEwo9jYAuhv+6v9h4f9+RjLdHCognMNIur6e7u+
MtLEV33EFxBglZOxRlrMVo3tByRk24Qh09liyfd23egHrtEQTeQBxnfLTbdfG3BQtF3fyjBQ79UF
L9A4agT/M2ZUAeLYSlMtpr7cKK1lkGe9q2YHMTO44ZwPdpc4/E307wjxgxUwWN6QHrMAXcyXvmRH
84cw9gpgnBhLAC8WZFRyVh0A6n61KWxruYhrwxMRAv0jGi5zaKW8V6INb7Yi1TJQWIKDaITETWQx
B4Fhw1VYN9iqHz8rMcNoheU3+zQBiTWBQ1reW0nbfWZnZSg/BaqukddHTQdLqEGOEpfLeDE63C3x
9xVpTW4qO5EiWtibgOPVCUkxGGHVHa9h+lvu0U7XQAHyhrNh22UT2+H+sneLDQKTOgXA+ywBQWeS
rbf2dsBJdqEr1vvIpOhMi9kXtt5k1UnZYYfrTzHxvFMx6lp8+cIoek79Ij+j+rlBIaeoOi19diTj
6C4TN7FNuywcrcbJHLxr/AKPJ6sRKeiKk0iZAG9AqVsUO/ItUUgO6BYQhRDGTF/yAJluo+iapY/N
BNdmkGEUTeoA9mHKeqpwiPLier/8dWOEosFZvRQNlfQB5EVa9FfBs7NuHjCE7P+4zl1MSTBFToHC
6Ogzchn/KwGII56bo00n9KuiY2Ax0JYeNT2cm3LPyiApDmV6Cxuw3Q/32lqKmVLHmcY5vlo+VXDQ
l3NOlFCQbTsV88a3WiBkpytyQtduqSGhoVDPj0wSfV5WOBGIqP9R/z+X5RDX1A5TCt3X96zPyL0i
qSVCG1NV4+0kwHDvoQtLZVNdCrvWtq1JipKZNmHr/FHGBBm3EN+1QcEdBRhsvKvTAF+zrxBx+qpr
AoHZUpeGaZtP0VN/yeoD5ixmXXZfUOCvxVUFM8ISsguA2pKy+Nr552iyVA7xMYGYzzVe9jYo7nay
6TPA3BlQc/pSJp0vm60Xr4fr2Fb5Vc2c0AFrCajQnp7QDWloreAe8BoLioKxEJdRXAFr/Z2SsJVg
M8cl5eV+VN5hJwWvcPjsA3xXqalYe55oe9d1Fe4O6QyLv01aIqY6sjp9WZpsGYqe1VCSbOiG46pH
2LfbpmZtuA9nmEq/su//aI0+IcST8om+8DzgePxi3OyIB2oK+HyE/6AFPyjtwM5ws60HvIchbekr
2+G7yWTT7Tj3ikuRAM6kaLsQM8iDwTZB0VycULc8B49O8uzaPCdgBqo8TrgSQsCjWv4lL3R8vJ1g
0/K3pV5lMxtvz9Ja6Pcc6M1ELYWQKQtmqcwiqV3JEt5f530R+232y0q8C0lBhh4cKjJgv6mW8qY4
Bio+sH8bJxVHmMw5OGoVwCEyg8VOXgphlW5SOcF/VormDJ8vYuXksWwwVewRhhX/fAbs3OIn4O+J
E23oFatWh/O0qsWlCaWulG4QY7w3A7X4lMRf+JsFPUiz9+G1l45VdOVQfje3u/tALC1otkoFYVjF
5kh6J9brQ9rGWOLLdV4i4QmzLQFwo9FZEtZ1EWC68A/jHiWj69y+oh1PRkKh2pYJe2irCrsR+YLA
Sq1Yyes/a28O1P3qlz/WRZE8MEf/dVS8xYhUzOHektYzlXbW0hYTRNRr5Hedqi40Z6kB4hrkyJ/6
S0GurE2MdDeZtZkmL55VpDFqc2Bk8+ag+AI+418HMr0nuvNua9IM1gnGoQH2y+KCtsSGHhDGn9CZ
DsqYc6GJZ2JStrVg6JKOsu/osnBjzFSYRjX9stMMxMNHh5mH9pinjooe14MzLyWwrY1xkFnKvquL
Z86mHkOp2PSG9uxWhbLn4+ESlb5Bg38wFW9bi3prQkE6J79tEwCEnKd2TbuIV0cC8jWrtaf3UA6r
m74KYbjbUWwm8aY8pNGzE2AC8zA8vPBBEgq+WPS5twiyQs94MZuv0fjlUiY6WziqAYZO8rgLyYrd
7ZREMT5o3H/rUWHiAHNtBBjZBaH4rNS5uce976ojIUWwTSDJPtvVOBBU7sn/y845Joff11amsUV8
F2/Kl80I4O3rWpX5pTVhukrfEaEfPVMAtSUC9gDoSp516EQFA2WsN5zkOAnPusIwf9XgHfpLj66z
pKV/tuI9jTKJtMtgTDjQOuxiNuEFloKb+n19mY1Ri9cF/DvqnFvXrKujlRypmK1ip3WoiccbzDAA
49cFQz1BSMiUM4j2Ywp9u3Iw9Sg2TLcCCZc8Y/AqUxoq5rhSdPADMYfMneT35BjKfOf9AiUOXube
YFENSYFRkv5QgGn6euVA4E6JD901MUoI8iq5U+ofPwWZ+gQmYu+LfebWGCqVQmj7S2pecA1gZo3i
yC3Ex/RZDQWjFKiU2ORE3/0KIq79qP9GPpYqmYmk1r2r/HRncdRjzwb7th3/xJ9Vc1DDNhjZL8UL
uB5AkcgXQea+sb8e/cHevvUzGErRfqIswA8yEednH5x28o7FnCZ9W/S4NvmxvMrgg13yMYnhR17N
ncphBwmw2Bch47nSrfXsemdfcSiHsNgrrfumnJpnHYirLsQQSX+elyoUfaL/fk/AckUWrlq/Dw1Q
MeiZPagsV4NXUTWTW4yhcSg3kqlOnQ+LDMxZ/SBrhPcCBdUoYLTGzrOFz4jZs+Y1yr7zfrvk5TXl
yl8a7YJyUcOcNXcr8+62gLV/TVW8vdmZ3mfi2flAWgFRbN3/R2cn8IC3P1Pyaz9tdS0k3l4KQgGL
F4VkjiPOkOGnfoDG/6zWG1T7Llpnngf4p1tnR7RTiyoT/+xpHMnvx7lL0Quxd+NlDXvTwuJYzCd0
28tYwqm422N9XkHCPDfubTQCVuS1BW42gbYdzjnjHBoco3wFxj8iZPYXjeahjrcbWP37lz5KGzR8
SmrM7P9e/7ekQr1r7MN0i5iEnTlnMbY50OGKjP7g3EVIGmJ4QqW7K8GxH8s4lrUm13Ya3lRrE27X
oxIZEh/5clyfELjgmrcQx/OyH3VP+LXw93ZLEecT0MjvMJpiztHy6bSEwNgjCyz/wbEb+u9DDwo8
+7x8MNtJ2ny16ggZTbiJfbCazoWS5JHOFdKEioxIuoe6/Sam3flj5wF7iNjQXwoYeo+25RKkNfCm
fRwD22LfGBHrkipQM1IfF0SB5QCP4K6QJQIX/tdyyhXjCfXDgcxpZiklunkEmE4BEmtlf1hRXB52
v384Hh7BN8GD0bIYcK9w4zGK3BFhip1hOpizm2H/wJVjXEHtwq52i97MNmhL1WpWFZ3Q6OrDzIxs
/yOAfrczi5wDek7ocyEnXlatAjX+GZAZahUjKs++tgBIN1JA8X6ydM1HFsnioF8ZIzAKSu+K1CUR
8LUvNncY9PupnSD1drkEYee1CqYYzk9TZzinS2AwE0M9bRrhi8Re70R+QH7ZJeZrAYYjcJZaLETC
mzPnxQuqQUMV8YZTitd1Mh5jc0xLhCa2HTKev3fk5U7SdmcgiSQjum/vIn8ASCYzSojo49+sQpGF
gCI0TLtid4yZmt4FhgjzvrWHlB6L5M+oaBbmN6AgEkNfwMhj5by+8rQpdgBzvmxPmkFQ0Zo6jWDP
YTVNSsHVUv4FAKWTikRnD3/yUVxY3spPLE7kxp8gMXzxyqrL9X6OUV33vCCLnZYBwMDf06g5dfQw
oKQR1hIsb/9g2gcw1W24j0QTeNKGnvJKNDHbislp//JaiEgchfYgb9VO/Th8VOTtwOwnTRTr6is/
wW1kVOk5ixeZker/uNcJgMhIllDg2qyZfiMDqfK0pq7RJtPFNzVdKpouR348djfOTgkkuFLpVS77
2W5BXo7hojcIG43Cwcl3x0kWPYPvbWYplSeadVwhhHIYp/yD6V496VK6VXRcs7hHQVrTCD9qLVv9
7h8YxmK75TzUQdIgFzGaRIOnGfvzhagqCKLivoEMOrQpb6K9MPcEF13z+eBk/H6N2GVlh/JwunkS
MAfL40LMJJv4MQwdI9WT2jda/Xidyz7thdRqIzJxxayBer6TurJRWoOjY480QeE/W6LnX98JlN4O
F+kDiiW0wNF5uEgdwjQ4BQLnBZ1zo0VROc7wLlACFT1pagjtwyDoYEOk1QNUr2YThmSivprsVSyr
yRPMGQFBHuzBksHIAYcfdlMxZkaf5ztcI5Q0OqQrFqaPbOfsHTuzWVBNL+efOGm2Rj0Qji+y2D7c
aMue8O29YElmih1dKZcFF58E1a2qFmYZumjJrsR2DlPkgizfX9ZeuIDNlNy8H5Y5yh4beFIzaXJg
8NUA4tnzMA8iyzwJ8KxQ3a2FMYFDCivsc+oNr+JCbqhRcZKvcvuY6gU+OvNly39GNcrZJNnbhksV
9RuMElOC5ANgP3LRPRi2HH0uYroavk+NT6NnROi4/xDuNyKEdlSx6BFjDj/Ze/PhfHsVbw+Qf113
m5N0kpRm7nS0y3sMwnV6B4Sq0yfHh8ejQObLbPpDx7o4knQz2aGFI/VojAyy6sVheWg/BZXN+n+a
5SDCRgUr3Bo6n0xMZxb7K+tkoRurw0rvuBlRLlx48xtGEf4M4LQt3k/xxU78oOsE6QYIgGUlix+I
r1zGOh4BKeA9dhCvIgBs1ooGMExCszImdjktcoukDmxKjw+1EeOHn/4jxcrE4qFIJC8wizbErSN0
MytLKESeT/njo4oo/SgBLExYmcG/XwEXBzEO0Oi3rhB9e2Ed9ThpxUz9RdMoqyKaBImRl4kg2lh2
Bkfdnk++/Dhugi4hQ9DSVlMxnJmQt1xnfjNGRUD4mYrVez6hk7++OSBNMt65zwVR/EKUSTXqJ+59
XHSlBudPyNb6EpaeZF7w0AJm4TiYb6ej0+bb+ItOKTaggt9y60V7tk9n1whzROKgO/6oGGvWQLun
viH6x9jVFyhqgQyRy3cU7xlRStFSzW7ga7HB4r4kArI51ItMECMtW+Pc7t8Y4L8RAbeP75QNeVLr
A7Z6rCLU6UNy1eS13eywAqgM60ygHOYzC4hGiJAIr4KAZtJ1i3rcp3ncVlbijPh3U0+zDnbaSEMU
6PauAolDe6knNuf8ePhI0Yt+KMFgX9mgk5OfmujHDJ2a7Cvod1vFlZd6g370kewxCVNG5kUWnjMM
YecEVSEK/A3X0eK/dQP4SQZfEif+AXUAKaS98SE3ZxwWNrwLxvw2VjjOlzvXAd6mQW1jqfluC5uy
EELY6bofnfgSLBDTvz5wpJvDIR8f/3IzmheJ6f43c4CfuB7KsgGREZvetN/T9auFgTNZO+NB76nT
Q8Qc/hQMkX8jXxZUXFr5imL5OgF6tNbi5Sk88DfFzZCdaF4sR4TvOhhTyrhaWfSbsJpfdGHj/N0U
5uPj438pvvM3JneMAs5R8gr4Z5CaL3xhLURq0uSuh/RWYOSLapEnirb+jjy4rnYAkI8ti+8ijBwo
cF6uq5CAkr+ZVOn1/Pt0SKasgTMNXz+/GGwIpDRd8s+SIW3E72EXi5jYl6zZ5ql7/mrHgjG/MkmF
zdiNuhosLbsd1n31M5oktBLZCFt8eeiMRNqPciRexSHt25lRqNO9GT9rw0cX3gXF6memCoFnnbve
ApWuixCXxa340u4SzJ+bdtxaeI+W8e+D9axPH8w1qh1UdR89xUEU2yVnUomadTJeeQJ0y1xVCPEF
UHcn89FIofyJchj474lZFC+bOV53ET+xfBCW9H7rwHZKfymOiKRpqfpiK07zEvG488w37DVwUtM/
rDWf/vvBqC37ui1iI/VmknoSdLOUY2PiO8ZZxc3BcrYJF7sRJjlI0ds8NTrFP9uwOliPUfpFA6Ah
+bTp4JQGEGOXxyLoPSY2FWyKct/s6i1FyybUe9T38yJcxHwBOZtiv8wR6F9S5ciXBKQGUeEfXP8S
7eqjIgeYxacWcNrHfR2Aj5MYwCeeMapP8fTydYY793PBNvJ7MmvBLgg54czrwjlguSeVaRiTfR+Z
DZUpTKfPTYYKdZH1V32xteCtDLoxszxikSkOE9gr+shRfxJaTkPUGZgmKJjLhHv74Vk/JUdJVEFW
JLjH6ybctSyCQg8xquRUVDKJnNnVlcXZIaFNuexSmZkXXjvkSe4FQHE0bc3qLFwdTMjZeudaUwkq
l44w64XKndWfRNijLo07BQ16wlnDYMC9mYbmgQloglFfs830hJ2PvxoNXm0EDlLXSPVEyO8DKXpu
izPf5m2X7sBsYfvuI0U+hSoZVjTS6xjt67o7NhJ8FywCKnC609NFI6JyuC/uoEjh2YWwi56LqcSs
ps/+rLVYg1eVUDRoPhytD5sBvwxJbKZVQOI8tw3LNx2qdZCAYeteAGgYEMP+0yg1+/OOTvSYaAv+
hUnz6HRstem2hPIptQWm/CTOHYbX/cLExBKSIQRuFR9ja62osI5rn5h4aBfQrm2uFJL+/6mLHfLz
ErBSYnxolXrWrnMIUXvB4Hi3J5zqaMR780FuEA9NJQQXJ5E091nZ7M0u/OhK6eoOFYYQMYOpKHHo
wzqUwE52/AJVTa1QSudx7mvQ541btuf4MBwca9Ksaw9XyGDmKfxQ4uzjomHZyNGj3jysChf44oDf
pDgM4vk9bmBbP2Rcn1yLP071kha4Dm0NMZzlGtpDljZr/N4byoFw9GwZq2yiqSY/vIrTi5GmsSwm
pYomLxCEcWP3u/uo9+BkFanOcqSpv9EoZweK2qdmI1aarbEFfqyMb+7KK82ceZREGfdbg98sjhFf
vTjn+LeVNnte89VWUDzwcCwDU6alPPWld3J3A5XEawSPnyrhrSL5qOj//4msh4INbfsdilbOAZMs
CMyAgL+I8rO5Tcz2ijmgz5fYXIlhE/doai3KP+60hWE42oRgBcPU9v+DAaofaE/7pUNP6XScSEpA
qivHvwNVoPHyDWf+HiyD8GpFqfGqYLdEWNsBEXCZMQ5BsRPWZ+JRPpAeg85cEYkGJaZVsJ0NLWOV
aoCmvJZiEBGQydIa18+yTLo6BaNuxVOV4XzDKUhjYQNhz+U9qVLAT5F4k3CNeaxK5n7MwN68Z3DI
HC5BU9CbG0Nz9mipW+MGei4Z9jWHtQoAyApfRjErNwnbAgRl0xkp8+2lK1JmqK9D2cOH/A/iSEhJ
dO8gKOc+H3NjXr8ukgG2xV3avaA/MmF/uJWWypysbOcwGwPZqWNTiw+5EqkfAx6p/GTrou9hW6Z2
qfmF8UvMjVSTidOYwBJWYNNxdlEtlRG3tyz33kUCq86VoHrVtaowXEf9NxV8EFswvY/8Dn/aah+0
DAM+yEcpGdPvWj89v/8GnuOKKnL/VlcIZ4Hn6PceoZHZnjJv5zzq1YpfEpkEGKvYa7bEnktgmZzT
63Di3rUoOM5HRTseXbYla6Xd5c4g5bRKEaFr0QGspfcpPAputKI72hJYgyfLh0NpB1uUpw/6bmaX
NOpFS5qMy524UmKic8Rpc62/6elGC13POkZ5jm65QcW6/gexQchTfm/8sMwcPdakXHyrthJfYvvG
MZhYCMMtyDF7DJfTgS/magXycJ3f30M7EJi6FZMOFYBdOPvJQmeHQGT39F2VTCZjlBAnTA10g2MK
Ljh7SWP6JTOiTsFJNDb2yqrE1EZm6LdcpnVx2ySwf2NCUEaoikSC7vzlRP29GlO0A5lN23jLpsUq
rGKFuEjQiJSpGry1kjZ8pbVV2IhoTRblsaud59OWmN2chqz6D2409qaRRCKWNKMkn/3MBxGtrksu
EKcqSyHkrN2jsxIx+UML5qdvheZSPAfx39VSrgxCMPutROH0bCrJ6PHHrJQI1VA2+UF4JSA0iHVR
7ur0xE5TfAg4lo6xsRaLUKFd5P3a0117LXOOqzx6l+ONI+kl282QoYPye3Cz7WOsff20P9jWaqdi
wzplgIe3B5rusu1N2wh7JJUtBaqXwDiRzLeQmLqRzb5s5+F5xUTQRTwgx/tOdrL9KV9/yoXq5ShJ
fGYY7RplEZRlmeAXTxbkjst2xIwJExAeZFALW0zd0+PD5itNFqq1Y10P5wieHgBudNNDtJZC9kCS
P1JlOO86R92fM/TsxcINiQmZ5ZAwT6xNJldO7RiroV7b+iTJIH1QFRmBYpg8KosFlOrRs284YwK6
fS9dbGdcktaV6ugqMfbZjfiXEDZmtBb/LFN4Kf0h/hNlUAKHOv+BnQLiu/qvC4OACOXy/VmgU3Rx
t7880Clmnib9R9xeaDX39z4eBUilqLOrmjBSx2m+H5zanufGWS0tznwFtlhjKXNg9DKpeR2OPtGl
oSG541b4aH8769YetbgtVNhkCD4C44YGwj3xcyIdUoHNUKjcdXak/jkB73d2uzNQcD12DP8cSMKn
LUyvdSzCFspQEf0wi8JRfTRT9R9ZvCga3VxWF1tQ1EsRPMVdm9Ei0GWCaJd+C0vLgFvhqagPcUYQ
7qd9SokqhPS7f3PSHZKX4ucH80CaaphmUHGUCXDUGuIOxV9Otmhgz+VHP3uliT+znB5fQB/bVpIZ
5nbz8KGffA0+8Bo4eOhJ2u/u62h8RUulSSaekSSxiwuUv/Xk0n/5AzWtgEiAnaltsNjU9pZi90s9
19iMSBYd53q8g31mDqFFyslDX5BcMYBdXnm2DuRN/RpSGbPv21VbzT0aZRja5cPPKY5ykdEIonyP
NAn8M2BxEGsJUbuvC3sk8HP8qo0RNt/s/E/YNRNXmwsaS+3vQObMGbU/eBFn0+HQJZ2jsa06Ps1s
MTqr1yS3tNy1PDs53QIfSR4tU9KCVxiKmRHLyKq57d7Vp4B1o7aNQxKzdIsgZ2jOZBxbhl27sk65
zImk5xdfElaev8UGgEtuNeNoNr6FALS+LAaUYz3IDUZLSOrdjeT07KlRfJJpi+BotbyRIyfXfKXx
B9lhc3hOZqy99CwgXbbAIwpnAJvPHbANDbIK+pO7pflSq6qrb6GmlwGLY0XCVP5WFqXmWfPy3cPb
N99NXzkXCAiHP/k/RB+XrEqRHWYRf4oPM5AEcgy2jEtE2WTiz8jX76c4BWjhrnpsSgACoSYo/5Z8
wfLuqAZrhrKW0FMhfMa4LdGk7b4JrTlN3k3BCPSVUwfUoU+li3F51kL0trCG5eFzTuF/gsPSP3Jn
VaqIg4cqJcJvRjxAJiyc+aEjDq1kmMoLTQAcQJ9PvHBFHTi34q5l01uRIrYX4MHhgt3VA/tmW4F9
DniGfo90DfinNFSXarYj0+muWnqCSQLsYhRoudOFQ/Db6SCkCmL+9r+J2wIoPd/KF1kbz9VNtNYk
/f2n54ZBQJBNdBYwp4uIp/ulr9Wt58d5l6L68ourm9p3bBkaC/FRWdsPGOOmP9zaWmMnz/bP0Wvb
ZQPcmcMl6ey8xOl1c8tK4caJd29DXOc7O4W6sq1sYPGll+yU5TXck3V0KfEHR05n8/Wkb3tZZJAk
xaE0fdrpmuy9M4qkAEk0EO8ISfe2zkGsKzHIa0+sBdLDH26WLoqInL8FNUcOqFmBZvTFodMpqYC0
RBrYsqX9u+qc/5FTcegXiicf7w6mry5lWjZIJ7yEyLWKH/7UsPqgLrOSC9476eDdscOmlTFaScC7
LMAre1xXhk2RXAPfzrd6H85p8bBfH5Pvum64UXGJybDuMg7b23CJ8n5gkxEXBauOhHONrA1JQ8nO
hTydF7hGcRH05aq0Lc3Ek4GU5CvaMttkV60R3yT7qKSHMwbiGCy3SoLR25mID3nY4+dKIwe7/ch8
xn1WDMer45SyUxzqsp5sWXbs5k9c4nPz2SFq0s7JZ8aPeh0cbcy/GI0pFcu87dxcvurBTYSy1WtC
8bHiWpFS3+MyxLlgaZoGiaL1vRJJV+B1XMIAFjDl22gKJkt/9GKMKtKGXbrfMHb3DI55rlsUPG5M
YF6wkNqoGoYBHToJiInsADaH6TnLZmkbK49PaZuNZx9QGcrWL+ZVBV7Hv4nHScEQLw5KAHQTDpC+
4EimxDcR+OuvQ9JTeyOJRSr9Qlt1+MWsxYYnZh5ofw655GYrTEKOWHdZ0CUaOpGF1E9nj88DB0GX
4j0fmwuD7R6Edaz52J0GDlyAd+i03Zu0e1H+gdEvXHF8DJHetGl3qBqAjJUrci1hD7ykYQ2bY2AH
r8prBDipe2cYZkLkAYSrc2DaDmuGYI2YFgrxHyQ6Hv7QLK4YLYrxq3PCNozXP5vLcW5D35M0OKOO
EzPU5py2kubL5PJDklaSEXd/fA585W6E1966hH6AIsJ1+ajXUTalVQKiz5UXQTNzDbx0pFYrSH+w
FloOfK/dybvuXln37BsEjaL67lIndIUy8nPrTB+TVkvFiCk2tw0+lUZF+p8VF/1fNaQbcn2cxntP
RGpCR5ZmS7f4yrMUcZhOorUH51JhLkoNb3McDdGveBUDI7Z86LJvxJ6eQ9wxvsI/7NO7FNXUBNB1
cKRL/yWzHO6dp/bUILrrzMcgwfDsFv2824TgSkFXsmgC6F3Vw9G6MuQNqU0VInkWKyDErnbSr3yh
vIceZY2fAn5pEjW1f3CjUm/tHYL5ZEOBW+uq454H+SHnPBdRPjamUAIc/UVI4TyOv/11GE+7yNaD
cu90QUSV6DOVYNVJ/JOPkc/jbsXShpckQ3daAYcAWUf+M9i6cdNhWS07kRtNnyyCQUX5Q8tfrfsH
WglgF2j76j44ofSggLkPp/c3vjsPWplU48dDrchtf/eKT06spntTb+6BcaSXmN6sXVVCMRG0irEN
jgtIVopalHp4aX/GlRaVXHqCjIqVj14TAt7IIOYXek4/QTqUk0MbJKq7o9SrWCN5NL4wNZuAUE1r
nubGPaX/i0uH5LUiRXfE9mIxJyHgU3QOXWJTDs7lUC7Q0L5rkH8qc9Tr4FbSYJjK2eOwJFoxELie
eGtmxtFxW5dwcq9UE+OpxSdlNfrPpU7/k+aYIZiCudn6xVf5SKoesc5oi0B4Z8xYycfWJCz8eiQP
9K4j5RoVOMiykTyYGtqvU8WDYjbBCo1CMMhvmg+un1xTPJIBn//W/aed8kSvZYYyXdIAmU2wMQUs
j1ubKtZtEvZUM042yf5E0G5wG+aATcHdk2e4HWtzTqhCXMsV1nqt7+8dG17ShVtEl61z490roR7F
LT28zDUaV2EVJ6PRQP/NYoeEJ5E5LlteBWIbp6NmsIaeQuPNuX6BivhJqmu2TZTOVxQux2bawnw+
PygzBfbo9F+37vgX7cwQy3RUZc08NF2eQnRjuJ1s7MLzpk9H8XY2/0hm1Wrb6SfCxRQrIya0CTf2
CArL7Lf2lCVKmRt8aS8K6sdfL9NtCxGzhzzw3pLEm21wVs0twpXV4P1kCkJLJuuq8wbOZJmk1Vi2
r2FY5ke2pz+LV5lRth7uga5N0O8FMcnsBMlkO6aeVT3+8bvxANqeM5MqpmaZcPEEQFie1Ws20lC6
zz330CFoFxkvdvcCycJPn6eZFbdPIDOU9/G97ozUncVwfDcytRk0gY893TLySiPMmVWNSs1MrvxV
7KvNDvG0T1TMGuBkOmq1HQjzz2o8qYBmS89LtCMzvroqp4+YnQ7A1xgVCmz5NnMAu80YUQ+k012V
TBAFKdBL6k2mk68dBFerKoIFM7Yu7SW17B+LZwECWNF9CvDYs4pJG3dL+yi2ufJ6sevClfX4bNa6
DHJ9Ilp43LGo46K2cQ4V5QRHYmtf08v3t3/IlPNKUgBDGRqUVGx2Y2l7TxUQtIyM18/ak1v8P2CZ
cAqeCCcuQMyx8GZEVFKkJyHxOiQhh801F9CvTpuREO3Y3wfz1a/kQtqoufcLP7/Zfk6B3TrekOOc
0D8EzhXl3zzbsz1Qur2WW2pwFUMMUpfgm50hjbfY9J7Sqb+8WKEutFWcImCHPkFLFfkousFe3o8g
Lmcoq2Ix5xfIGuz1qYJVtWTabWjYJHOpXARMycGy1+cV1Oqo3LV5jnt3/ZEZNn7IL39eD153v3R5
sXTg4jiEVR5T3RO5EnWY86ZLUoxTRJZ8WrmdleZ1eO/yS7W75vtx6Kr/OHZS7lL5/oDASieehHLl
ERCx1iibnPPh0pcoExVvsfIFEwcd2sNLcLBLGL5GklEZzdia6zpA87rB3w033Ff3I7D6LaFp1ZAB
NdoQj/qsK951x/YqGITeSPyUF6U7RWRJ8n0XsDLsiE0Iqop/KK3ekuNA35lFLTlM+6qU6AAj15pq
t21iKaWM+gxtzIIVsUCDi+bxVNQDdrZrxuva59jUD10eGmNijEiO+64dsep03I/ZP1e0dnRJDDAG
CZ9IZUKkbWc9PbCiwzvIGuPa8uMBYZde79aV6jMAI/s8NHKkaCG6VwYi2M8XCK2/U8A/l0Lbrlg5
DRw0vEloMxvoroOqG7/9vG7AUxJvT9fR4Qq3cSkAdTcT5rbsc1Dk8AwxOKlRUK5XoFsmfVjX2Fsh
d0LAL5G1ZG1C99RxICYb4MDLBnSWudjXrdwCvRRPyW9Nw/iR3eLCqMdHchMslILMpBaD5J+s0H5I
Ed5EjGIuZcByQ+OV/8hJSJ/yx3k2r4c1WuZcSE2d2FOS50DVNZd2/Y9Lt+5q2uY9Ujp6OjU/ULhq
ZSBqFKJ6X3rF54llCABlBSnJfk9L3IMq62vNiB1eH/ILvIGiFUbZtLxn841CYS7J9sOxL536A2RN
FnhCLMzhTJYcFLhBL3RWJkXYtZDjvrdKBtEbTdGQF6RuavLiFbK+VCI9EPwglsVa+vPxYHfd9z4l
Wct+doyMWQxd1zlw/fDy0WriH4SF9dqBvyBMsSbew1niGAU4Tpf39NgtjtcYgJtWNimkDylmR1VS
hEqUI//4NHS8ts8oQec+kd7rJndVGq+bFVgru3gKiyORd+MYuovL9sNshdsuaRouagfpEd1jdx1L
CIoCoOQdDItsInJ91ZyHzUpH6jWkazAPGj7litnCVd0QakGdWgFSw86CBqtcQM0WyjPNi/gZLaCJ
sXBUIX29Rwd4CTmZU9T+dX8J1oOI1x3lI67PGPz9QIrg67+n7lsX32eMAMyLITcMYgM1lqQyYGUd
MBwTiErEl4FNglj6sfRnS70QvDSv5IGZYICmrQO3aafx4G4lh4Waf1295B5uFnceDrUboPTFBCsW
/qZNRFiPUm4Y8yWcahq+5DHCQrBiPxy4IXcgrgBh0jLGDeYyFzjiLslJijj1M1z3e56KIsS5JFKd
thFMYkGCEeJJY+W9RpgLop7HTNVrBm58Ku7jv0ec4WZcBJeNmMvDx9+TWq2BCKT0xH9i4hLbmPAk
b8KywFmE8CuAhqqhQfZGhKSYd0rYTiZOioVvCghcxDPAH9SdiPxcysTmb/BOTqRlP4Gw29g4mfEK
fP8xFo5gxy75EUO7RFhg3Z/71gN0abMpRPOSiv8aphXcehwE4A0mUGOkFrZ/2oHKqc1elkH61uY9
QSQtfTHQ3AtMTqJS1et16CA9luOITJCpeUI+3TfxhzsaLZS8cxqHle5T7pOtFdSaJkj9QFEObjHi
LScRVFdxmpvrEeTiPP6tIVOYGOdDWN5uzMAoN63xiMto9dXY0tTabCY29lQajWFzxpSUeDadiF0U
cl6zyMTEbch40sB/WLWx3YN1qppQJcBDdIhYXwu0qhr65PHFxdQiFihYtsH4DXbz9a1hAmxTLiwg
zhSVORO7PPM3XZDL45GJkWed2/64v8bdeRWcBTZENvBNAXZA8ge2YL6j0h5yJn6susCxHabSldUg
m18J8DmywoINwV1YcJpo054WeVtJlOrQozHF10nOCP/T7EpJhNHTuuvxgDjZ4hiuvm0UTbn8dNAK
LqOgaaOPCegHnlH6yPrd9KML2FWI8+xnsupGquC9KDqUWrWIgU8CsRuLMjODCWM61Q253PCskYRe
XeLMM/DD99HG/SVgdnxLjM7ewbHidrOJnILgRlA6yrDCueSdiu3v8dC/ieWM12MZ+zEl+hLMpbLp
/EtlihokE0Kr+/Mdsz3/S+gcV9B2rUMrL0b/EVx3nCYQxDZggCHL5UTC02wPQu61a8j8X6QIDVdV
ku309pwkCV9B9+vAzD/o8SpgUl/NpU+Xh4GYx3g8bwGdHL827lI53x+U5EvcI9Y4sRr+W8hv4VZ+
/wHTOQgKAOBCbsa5FehjX82YrbvgFAiUHw2uttlh9Exl2w46jEpjPvdsjfh3SSRruMlxrNJ77xIk
vPT1UnGHOgmJZuOJU9Yj0ocu3jLpDZBGgE/w3uQncI/sNX5dlg036JffFfPhUwsSaiZSqX664a2/
TYaPh/InAGvi+RUUuoIdXRmZxy83XBP4HWkAAlK4IiSqNW1zAURo1monXkvzcME6xJ9WD8FvPl+l
x4OCQQHQL0GQHEJIoCbHaIxqsIQGGzlkYMY/ZHg0IQgn+8D+J7tKXDvq9L3CxghfYnsVgicZmFWG
VA6Sp6q8tG73LKbv18LNg/XOniZPYp04XInLVjs0Uhf/PnTHmIZDQ6ou0C0OYZSeMObmmSZR9RId
t87ejDmTxB+r/Xhw9+ENeh8ds2czdBi2gTrbzhudoB2oeLOc01eCzPGSLY6tAZlNeacIIQKJmGpf
ZA2NlT8sgj9cipk9D1XuaFYbXTCWLERjJvM6ZO4n4JIhA0eb+nGJswPJmH3OiELjHpi/pbMY3RSt
rPBCv+COmRcu8gjnL6JsTr7pVmtj9euud+LiZjuNRe78zIXwoZSUW3/P51qG6tC4nRyVb8InlXz8
BqX0Vf3faW1DGT3IE8DL26RL4u3z2d6OMpDeWFUBgq73RWDW2moYsTZ6PZGhC75yIka6KJGfB+aR
oLhPWhQKMDBcINCcXkh1CWIVve4QVvQ9SSob+A4ZxB4FjEfMmX9gFHHxKSQvk0Qu+/RqkXgmHN0r
kRRbmqgnyZXLw8oGE0Z+lKpjBMMPozje8GJ2fLRVEb8Qzi1w+8bu4Z3APosheQRPxAYypt56KWv9
ODNHdKr6iv+4Pw2WXbgj61nqHcXNToiLtHy0TzzgsQyNk23YVuIwDYb7pZMnlVHu/pu3QTsId1FJ
V48y5M192hKWSnFEWMDqsHtWqbl15BJn6HzUSTzyySxzZ2zcCCC5JAUtfnXrxCsYVSj+Wp89yStX
emBNvxM2muBHD/hK+I5Y/FJ66ny1qM91vlMNfW5okoirpx+p9hALLz2vm7TD8pl7PksOsjX8IDkY
2IZvuGYR5xMsO2dcKLupqLptHZOQjZoKcP1KSX7BM93ANUdXsU7SgLlDmn/FhAAZ4nPs3JhFsfXS
z1Hu9NTy1TxBKgPNpz2iITAAA38ASAx1G5Q9Ieba3lLDi5GFMlRkySyPLAnxsZOMOSMqvlMpiqxm
tg4c0ffVxCqWkH9/Q+CaETTsABU8ifwfXerVmWeYas+rvHYuba3CxeZAlJJr8e4AtMxXjET1jp04
uIioTvzf5iTIlEveemKMo6cuKAV+h1ZSjZDeHJsQYlvmMEQH5Gm0OoKblRt233aNVg+tFFpvlr9V
oyyuuqGF0Xdz/Dq88/ADEldI9cZUqWLkL3SuWksb0yeKhSw05rnJwO3TJ66ao/yjuE7VNSIDAFfG
1mChqr89rAoH4gbfMcUj2zfhAO8gaKrpdD1oSMZh56NiSToCC3Vzjn6ay0zcBuFM4Qfy3BcMYHdg
jEbgGfWJWwwYm/Cuv7Hz597seGL2LKt5yzdQsATVKdZjGBX+ciSQjdEWRgVuJuNaXu/j+ZSHW2iG
QLETnKT5KmWqrLKhaSAE0Sh1krgQABaT5J06eJh9fIksvTaaYu4n7JIBUcQJMWaMTmk0d7Rb9X7u
bYxVc4mjYTShsSm+LMIFzoKnQ2PGDr6qfafiMQ1XG+E6HKBVVVlSSdJaTtxlkxELICUG2oxX1H2G
wINkFttZTCCmLUEiEBCyn476ojyfbQd25kjif4NO6yQiEk2wmWbiW3kWydyWT5uF0XQqx+jLGm/H
GBErJCNv0ECHia7yWsfYch80s3jY3ZfnTeOmTdSAio9NTf9G+0MpEH/mQvbw2fDHjMmHKrphYnr+
VejDWQWN5RcO70WB9HAQ+p+7fw/S5ctdshE38kHTD+ZX9Iy5VzWiQ3J4byiirKZuDoWcKRS5aBja
P22aZKG2MZl4TaGtbPMiEaBT44ximhcKlalWj4XkBHE6hbr2LAGVFgj/v7ii+CCzkhT7gDqBCwN7
R9xTT2imsq5G5b0yFdG9azqTSpDu+sRWVG0Aqji6XFnKShePevxwmbzwB0Jz8hqH7xy+fW+wMCVL
lxFwbM/QErnd2KUb8y4ErKMZbAHDMQyZ0QJ+Izz3C5ItjO9aSWQa1UADYIFlsOk+uJEQcFY4hTYh
FUpak5Y6MzjQAUr5PkYsMVMyN2HRhxSH5IPvXMtwUPvJZbILlJZYe71uryKa8RDYbadsA9D279xY
k1TD1mkhsi+xtkjbf9DKWuVnnm7b5tXAC4ifGjDdM4zsNQXiv6Uj5pNrKgwgzFKBV4kM+6J/lz1G
kXRdCB094lNF2OycMBVmbr3jecQQFmVM3lrZaPqJQoi8yVqLcz4YmfCSBtS1bgtHeBDveH3CN9lj
Y0GO8Yd7iZ+7VZVu+WMQecXgDO55M7xYGK6o6kOmmziWASyAGdocvuJOOoEPg3vt9lexZFh5OOEp
EblNVECoo0uK3RmSWdjhMu1AzjDrlg4X1QA4jftDJmOSj0b1kgyRYRtZoxFqxyxdxHoi3Ax7Fs9G
wgvO8Cu32mfubranzgp9f2k1Tcr0D2UUoZiP5HCPpCxqCPndowjjaEQlsKoP3VE83Q2B3EHl1gp5
uLJtA/NeKCpgRfL8K3tdHQgsA8WkZNJK/kp2KwWnkEIQxa9Hp8erNj6VWVFpBb1qyKa7XaGDZnHV
YqHIQ9snUNMsymYESRC9YD6BLsjEMN65xo3GfYWIRKPvOGFo/Chr4neNQEWYq26NMvOdarPp3PhG
wwK6UX/YpBPUIhB1pqKiUWkuM+3XyZwn7s9GH3IU7C738BrZtX6LUn/MULlDKQIu5/AZhW/S3pYv
r+6LuWjk5S9DbOM81tEVcN67E12QTzrh+ySndWpmhf8LArjjC7sZtni7GD8iPcvdD8UE0HRo7W0W
qPZgiRKnHzbmFxhSmxJeZRjvzmlDWn4en5FrscalLCYXLEYTQ5CrHFomhwD2PcE0b6C4Q9uW3xFW
g/LH0/ofe4Qr6HYjciBGiN9hydM5fW0qkGBeNEREpDFkLhFMTPJTCTeW86alDxSK0sYiLC6OGhNr
Tt7Ytq/frMiCyTsSPACTiEuxQNc7WGVEGDLkgDz8ZSHDVA3qy88y8r5qxlCIkxwSKc+kweCO70Yw
mZ5QWuXeS9Iz6ecfZrRWBH86uu7pSqLeDFsi+jIpUuJq5xDp35ypqaF6WCKc1HwN/x5HUHELZz+/
/aFyVjk1kxZUE/CeI09TlrmifjYfeUBoZF9SNZb9M2C7buxgqPPZdk7k2QBtbCORk6EhKcq/i8PI
jsUkbfOCtK/Xd6uIhEeCEEXDnEsGE7ZnS2YUmrJ/tl7OKOw/vbJRgcUxWFIVD89H0itwrvM/KEeR
ZCRrJ/dTYxSSp208vltc9etBtUsnZJXRo11PqGYzBH+avxgeZ8mXaWUr+DQdsNICJEdfZwxkWznr
5zHiSOsOtuNIbzT/gNS4o3wj1+eu63299xsTi8eYrWSkG7jHpru1+jblCQs9rwLq9dv0ZDJvL35Z
03oOsx7V7vGwOjm8VivEowocjOUFX+Y0Y6wki0ZImpS+/FCsNSdI4tpp45EmegNbsUBUQ/5xAN3E
M5+AklS2Q1Tc1dUgODIrc8hQqHtY19xc+k6N52uhBDCBArHrDmy6s+QSI4e3z6Su797/9HJzzem3
OLyATUuXI5W6ydkzAxjAHZ4Cf8a/FdfgVhmbaATcNgTwA/wdWInxECXe2CdGdQyvyJH+jGUu7UNZ
/2nY8BE5vmm+DZv0e0LNzAGE3p928DqDPK7n0Q0W1hFBptoksVpgUpnnqpVvvOmjroJdMKLhms4l
+AKIVBvwgm+CZVplR5p/b6ejGJmiOKiWfuYyQrebtmQneWjZ78D41EAAWxD9PBW69ZGLw3GZsHTe
2u8zdzG40BmZvqyoaslkzBUqLyyzXQqi14Y40SrkITIPliJIUZR5FhtkPNZJVY7TzFxXohyAMe6H
/tkapa6M4kN9pWyLzRro+XdRL0x2yWZ1zM+v499YeZPPUlIc4okpevfUoERI4DUlhb0S97dgu0Sr
oAjINEsVlITrvpPwYEoS/NFF5plqomD7X/zhTEstyKASaDBoFIN7+5pUlXDOU5BlVS3bTJZlNgmK
k6jo1WIbnItXNh5m23ucfee8r7youG11SH3u1FST1d2g35fPLnx/R7ZezLQZxNlWA7ZNa8FLbkjr
8v8XGRKWzuweavFLYC7+L6bgplM45ohZwpBEZKjs1ZjgmvLjkiUbqkwQMKNMDbbC684+8Az8JNQw
oNm1zZ8Lzo5V9L/qjLJ5z6RHqAx6ycO6xdnW0w2cGlGfEC98DW/t7+F4cDNWNjV+5BQ2gGbLDrki
ZYrClfnqJRXR8aR0WhOkQMMdN1UiHx4pLjDJjVppZsulfFNt7m2ypgF272xnrUzNP3CkKNYBFdKV
S9W80Weip8VMB80rZIIMZ/GhyXsCH/JBQxnCI8sK+W9ibN9dVzHjaeBJmFYQ/kfDTJ6lLya6l0vy
p9btTaQIEFYv8fyJQI6wsPmesZWiQhXNxpAX8TFwEp9ToGYTtIFRBL+Wqfk+ttc2AstOAZY1fxEj
lssfqjlelxEFk088BBjisPwL9FD0+WWzXFUv0YrRvYdU/Y1VE3xD+Mcobx1YP3w6g+BJNyJDB646
gjn4eiElbQpdCGPErW/aWGLoTqT/UjQbNzGAJG+gABuJMSMMb7FHw2+SaTiN0gxt9AzKPtKYhk1m
IJ0NwqOyGjlfSEaqlsKcfD4ikw9iRl9dnkLt98UHppRG0ihvSggAoGhq8AYbF9dSyDpH0IpEHQBx
04jMe9FffgXWJoI/h8S51G+Aurn+5ii3B1DwObLMNXXHhEbg5jFjyX/ry3UrhqqZYdLsYWA7w+Yy
UWbjFgs7DEO9SyhhhQF55bi+c/Uyw6C9m5d8PsHeZvjhI0x8HAEox01tqaEiqdI1qNsMoNoSSNyx
tol5YQYxvlOMNhSABpg/t7kAUMvyamGMk73sWeO88j8Q+oCYcuER65klY1BSMLvrbDfintx4Ozo6
lQhwLjk9B6Nht2PaLFkkuPHvYvQjWZjfC69aM9oCMuJ55uzOFtn23m/8OirQqnTwb1zQ69THxTnp
iK23/h6h3BB7Bw2n64PDAwod0BgnOTEFjVqd9SgrmDztQiBOtEg2tXj2kb3/oLS3X9icaes4dbxm
950+EXyAE7f3/5T2reeqhOr6mXc0+o+bvbMWvR/K9DnNUHmo8Mz20p41Sh2joylezNCHh12bhkAA
ln+db9EvFUV6UQEj+dA2bulJHFvd5JPd5npyzenQzDUwhMwqCWGzPKuSp83M2sRYQr4qhis2Ulru
bZ/fpiT7EQ81b7zhex5wsLg9JelDUvbWNawbMyp7y4lIDQzHV4xhtZaESuBoNtGLTsM+xv91mvFf
qZ6gEDczRnboWjTXmVT0646vLcA42Yyb2/GleJy2eXWTEkTGZ/CJUkhyF9u6AncTGJqEbahnM7NV
v6FVULFhVsSuGxOchwTln60a8qSmljNQou8ZFn7d1Txu8JfP76MAVhs0aA/k7DG8u98+OqJ8cqCC
eUNyvHtHaXb6Y2E5O7h79lEyMZUBnFd5QZyOL233DgnqMC1CGjgxY+9P7wKNe8B/zvmdEq+ZJC2Q
uRxJ0//Wz/sZjJCqw+mbbsD1FPHkZRe7jUdho3fVpErCsadW4bKRryT6CuoIpUkqetrPyMfNzhCY
jpO4SDfM/Hs9DK0LFMwLN0viXoyqEP7fpG++7nJt6fMOlCbJcMNp06keeBWgjnoGh92tV6vHFLHV
4YVk8KnskJxzoxsewQAYPZqn825PcmVoeMTWqRL5xDuxo8JAh0ha5MJju7xoBFPTDzaFWDVkHewF
HlV3hM23rLSebDV4c78yXdWcCFOlZhCzBGYqksqjSYQNne8U42zwIN48pqNi0/B5zQRhcKRYHhoG
E4IgOJKVzESM5ESW83fQeL1Fwmv1HEB8RlCYAqRijO0tEO9Ne3KB6+ZrRrh5kRCuzcvFHEhPhyZq
AFReBdP/tG7ShV5NbfNpBOs3oVgaa6/PRuArgH6u2LnDld/QUiyaA3yiIxsUtzC7El7/62e1/XmW
ra7Ss/k0cqm673XQtRKspB+7MtpcUMHiI5ePbIKMfdaNr89gxSCEaJ2r2+HOk5R5xsMIbdSzwaPA
lEQqbNVjcwB0cGaqW1gq8kV4ezauCLSEPiVPbu+hmB3JLiwO/wP5CXU9QMo8yyKGbfPORJGbgK4d
HAvpv90++CujLdzSnd4yEyCxMOM38KieZIGeNpbCDGMG8C4qz6ysAQlfEG0Gk8o6xiGbcZsA3gjx
huKDL4o76ugHCKSP6wiB8GUQq6VdTDKZqyNtLy5z8ah3U24qvSaGg+wOlGSBlG/uw0gzZGEeGvO+
GqmxDFkZ0khq2Q5jv4nTKNJhu2WC3TPfajDfKuQHLb98M0mTbzsqRBGcnICm9cHQzbMRDk+C8HEV
cWalJZJ2aJg02Y5iDCnV6pjfG2Gh+ioBsUhNnSI9cwtlDuc4o3BprnzlsC+6aWScoVvcu75gXHLu
CBvrWy6IFf8QnMbT2x/eLcJ+WGjsjKAJbI2rNNQWVl55MJ55nJPPGt4hAegt88p+7PDj5vFK2VTJ
xq7iKrNsFRMlowkxUmsJG4tNshcrpwDLgD9McnRejlypj/0AZ5M+8G9ERGcK2nh8y/R4tRorKpRb
c37+YS1MQDqkgpkxce0JuiixCzxGXhxXMIZTt+fpD5SAmE7EoMbnxMvPjmSxq4tlt3wVAgFRw1ZU
KfrEgJljSt5dvnk1Ysi8OTF5pSWpx69I4F5uXfMeQ8EFAH1GnLEpY9xkfYFbQT8ecj/yndO5701z
x3NTTqu8YY9q2dyc0JNIbFcGKvKZ8rNRIt/vBxIeH3uev0dr9f0xyK6fwrOXUZ9SRGteUODzY1Ej
vy50cEswcxsBENXrNoo5x5Kugt06I19WD4vUhpU7Yi3jDoAf6uZOSHg4jF+MSwNuFXR2fxM8Hx2O
ZtiEXBsBwBif9Xpf8ZgEIBJzR7iNzQde8pVXYs3BBkP5BXW7/OXzlxTL41eax7Yegz+mlq8UrJR6
ZLgnq+fBKs5s4NxxYSiZeSPtBhC9N0ILWszEE0f2AvTs7IiLswVRvVfkbmL3RW4qlqmXg37GQanB
YVyJeAD+LcWl5x12xq7Dz7IAN/dJ+iMqphEauoYqrmK8/0QFyw5dxT6a2Cy8kICPnDDNHNQnZMcS
kx99Ozw0gZWYqKMm/ujVBc1i6+1urmv3ZEy7Bcgx02rJtPGKFkbJzvNmq5jPVfRJFtt+ewqfta/T
RIyFYdgb4Jk3lc306YDYhqRfYFLMQmizsDos1BnJDdoIJz7KYCbtm14YfKrsHV51Pirxnuk3ampg
skC4pAomSjbvLEcMqSkh++2v+8B5llFbAfj2FPadefslZ+lLQWNvxd3zv+XxmPCd6iQpT5L6u52u
a/HCMsVKcsx0Q7O1e/seX9IUdX3XpMt5NUIqoLcqH+q2+pnhF9Smex2+wX8LXGPTFeF++YCeGMoK
midJFAZn4+Aqt2HdndomjulPf03yFfUAXJSjKbcG/GMjF1iQQpqfZIuf1DBxE355oZJlCokMuFXI
DFOcwUW2lMnjXynq8ElNDtDKRRIoRD9qx1c3aK1pRhCW8nCCMUt+YxhO1gj5p7Xsf+//B+zplC9e
JifcPlKIFdLh2srZFSOy2RKhbOM2BUuHEDZHnNdpFdmv5DGEm5YHcNZfTvZoZGcXNpCBGaQXqdBO
vK9sslKPvdw3FYX1V3sqVJYOQz76dvDbUnZc9xkZJT/bBfMKS+onVSq+KxiJUtsqRb2o8talbPM4
OwaL2sQkhIas9ZxJWn+x8e8S9f4bGGyb2wUuTbyD9a8ciM2LNYeTEKaiqAcXlwFcispNEdqbH+ga
bUrUXwka464NSQ65588ZH/WCMDOe7naOMRvdnSkhqTAbO8iiIBSIypHFYp30wGgtiASxuuy9+ZoQ
lSbdvERE5Tv+WloLzxWKKvRRfxhWJY6iEuTfPSxBoLSe0CBviRXCGteIKa13JumXWX7RTMp7+Hl5
/xs2+gndOrbgm6YmCCPYv7FBNfSOpmSa0Ybpv2xUGrLVD764TvshVbjdxJaoVsq0H71PcTscWcJG
4kpz9qwyUwJZZePCYMYF+cRniQMMnM59IdsgC6bLasQPvRRaogRLld5PcK+nPVFtfAwrOvywYfo9
cIC95PfSaMmEcnib3pOWpVb5pDiOphPJoJML6IoNA21WQx5ApXIea3uqL5mHl1OHGbMS8zMryXHq
poOBKrYjz1p4n8o4JVuJE1pVF82R+9Ybv0nZn+t0s1Iv3o942VisRpNR59ccJ7yWMVBIT3i0qU2R
ABMSczS/uUbUwwEYjEJydSSdXClxdSUFnCdLEky1eXTjFfqIEegs7PkdBDNdnHVTKhPXe9E2OYbc
kE1mOAQZ6VKt6SHBJMmrxQvdohoYwrdcFa6Cji5OP6anQB+GEoXqp/oZbWwGTqIIeuLYCPxiCcrJ
sk9Z0Ip9WVfddRrp4eUDs6qmuXPjli012sfdeDe1xcdj0C8312lTzYTY0Ms9p6IubmsFjohJBvin
g2BVBRkOee0ZA0XgFKzkyyGxwfX+x4XRAjmpw397Qx4XN1bY9fuwxUbZwFBL9hjKC9pZtcL9EBfV
5pgwBMXR3jfC+2yB+kA6QYHS6xydVWP/lsCl/x5uFu81utEXa/zWzv/2i1c8tPW5p9qcmHTViikm
ulMWF/8m3wLrf4lpePNFauq5uLrw7mdxDdI+hYUVQd0p+uz28gJDo1dp03bUWP9lZnVUQGcaqXMQ
EIHkJ4z7NWxNzHbnophlqLw59NU02+jWd6ZtexCrLz6Ip03proAdDUUg4gaZVye0bVYQVkvstYdE
q+Fa3b0Eu/FniXIRi0MaMMDqM4rkHD0c/bsA36tgCYNXU/xMDUCxYIC6/zArWSs5WsQcYTKEmoOs
FLwx8caGjZO6J0oElV7SfbmcW01x8MF45Rli05DRdAtcBJfjR+izUZ800l7srKBoMOERZb1I0Guk
zM39eeG/RlzvJXfUZ7TcaGXw2TkSKlUDFQtSd6uPEMYu6LOjIQInkHKMGTmCef6KfZHF7f/pHShr
wneOlYXrYacnMrfzvJm+wzslSOsdvmuR3kl18Y2YQ/U2/xFF/HYaCscVSzMd2V+zB+hR+/j/FeTZ
1bLYXnY31+cAQ0H48hgWRb8v8iIHju/PKqCAcO2x3UnESUuGyAkoYTZEdPWwpQJ+QXsvFY5wgRk0
ftoPDSNGTnbs2at6wPx5/DODKsjG4FH9GTz7b/JhUaukZHTKMGIdWTAXdA6nJSOUsn3tZ9R34XnK
7h2O63s6ZhLGDucm+j0v/n+AlsszVXjetfTbMFWxz5C5utec+nFsUBXrUrjc2MEX5gm807cSDwbE
UCLPRfL283u+XYTwlpDvtqZJUNhWkvB7gZjnnhGeUBVnJ+ZzuEKwObIB+deiK7H3Ol/7M6Jt2Vnk
WxqaWexrzNsvScHpav+zTCH2K2h/bwCvs0tuckuxMDhVhXDRs1R4bqXTbfdj0C0jwv/CEOn4ykix
yRCGJjz2qtrVGW3Tip6gt4UUoMY0rNDy+8hY2Q9d0Dl5jQWoFVsmz2yJVhFZ5Amfh1Zu2SKd1akE
y5jAjPFmp+i8wqfDrHnTcjnGvmhsbkaQD6x9HyqzFY559ON+KW74hTzUJNRYQVsBLT13hPiiqkQz
zHJg1PnMYSgM2qlIbgOnXIFB/xkwZ3ipqpdMyLxu4hBQKB8H9QiMI//SFddZLSwQOJDVEeLUovsA
suAfPO5aSc1335CAg4VhQzRLqksDeEM6dtshvJwFLCrTu0+lSO///sY6SnB0ck3763tQuwK7Vu/j
8QBa78cSxw+k43/rKDcyHsW9pjjpk+DO5bmruRCD2j0nTCV1Uf4BFnVFQXSllx0fCQP//FazvP+/
y0qOR8ae6ao5XrTxiBBle2TFP3C8uTDT1dN5hr4AFzVGuUwqhvdUBFceltv8FY/fdT+79bhMKL+j
ji1LeKjPPs+WLiZ9X5EYSqmdqzkZ3SWkn6Kr3VwiPvHFV1N4FgV3NhoD2Tp4pK09BxJbEL+A+3d6
Rq5HB0WYg7pSF43xjKFHf6it+ji7OE4HCSa7t4EdAJx8oQSFpROaYG49BZ40NGd72FbeS70a/GOa
CH/JPZpHBCgezx4aB0GpOs5yrDgsfVljlRN9BZ+6gdkmxMHv1iD2RS41syfanr418PJNQwmXGLqW
OmCe9P1TFjtnufbFYF7LuugBAmMgutgIgjNzYgZIIQ4OpT5FOV/mOD+NQ7kHEfC4I4HKPY2Iwrue
HAuDyeDZC90eWxpkw6gCmt2MOQ/YnPVnArHE4Fpx5AO1uI1X1SPHES6BEB3uygD4h3yAZnjsjM8P
6bJgqjXRKRWnXxb5CgYzCVCDxIXIArSTGVJUmBOeeXVVgVv2Ix3jlawZFsJ9g5adURofiByjI5hD
T5vzyT/QZIYoVOLmm9Rz+8sFjbww3xy3P2htIeaqvSxvIS/+dA+9mEbanZLGMy4syGQcQQYvZJfn
MWHdZbXohR1Ps+lD0UD+U8Qyk9NeGUX/D87WeaA7Nfq+GV72QdEY5Cj1HxkMRajSqsxVdZvRE6hj
0/Hebr2HF8uKzdjTR+Thy2kKk21UyPqdi2fJBozmZ9IO4RJVXnuqnQZ1fb5cGci47qdZL2nGDlRH
fy3aRp5gd8JfQX1G8TwC14+Hf1fye8Qg1PYxUIBwbzsipYBVgJjXPMKxEt6BlkEAOepJHrZ3ilvv
3R+QaLLKdPLPkvYDHKCt1kHLpTZN7I8SWXr8WvZ/G3vzt7d7Irjv/Iz098KR9AEjA5qmw6o6tuQH
ALtyBVqY7A+EA6pJf2yr5G0UCw+XgnbyvlWQhrpzBl7bqMPb+rQecPr1j5bC06rHEAX3REDlJGXn
xLgVzzSn8FwdPGjcho06GmKAx7gkTtRlOkWTcXez2scIfynmu0IUyDPf+mJd1MrP6YPa/jlWOTHy
cegrsyqO8oysuySrpWt4xU0JryzLmcFC4p+makze54qk5soTG4tIHfnNjGFYD7NN7f9sNcvpCd8k
f1TrKxwxLoKHUaZPjiTbLbQeurIg+Lw7L1oHV72+ytq/8adijLknUyerjfOKo0mRkZYGaBgsTASC
yuPLPAcWS0Tjvi4Du+CLhEk7g0rM1FDqfKzQClLrML0Zg7lkA9RXfDvDVekLgEJAZk8KpHpUtQmb
q5pBn4xc6TMI5nPowEDlWtwBaKNjUa3XMK+4YXYgBUhcjI9zZMqVXgjxivEJkQ5frQ8uoiOOQe+j
eBtJGvPfuej8TtLV1ksagv14QMmtvfLU5ET/Rnm36jaw0Eo/Q2SgL+Qn1CJ4GYFT6nrZkxCezkSF
oE+4cvon/1YUZj1jz18rKlk5Z/daMTAbbDOkLZLWZqlFJLCS+RsxXiD7+N6zQ/kNBnRm87rTOk7e
tRNSWPIY6I99VMQ7CNT6X+MZn+wUPn5CfW4mne1h08KYvJv8OKh0EnZjXzSj2DuKtNfG30afhMsm
k3c/K7K0Cu6KaeKrzymJZWoZ5mSn69Gga6/lwWwHk6KYDziBsmmSydtyTHzfKaBiAxdoWuiqptNT
zMxUxtG2e3VdwBIEyltcU0z/jhdpPO4GF160H0+pxKvDj91XIwrQL3P8/3fX9p899vSIUSfm0Kxe
Zc6Zae81FcehQ1hhok9BJNNUZJ4h/G1OCj6bCvSfA7Y3noOT6A7uGJEnTL9bU0HUmybHGWqeGAzz
qntG4hGbMy00tUOQUe/r3ROsiF+9sY6RKP1K+5bYYMO4gB96lrJqgHPLItTcL9ByC08ZXivS3BzW
fjq57NwhKk3CObdfWq0vzkkagoSD+3Qp0MgH44h3F1bXeD0yPfx+kdsFxvd7uxemG3t1opibNvn/
2mqMaAOe9L15JQ/CQYHOhlxNzqaOCKqPYRNh0MlNaDfQfBKJF4jMhx9gNXftFMsvLHkqCDkj9kJ3
ITfHigPOZa1D0Ae8xvkv/Y0b3qTB2W9+nCfqqrKdAtRTOlFG+3cXtN7/4KVJ1BhLpiBsaM/YmUXU
P0JsR7iByxyA4T6y/3/6cl6MvAhBlgQS02f0HBj0co11yiOtIVmPDcK6ljjESw/NVdY02GEKXbPQ
D7Ic18vJUSDPOtxUU0UlqbE7eI4RtggmGXfogNVdKduWZSVpeiPai4QFUNs12lQRCWqox7AICRsh
PyGdAy3wdC0X4nTGM5XEVm1u3Ne6AEKz/Ta/Sfdz7bWFF/y/lwfU9YbxTLyjA6LIs9oZIxPUkuhU
QpYf4cvh4LJpQnEoc/z/TqK1gJcUqj2L7iMscGxayxM15F1N9RpCDlQsARhiO+E7Zn/TMzVC3653
OER+8GEdCAyUunfec81y/HTYjhj9IcamB8RXi7yPxtPm6q9Be46nJrtDrM01+7pU9bZHeISd2E/+
4FFpfM4wGoaPC/UaWsOAK8hLwHY91ocrr+oaQXp4KoAiDReD6GExf/2Ek2Ox4uo3qt0AhoM+kU1i
FmW/jdG8Rvd+xIbgcJXDUCCZ2OupuIW3+TVNEOrj0ULomAAnoUMQyRsUdC5WH6ZwnSH9pvRvaO9+
+GyaDjS1ehgX66abp67bHYogL1lJ5bOYkKTmg0dWOdMCt0HjpKxig3gAYMYhZfp/pXOL7JuHbYMT
xWWOTnLJ1YIXL5wR+qF05sxDwHTvpcoU5SfZDEIqS6795PrWqC4OKUeM+hEp3dVWHf6ZU1t3jqWw
XrJATnLkpYSaepuhKbSIorEKRqpIkYGJ2Cwto1J2PGm1urlGUUaMk5p5+V7u7nEK8EwEe2bqJcKO
AaWIhTZ41054CmUreXdiiBTK6oSEdsY4WLANWpedeBOImsGpkmCG97Novc2L+MjB1WQPj9dYL2XJ
ldpSciyM6CJEt0nHsrl78i1admk6O2ZDwixKc9wRmdzwf1L6b4WC94jRo8N7fPRpHJNyhrOSxJ/z
1z7yRZPCucuBgNkL1cLq45xsxDzJoM0wBIMe3IuRvwHH23z+eIVPGbCQyvZKr1WEgbmLfeN+6/A/
G4GN83Wn/niLFpjAX2LbCwiWdRL8708lDRH/PVUdJCXTzgBQ4z1ku7/D7J2kuwiw7hjxjihFmKj6
VJrPoAd5dQZAqRmchpNMhfqQ4AYLrZ82WUjoWj4WRyhXq3lEwJpQIbdGc761tJhplyIaWVa3dhyO
/K/msXyrT8tFWB6O6ssYDPM4OtfzGzeJbN3LWqkYffpg9i6CSvoxWGUMr+QJwKWxe0PFebCppMEV
BSzIsjH8arTNwo+YDmivUEQfCD9RTaXS2O8siw4opIJRo4ak6amQH8AAJv70wjjHSHpA+s9aqJ0m
gT7D8P7IQZHo1DYJUT6Y0M5r8YTk2RREhuf/Tkk0wC/9tUX4P8ha9l5TyUws5ZNBr+Mv3PyiYJ71
1ZKUpU9OZwl7D4sKKDXKjG+aFn1J0bkw6vedOigYGuIiKZy8E+GnRRJ7/p6adNd4GK0OXeCCwZ7s
o7HFeBAjAkqx5gpepvYMRo/RMGi6ASWtXSkFWwtv/qZ4By+URUD3SekVlZyzLWkvHs1YyY6IqUoD
p/sRZwZezzZkOwFIlthe/Q3YLoTFEvjtjfONyhpHg/XWY/7gPWE9kJinL+t66s+3+K+hGCfDehWt
LT8rD4csFLYOPGIUm7CVN3OpGlMkn5Xmk9TL6PyKjhWfIS+QRqp8knF/tHNqDYXVjeYHeWkOWDVw
lEbkV1YK4vYCOTs7u8ZReYqloB5BtbzgEgNEy0aVEXlsRQpAamHZUXvjw7cYttgE/Hv/4h67hmOx
cOKL8QZ2ArdvXqD70r8Xb8wvbMQdS4P4DgiKkhfCYgolG5CUngYcmJeDCvZYgFotMQnKDoWq7np9
MmiCPteyk+RXc9PS0dMofBH8mSG7ssEWLgoOB775wr/+1iBcQtgXIlus5867bBKsYdtehXT1lyD6
wi5yMlPtpAPxjKEF3I9GyGUCEgWyUFzjd7R5GpJzXrDB31GBwR6hgz5C6LMwSYbBsLhzbKEoQX/s
2/YEi3wVqE8kdtKU5N2bvPEiBds6wknVfAUsKJ4SwdXXhGEFMDNoxOHGb8Yk0tZA8JK2o4f12czg
8qSakJpEZN7e41lXckcsREC9AljoYkRNMPA1ffUIDkfgHINVgPthQnX7G8GRXmWv74hiA4MkCmbo
WrIwfZgT5QxHTbw8wkEhFujQbRcTBreN3ciCqqOHOkF3NBT7oQv0rs2/aVDn3ej9FLbelCOKQjGh
E9/NttFWfxGAmMSk2lRRu5HZcoA9aB+UtRqDLc6f0l3uMPDQ8g15+8RCHwo8aPWaT+2JhH7l4px+
peTTZudI2EILmte/0D4vQmOA7T9/Ep/6hVryGbfzfrzqwJQfIp2T/NVxYQJ7Okyyp7A6cpoZpZx1
kNSrarjFuP6TacL1ShWzAYhC8uOwUd3qegGbeezZs0NiH/EJoSJj9c+kOzjdBBmf5e0iTz0XBMIv
mZr3AmmccqWOc/ccbSLJyDG8xAeewa6cD6j6EQcBDuG0An31yBFLgDutzJCJiobi30qhr1KiwnoZ
YfSCAQPDpkSbziCFrwuMXQKKWqUqjc2P41ZGHNHrvrQf3oOZfBCqYFOhxzcLKJc6Bxo82p/B9k1z
L2fkzr3hAHlZT+yK3GAs6atGmKqKB7urEc2rb1Ha4yWZm8N/GhZIdZBpBU+MPvbjw4RdFpqT9g+9
G7JDEPoBztRW5Ro42JvmU2CfCTLFntCnFKS7yD6BxuCpSo059HtKXNkT58kopT81ASnPsMA2SF6v
JsC3YvzC3pN0plBH5Sd92OtCKIqjoNhHQDQvFn12++2xSDzRZcDCanjgDfP5uxZx1HNYaQEjUx46
8Ik8sOaQ4NIoCOXASepyvvD3EKOKr1IA2N4Xtgx9yvCQsY9V3QAW4jPXxpXIXNLXgN9k3d+x5cUG
6ImRVDW+X0g/cxF6LBUzNCJqG5ikYstDFtidtF7eClAXQJKT0904tt7eMBIB1d6Gf/UVn5PqrNER
tqdVCDzjzCsF1oEa34LrnVli4f5Pa6PkYFoN/vhW8HrWNQZuo8BCdwYNRFbuRv05BrB/Bu6caj5l
0ZuZGdcq6CAqyUYu+aJMrbgyPxaXvjW5y3jRt/CkJJjrsogKvvDB5Z5torKLxnUGhg9c05LRENE0
9ojJ67nd568Yj+CxY8J3578i0ZJlGQZ/w6UU/RBPrDCIf+5xbPMSIjFA9Jauj35Tj7XULntIaMpZ
FwJ8rtURZ8JD8HUpsyib2ayb+JwzV6Eo7ML+8hipbielszXFZwk8Q1BfrK476Ae7hvo9s+eU3h7I
s1Oz3Ourk6oxKjxbLKvSLEOS+o6BXPrkPaXMJlp5WffCokcelEfOBeAh26t5O76UUKwc+ngF6eyH
ApgCxnGuNO4AgXFZKXSw5nBBUA5GiAXH9QsEioFJO6Tuhra15n/3Gv3996xrujpoJmpqvup4dFU6
v6GWP59bdM7qscGiAepl5LZHSCtUO5P4Is8WCUKGk9vbtJP/Mjp8cmTIsWt33rAoKMUoNZAGNyve
iuNFvp+bcB/OzCzbbEMB1LrQGVHr/iiOXmg3DQPNFjMKw1lF0RGVpiymynVB4Sp7pr8vkzmfJFJY
y+p4t3FMtefKWy6QY2YkOSMTmg7stxY1Vn6BHaMRLE7rpsOX1X89Vcw8DYizwOk+1DBeo+M+qSz+
PglsGidcxsuBgM+oUs3ycqIS2oyHgjG1DK/mZF2cMj6mKvRsUAlXxUnFExjv5Fx/s7DLuGdQCyDQ
uH+vfyO3BeN0p+lTh9c2muyQ12yOh3MPF0R/F0oQbYJ5SLSSQibLvhuANZeY37pegeuGnsvUpdHs
uD2d4KzTPoFCf2MXkEa+VGxHi9AR94y3ImrBAsWi2sSNdrHvMRlurP+kU2C/eV9EHZTdoRYKjV3y
gvaUqg4oDiRo5jnDY4ek5o5VvVBLULtmpjlhPzXRMkshP/sQ5XyVIlz+ZrS5wD0PvHX0fL3f6nCC
BlHrVwC+DYhJ3uS5Vhl0rsG4cO700gcrO48zcTwAiNYAG4xDijff3rgHQDP4+MY7o+Ef+uJXioRZ
Ma0Mu6y/mMnmL88b97HTn0KCuSBLdmNrwSq75HUEuZAVcREot3R2SFWHxM4TpBvIcHYfIo3UcAs3
aQlCoNS0QlKxBdCAzSBhr1jS01bciiPFPvXC8nf4PJZ2DOMt1C8yWbgSit6MMpP7zKxch1EZhMwh
vrT5K7yaQxA4gV+LpI8wNJnp2iYMU5Hjoi3jxymaazHNmp2ZPfWSb0QqyXw6K2z0rbJIPKn7fhHy
F3bzgoct4p7vw7J7qLyesAzfDNMN6H7PtLuAd4J+Tefigi0nddOqifluMkKnS87tgklYnZ2RpCub
T9LTq5x9DIy7po79h9r79ni65Y/pVfKEZLWnrjPbvxooDcCEWKpdHke6fsdVBTMFawD1DBKUmU9q
plVk64cR2cfrWYlFfQxTNut9JPhjYRS/7zM+zIde3O2ONvRHPFbTk6fI3Pg3gBWBM2RcOMjTY63m
tR0HVU2yoKct8nYkFLiLPMZ7rKPeJSLu4tpqO1TOlcVyeATXSuYC7DI8wzj3BET2QTgdDYQLeJJC
E7eukVRIT0Wy/lWFKI4tniAbPch0amvxgQT6eKlKBYHKYpUt2TeFq36CKLjaJtLylwDR4Yv9Qfm8
pCAMPZV49d7ntihLwiMuFVT4HRoXrTOB+KA51ph+xubBIdSrOa262wlCQM4XwNgbEVpzYVF8PSsj
AOKgM1q+BMnjVfDMcq+Bws04r5bDCTd1zqaLJMtq+7RRPxOzDYP/sYNc5E6+wz7m/NGjtvdv6WPP
pyfQwi/zw52towDlABD+k2Bx1zWtKxz6vmN945s3/OZos1ulY6zv37In2zMbHF/S3BecnYLSXDn/
fljPsVvXZJm+ZG6g5VD2W2gp8cgxtdLZ4L9RWjUZGJddOeCwNQww2ayEy1hXSp5XUuF9rPvmxbGK
thiX6eMaecmg1FNR3snJ+hgDM0EXoqRxWUf+7jEAre6yeMAj84KQV6BAu7KsRPPR8zHpIZXhnuOX
NZxAkEiPhtLxzurFivNnw2KYhnEvZTv0jnSGoaaLrwJDx2U1Ebu2022NxjU/FMH9L1/LpZy69Ing
rbRzWx2tfTgJRm/20OG1M1Xvq+wLqicLcw3ASpyMHp6gSQd5bV1koKQuxcMaFNSpgJgvXHEZ/w0W
W0YI3z0fV5knLZofajmpZyvD2MSHKf0+YPvL/IiEfceVkIEhX28swxdE4Spgi4gkfTDTyw385j8N
TeTEK7TAfpNKsUJya3qz0VIMRz1xA5yjJmdEmKHmq7gHjpw6lqu3U12njJP4G/3bQ0EtMHKFlJ7J
HeHK9YF/wFLbJhJGRHTizFEI3pBIg/2k8qiTH/HFcvrfVRGY5J+F4lNiQl8EU0AG9MA4vqiHMex7
LbnhyUJgOWOYosUIEwse0b/Mh6fTe2xw+cE6Xbh0c0Zgr6+FGzW5wXPiGrh0smxAHNYE5ICO55XA
9UmAwYWk9ERYTMu9ixt1mwWidp4uUX48RBGJfR8ZHvXUQwMWy2u/WEVrRRqOfa7q6aToRRCyBpSw
DkZEHT1GD7gAGW26np8QT4+ulKXeljQjZCvLxXvAmT0/JuVvwybY9E7kUZrhCt2NJAzlJOSj6Ipn
fSgnceZ+9z0fSELVgllU2WC77W9E0WnnfV145IXqOqS4ZTcq4C1WG1FeCUePVH3bJWMQvpttc1Az
pThHCpLwe5pZ4eBRukHGgMmyY6qpU1kSHTf077aBP5+V/vUx4ewN3bKfVdLSdf3M2jjSk/TgMcAA
cvEF+P+gnJu8Vh8uh+XbAaUGl16G5Xo+K4BW88Ui+ZZQQUE0GY0bQpCpyqKzZzSL8xVN38FJQU3r
dH07j1aHzkXrS2y06GIzowFBQ5iSlN0JY8QnKSA+U94WCoLdttLbjVmLeW46H+ciJAM9A+KZ3k1X
+ZylBTlJQyrXFuUbgpWJlx5VBCXsnF7XG7z017AsLEiTyDoMzKlPgVCHeFo/hSsglWMCfALEVYy5
SdDZniGJCbS3hYXnrG7AP6NXwAmTXBMjNhKamAe7LhqWG1GK7eJpOn8hp1ZlyU0h6NrqID9V0wEL
/HAayW/OMujOmPN/EzZtl8S4IuzmNCUZi5rIay0gg0SyfG8CQk2B2l89V4daQFSuwC8ao56BvE4K
y7t0srJffdan1Giz6JLFKdGgFrBgSRayPw+04kDAO9UqZd4Cy4usYwNSyXKuOn927CJAd74l7Hza
R4UDwjYYz/+37eyFAtfokCND8AZSUyNobiQyeQ/5NeGA19cOBdUPBtsDAkR4gGAtU6uSuEXVX5oH
QJwa7+tl9mXwevXhL0/IZBvQjpUHHd9de+6IF000+pU4HAUx2zPBEofw3orS3l5kOBb3yXZHA7PN
b2IjcNdX99Abob+2rXZT81JJy8Vw2RNuAJ7hLF2+v3YNjtlfIHlivWvOJz/IwxX0HZc8jqib6Xl6
6K0omeTq/GD8Nim/rROwPRnYhDKA28s8oNhGvxe5sFd02VDbLr16S1y98qd6xf8tWrX7J9WXXIvo
q3+bfzRUKCFHhfnF4TqBhTznm2tpZM91fQ3NvJ5UZba2NkgkMvHfMp0CbXflJ6pOzQc1pj9Ja3jv
aJMxWvQrJ1gzcv77P0cUiz+0GpBOYkRmirkD3/n1LVfewlsJfZo50TLydRAqaEBvhf70auFFUgg7
wgJrCyKd97IPEQXZbS2iiaRdWTpbmDpzppmQXgJzm8+V54BWgwTtfGJZu9rQFNDVx77UUUUrBITf
VCq2lgnPUp0L6xWDgL54bvkSpYMPTUMZKeyjAdLpXzSLl6gFDk92vSHltOeM76CCcv7XpYARJxPh
JDDaZyOzRONU4TJIg9Tqqjb5g117BVDp88oesgqp4swI8uPzYq4m/HuR1CRa++Jm63LwVRFS8ZWJ
FJTPPUtRgbzMHtNNiHGFZ5uuctb12nAPSaVE1i7ceVn1mgjrrjvjmhyFw+tludMFZ+zwCAWUUrhk
DB3iyRgEDBRRXNIwIWnS/MnJVrTBJHMqaGn3l/sO+ayQnJ7WrYTZXlQcRlT/9EcKHQukr6qGf4Ha
HUXVeeXl5I0cQW9vi53OBT5nVSQy9/9y/h+IzcvNgTJEmRGrRC1mehf+kVXIKXi3deWoM6JXvcrw
U53GUjQC5bXhfURHa/9FVi/xRHCzbNcZ6a9A6OttO6J7bIO7y/x878ox6SehV01AP2GVvi8JHuen
iqeNwpXmZCrcKn5y8nrGdoNKKEtMr66ksk8VYdDFik7vmEw0uTm2XNhQPA9SZN2O3Wqowzs67+On
q80m8MptjiAtu7Zg2juR5dxjOd9+/ccz7C0NELai6GZMbIk62BY8fWIHOoH/H1ljhCHTuZfBWOZO
ReQvBjpcCacyFk4Pqvb9zvLVrGOjVpc9BrWeMP3+AlXhX+os1ZbKn1YbO2RQD79YrhJ7kS+YiU0g
oqEXniQX9XxLm5f4xnI54ZnRoWKmhSTCgudOIfneE+R7YxZG6u0ooOkJyI+KEd8iAb8OzwIbjIU3
eJIzql44uGOtcq0uCU/PT7VhSR7v7l0aUuL+zyVYcJQJCxyqZfNUHuW8+IBkG+97B8+Vl+GegR4F
gkeCxaSFswvO7HV4KpunYzsyZTL6IKZ9o6TGQl6CAdLt+B3mLpzj+odvSZSWPbJ3Bhq3NWHyrKkZ
RF/VmL/QjRgwwgGY9mqbMuc4BH5L9Wr6tavaM9XlqCiL9xY9GcerJKUPeGyZcrgqZth4jo4Sbzi3
QCbJ0CvE25vxUOuxu4a8uuNrUHK7MSdm/PsgZSnfMgvRZKnqP6xfI79j2XnIuZ1J8PjEnINfxnz9
OMBE8KRa9FrVj7qRromXmFvFF1PfX3DbDctDP2IdtHW1dJLHNbtSprckAi2NNAPoUHtCouw1ncDQ
zXNQ3m9cyQJrG1JL1GrI4q4VlGwMyZRp9DYS3s4UwxrB7G+rU2ivU/tbQQ0LmWHCWC7V+1yIRVn5
EDZGQGIyLfRgNEHUG3P5xd+rq2K18Ppt8QMDwv9POq/OYh083iB8yP9/IyMHVSedqyaZPSAfiyEl
hj6ey9Ol0FaM1aj+bGnCtWsG4EEJACpSsqbmSTc+OoOQjIxSE+tX/LaOm4EJpR2oBmFagsSs0y1S
AZDEuieQboLlVfa2V1S1ZdTx5P5XxcL8Xg0NsYk4MuSp6ZL4zoDq0S8X6A53cixbET4H0Pnu8QQ2
BoxsPstMAwXPQ8R8t4ge26XM+aXD+yctqVrwcuEVTgUK9MqHCXxHvXOaqwJ9xrX4ByRjWYN8E+y1
Eohg6J22+wUp97SHs1Fi8LmD9zb8xtRyVoEf9bDUCAUmvg8QGQLRwRAjkG8Z52PPEOmACoDAvotK
0vTA0NEw8dkfU2MXtWJE4NuqeHWk3GGeM8cKjUIfaFS5l2gAHsB5zBv4/AjBbMTFzrhLpKJTkbKY
tU48tlwdDpUEcCgHL1aD5htWqRUUMoWfqvfMYypexbYgToF7GTK9NPXcO1monMeA2r+2BpnAUNbj
wuFOoOGqIMWpAuAjfsWK1DAkkdrGKHlyUbVNe5sP7kuoon75rIEleFDksMvOoLSJvTUKwrBH95gK
Vy/gxKAN3rmOwPebSzPwT3wzJ7M5dQIFcD5USxrLuitbww7xuEbXc56I+MhSF+xXweb8OaQ6zRXn
GXI5o2bfaAcAlNR1cNFEQfhHoDwL/V+iLb5DNsFc5l4jiyLg3grDqTOxX0hLR4QY5bk2ZC4u064/
KstuFX6MT+DXTWaZ7VcInaFLGJvVp1M7755w33RNXRazTZd2TcddJiA8u02G3E59pGn2qtRmDRR6
8L/75423Q7awY03Xz3KgPbUhheh49qvY2VljkC+II0Sdf4SNwaJteKDgiXc+oB/pMrFHuEGeXC98
25wKWJEQ6sQVmATlTqGN8fYNDboCQqGynCxPBO+lGOJio/QywJD7ouB+A8V7jC6ikiNueF60V1ql
mkk81129cVzxEwzXY4Vg7JflO15ylgN9LED6b4uNKB9Qjxa7Kb21QRzlN37X7FxOHzOsSqrFRBA0
EMDnb2xYZTPkK1b5a941dUskNo+I/krFTy4OnIvUFwq5Wz9ja173iV7NZ4+N8nKaOHAkZ23yBTRl
AyLdZkIRV/qXbSU+u+MXpvIg8Pb8UmP6rcHnhhuq0P9xArAOB4ao7dtCyuur+1tVKNOTRwBv+5lr
lDj7MZFLSr8wPdFio7MjV7Bc0zNKifo72s/grEpyx2XFyrKBLrYpLn9hQ5340vZ1VkrMfYS1Aocp
7tZ8XlrQOQA6ve4pEV1rc/cSuhKDKFp5EIAOajqLRGLVqSlC6y/WDS+tqQwpCGP1xN51DoJ4jMOA
OPfKbkn4zWnDjbv3L57BA0RhTOYQBwpPj0gBIlV5ULHcXUVWIhBzV+qvBqgOpdInqvJ/8CS2mEBu
x24YcWCuVQtVzvq5MT8IyyrSFssgXg4341pjI4S1YDi4TFlGS9aj77zhYZ61ay2y5rjaWSpWMUrd
z50ADdCQfUd8UssM2hdgskQVTT7Ju3z9gDDmVglV1509Au7fQoqetXiFC7XeU725cc8gFUf/nK6w
gpDUW1irItVZzIjVhOoBPDkK5UCos+lS8KetO6ukKfNqfyNVUclXdRicjlzkPkXPsp3wObbTCZKW
5IhZx0Ge08fbXyTXip1TTJdAhG1ePAXEMKe0Q1XqR/4ABW/VYph5CUBEy6bShiJK/XGcJzEDNXUQ
2sOKnepAdjsxEG+kkeiG/dYyxpxEHzWNyuWOzRGCv++B/k1JM2dhOAIuNU48IxK/YEchTZs3EvmJ
XqYY2aE0VguptJbybHZ1TaDJm+QWLrvQm1xCKzM1oT1tF4E6F6cnOzsEiki3699yZmg6Q/18vSAd
rTsHpMOBx9GNHBwC6CXZmfwyB6/LnLn42CtDOz0EtP44ZuJnhInFWQyKC+La6ztW93YJQTd6/6mn
0j/L4FL1a7YzZuf/eU3/9Z34OZeTqM+ol7ddJ1yscL/exbCMzrKFZNHqjzjBuCfsOl68nUdB3qVC
q4ANToeECJ3oRchr7MrKYIfNhx58NSSgw/lhLNVQV1nVSl0Yp65LWe7iHn4a48lLlad/SCImn7qs
3lHsEfUnU6Cd9rUcrs11qmzHRVu8xTBY3L1Jme3ylCkNKAiuJFT/ycvelsjLYC4VWM4PpOdcnM8j
s72bE9r6MuZMTOd4AsO3ZpoD1ycogFPrauYS36PxivzhwgCDBu/K8rkNnawZ5KI4jSzZ+uUfbrcy
QjSifThT/ZhhB2M2sVpVFp7BqXV4suVoDJ+uMeFklWGhCkN816l50/42VuGxpAyeanr5ZH+jVjAN
QUA85qdAI3AlKs2YjGNiPBCJsmU0+TgiMxwAXmxwu09Ts8t87lDsvvS2tERy5O7ajOzB/Yl/8aOt
VdehixVnfIrW2/wcLXtBmuKhPu8nZcOWpAvV2kRQfV0LOjB5PjrxHYji4ljJu/5IYngXz3YVBqCs
RMIobDjROHtP+tombQysXNwR77RfbbOdNzECbJw6Ou3gsdDvb3ZKjcOI7qrdInV8Sc3L20f1cJtj
2MgaQy1Hg+q8+d0YgfKt5b+RQejvAXEypNtLn9HniJQwubaCLbrvm4/yow+8HRKmwek6EwdhWd3s
T2BiJidmWoFyKcdQhDPQmi3N1Z0SbaDbtjSiPkuO90Ij5+UjALVMUovG04MPfZOc/M0maQUKQ+1+
ZUfW83xX81tNV95ji/zdEEJIO/d6uS0rFSbSNtftMkcWDAGOpW/2++XO2jTVRRCu2BaUx4LnCWeb
vSi/1+OSg7flK5+tZsZtwmIrjViTXdgYAS+MmmEb93qSuf2wEYdNQfLLAgPcMzDNvimXGiIoEBfd
TFciSALNtHcfat4/STB2xflxVirs/itZ8hZBsO3gwNjBRQFac+ox5L7TeKx4de+0KVwEDT+iTyER
8Ez0Jf2vJzsEzUkOuaj8/N5MKh/IpMrRVxMiNlEezo+nKeKdMywDaAAv+2yh0Zua5AgWEADLxZ9k
T6wqEEEJ6TjokesZvUCRLZ3M7KeASlZy2xUhjl1gYRLsD2Gof9sOX7/+4HBegk/cMYmihQiFktx5
8fNpmjusCzP7ZT7Wlux8bPNi0BLQooWKtfa0AeH6/spZopR6humE6dr5jJMXBo0PB/IIFZJ+gULe
jPo08jBUOSC0iDdBRD5COoq1pmSss7aA0KnIuX+aSkVoe9a2NFlwCIZqKF/TfPUW5E5gQDY8euO4
MekCztILHRn3pckWmO2ns4aRWVQtB9O6t26jrR2KcCGdn7iIe6kGVOFvuwamue44sdMw3mPYAmD1
7fXrqcljW+2/qGPEg5x6Bo39wq+BmI/hT/7T8zso17pyUrrXWe7qUnYUCfabqSVJntdlgnP3HzMo
/1XOWMQ3S0MQsrfzd1VlftwBo/mkcDuXC8op3VhuMVYl2x4NlksHq/ThQ7varWHlayLSsC7fXfGJ
xtwJtX1iv7e/46xzCEllVieLS6YSkKS+PYq7rOyQzvoxYSAFdpWk1Jk15suL1R/dwu4xrKIvKWId
O5GBHArmBOFK1lLgEsv/hUa/n0EJZMBAs7TL6lhnN4eipkMoc03LOThDbZr/5m/DCSIUoI9TBLf1
J7p6g5Y+SxG/XHTuSjIrU5aNE7Ko1KEyabOKddnAcgKVG2XGAVuFsEYziPqCaKbHK3Q0BugUZFpi
NhQQsN3DWP1Qrwsg+GhTLsaE5TYomex2qlTI5gsOG9SMjcSoSWg8Vdfm7JL0SWojU0p/E+TTxuVf
B0sslmpWiGEY+vYj1x4LxVsRmWwiCM8GuSknL4f/F0Mhnr01DnNBl1Z+/9xzdDQ3fiW0TdtSNnH5
RFViKnkQSEw9EDIxlW3HvFxy9YH2QQ0pvi9gPUkJY4QciDn/p2zIw9Z5MpNfM3m+9iCDdHeif2G4
Vc+X8+NpM/xjg7P6GTxT+sMRJpA2qdQB2/NWADTapxU/m2fcif0LcKRyENdn95vkdu/YpoHa3+Lj
rw4ud5AzXHFfPUCWCxYDw+DGk3OsZCFnhvmkreeY64dDfqAsTFbpThqhWj6RfhG6tfgUGmIkNqfe
wd5Mm/5HTPR2DTdx+Ry1Evgz+JzdU3Y4H9BZ7e1NhsmhRuHsSCQd6djDAbG1/aAAUYJhsuTIQEwN
kqxghnh7eMr7i8wEWBgk7I65QfikDd0Ri8QYitEIjUTh0zBgdDcUBeGigY7+EbCgTE5fysOW6ung
trSVpf00xxJbjVWO02RO2kks82CqIJ19IU8O9FC6rKtkjTRJpjo63JUWoxZjx6pY0MBgFOmgarNC
xrYzW0b/ZuPiasKOFovvUwD64eiDSP3Kvc2ndh8JJaGbj+VLRuvmvWTpH8mM1GhYSGvjaA/09mrk
wrvf83gKgntVkN4VypcFk2HmkleGDQ9jFngO/vcvmjdFfFmqSjRlbMqZhV7UumqbkK+hw04I1MhR
PD0I1I1EcOkbeR1zOVlt5naA1yJA8ZnTSXJB2XWoCK2yIZS03zbCV82sXtR+kbmM85BZzQABEO0J
rk8/2uHrlIh34eXQhxMTXw2L43NHBBsk4e18jMoZmglBxW+Gmk2EesX6o2nM5AtgBdbVFi6FzN42
kPgJ3zHQkdfsHIspw6p07hbn/CPhxdPBuiqQJKxm36VM8EtZcS1DCJltPSCFnMmyxhXwXgdzCib6
beH6hoe1/r5TS4qnfsLHiPeMlb2Yp+Z8WxT/1gFwWt7o8Uo2jbNxbvCdUCpzfKNpvQyg274B14la
Ss4v4F6o65ZdsjObkkGOSt8R43h2mPTgkB0YNq9PcHPH2P0zI0vL6eQTgLCZOyEGm0c1+nURVEGE
XLL9THvMEDHSg0zpCEqbByd7ohYwlze95tlBVehMobzDO6eTt50nwiAbru4uJg0NuqhVvdjeLtpS
GJZW4MtOEsjXIrRRAmFz7K3NYEJFp5fM5B/aUDeqIpHGxQ5dkFSItz/lQ0l11VMb6NAeTo9d0/8x
7EEJPxdZu2zQE30MycC6VavSBQtJ6s1TKBmm+JeyxxBYbMm4gnOSZb6byTvBiPtkMvZjk7Jjc1F1
GNPH9Gru3nqlMvK3QKFV69xkF5Ll2DZMDr4ZYdTHSsuhwwX9l0asLYrTlzxu0h/VloS+fjokIN4P
L+3vTeZxWQqp0Vh1L2HmQiOi1AQrSvYxsH8tT+0+yJnvbdARva6gdZQKg0LPGUW7RpsRR3V4z4OK
+36B2WtA0k+r1XU1GYiv0K3SyycqqpwDShc/RXmKTJ4HaRdP1GBufJQAjebM8oD/SrHOhkss11Ix
qYHl72LFlmoT9YXHtcwAH8GpV1nT9B7w2ia7CyknDGZhIQ56ksyl2RGtO6JpySdcD/f6cR7NwR4/
E5MzSj3u/eA+nxcB0MAKiAboLIfbXff8RZ2aoN9RZ7rRcDjqeRmUFkt0+lGlVjJTBKzJQpdQ3Agf
Z2l0Dhrs2IhJKf1h6+yp4llbQKWoKdreVz5QxeGqgWxH/CkEn9jnWWAwhP/2L4BBH6celT2Iafvv
f8+vz5kf/iow27ewBcR/wLY0Yt6GYY6Prb1nSy8qGsJqA89YsEbUKj7ni73vEciwYs1ThexM3GJI
awCr5b2DQVIXiG9Zyb1wW4Ws8vZeLc8fTCA5La7IdcK+9A6/07ObM1l335G154bdc5vwM4A7EMaS
uikUtfEBaMs84EQiRNA0/OsojF0odIQJreuf209iZk6mZL9UIic1Ymg5pQiFvTPhIEVxm8S7sFTW
K+kmqAekDu+/+Y3uk460oLHBPMPmyDCw9gKdOE8sjQ2VJFfvYqMKet9u/EOkHl6TqJdmNUQHkvL5
yMo+l0Qf7PNuXaNNZpVciVssDdOq9kh6kZER2UEDIdWS2ay3l8zG5jfXv0xC3l8i16YMHp/vfw+B
QealN6xFfkb3smzoaEo/SFO5yeFFz7m/ui3yZoBm15NF22JSlCZ1Anj6FE4HAeDSvphUW5cck56b
Z+nIFunTxXckzfSCeYs/oUIzPl772ytIFqnmD3dfMi9PdNJeyz0fP/LvwCA9iBrEpl6BcAjL17x1
/SZ2lY4bMJYycyf0y0Ugi5wonckcOuJ+4amBCYv1SYyUpr8kRtKpVi+pPJ24ST/EuPDewQPeWGPc
sMR3ZRIvbpofYgNJ6CR3fgAFcIGpnOU+lfiwjadiY2q/8LUNXiDby/ZMR9mB7jA3+1VD2W+P30XJ
Je3DlUxGt9XuAqw13d1jBQO4DNdgRBpTjaAq5E7E3HxcNTBMkNgabIJnRU2KAgdvv2VCzOIt634K
qR+DDSDihE8AM+1n6fDgXGHyP5mgSkL8KVpYpUTx9+lePwMLgA4/46l9uYniu+rjURbyC8PYfqTS
OzUn2aDIDGh563uaHeDSJbSll5ZGDxNZAC6roOxTBzAxOCHwe3V6FQsuiwbL+DIpe/T+t+YVnO9z
CWJnHDfbLRN9c7Nr3mnuJBRBUkc9oZg4qnCaRj8QoXBwZjZK0V1lMyAPduCIpb2XlA5fPe+IZbFz
divkd/d55RGF0Mec+YJOmXQ90TgR6G0bWbzHEfpxQuc3ESERlAZ0f75ARxh4F2I3qcLF+X7NNF2B
+JMcpCdOfPbJnOUS645iG2Pbftgx8ww0gcEUgHkyZMTiHRTIvoG7o81JsIDn6IOG8I8znJi9D6Ay
wUjXF42hmXIaGwtd9NZJwMnxFgL/gJgx0lpsFnfdc0YAGHL9q8++NQGOZyqOs7oDpLqP73MkIZmM
k/Rx9lwA+C4/Qi1je3Wt7V32+7JS1tckfW5X2mH8FMFMo09BGGdpf3wC8OLVioxut5EiePeL2n62
gdiOnnUPVXAU1701tt+PIt8Dnq9//cqnHDSk384RvayAn22WgOzIgyg57a6BqddkRw2OcemQbO9a
qJYbPe8WS51Gm2L/5R7Ove0BFTpdrFMSwEAU8bBMSvksRW7LvFXaerlcwWZDlTPAV2l3XK6QshRW
89ZcVzK1DawSegg3TlSF+/ovQxYRCRkZ1AtTFLn4Q3FWXq8U5/i5GXF5DfobTrmAp3Gq7IY4T1tL
fHzg22O4hNyHqQbEUE/+S8xKczOW8feKl6fwPEN9Ure3R9S9dInF2SouHobvX+g18G+zV74gbFTA
f7kemA0t+B+tdSXDw1hFcIzRbYyGSc5XKTTm2Ocd9zPEVCTsyqIe0Ou7F+lf94fEwPwzUDpvz4pG
mmDf0gfuC2SSe7Q9gt40WdaY9Wqm4qgPRUjGRTDzT285IhdSr7CDc1tmxlHfyclpA+0GhdBnDZmp
DNtbMgHlYrD/AyaO5EmL09hSGbfzuJg/Hk2/3sNbtUOTbTzXpck7JMbGzCRMj4vfh/sFtPzNA3aD
INshvQPwSMjn1mrfBxqQS7fqriVZU4iVk60bHDvUedyGpieGNc1U/jLIMgPfw/qX/ZSA9dgIk03R
XM6R02XLZS7DDOXgUXNOl+JiQB0P/DGgkq5khtUoYRzW5S0NdExKT1XuHTvle8HKKGsJWgPcMBE7
4mZbMOUBlogB0OVN/s5yyeqsDUqdPg4O5mhORQ6Ypeyn+8Mvxv4UhtTBR2D3mtG4uybsQhQX7wqx
+VrNamC/Ic3j/rUKdqEgGDlseysQZB/x+kR6bXN4ieTCEI3Mu3ckTOuOIGf/Sv4SV5YHYFanwZB/
uM7TDjN7yssWHaVB0tbMUUG05SGx53Uki0IwDaDA1PM8vDwM92hWDEtWYEuaCW/D+wi3rzlrnzR0
J2QABeDNo5+FnE92frm+XtxWsLiPgq1tfa61R8G4ROTcNOdnITYPdk5XS9qM15VkzsuSpeKzZof2
kVVtj6J7EGDwxXDX8YK6S+6oD4635jpv4nLyoNPkp/t4yqbnyAF9tgj4lNd1yQT7igyiZfPa19te
pYx6LTFeMwkULhMW1LhyUa1V+Qkq0nAPdYhicYqchRy0fEzuEurJvLmivz0fTJWnJ1cVIWHwHfP7
axuY8n/wxAynOWkIBGy498lbIXBSLXJk0RmKVpzXKXOYGcH/Jgauz/V0mmXmXFCdWMOeIBho6w0O
AwOWhM88s+PnuHRM6+5CrILn8tdKUdZaXAknwxnw3yfmwyW9hANB+PqbdSt91UYzAmBvXKuxrqxX
OiygQNCcjaozHdCHZZS5Om4Wi6DPa5swWZgPDNmuHJBrmwBzk177oIeCW091AphbjyJ1LToIYaA5
c/WP8wi0SnAFs/ztndJEMaWCEZhGVxFiXUyfVDXHogdeHx5ojFrERiNO1EwY7ZIyYc6g5ooop/f4
VprwicjR6RpR2i1Cl58s1ZMgQgnW+P5hmtEOlO8TvKSqOcizICy5aVRn3+I1PC5eYk06n5qKKalu
q0624Q34VVLntF/9BXjt014iPDMLmqt6WLAORyYSe6+UUnEdJZiNEJdxHfaG/HYIg56MH9lIy0qV
hieNUiurMBjK+/PwPZPFhUgy0QqsEa+s/H5Vw16VZpBm9TpzzF1JTwsubTq/OTmDyfwbEkPdaB35
lQpv2Rlg2MQHyhYGN1HglVf2WU6ZqZlDyWsfSYCUqITi/Y6A3bm+fcF9tn2nu8p0P39VqXk7jrB6
0bjbjREkzN49i7Sm/wvryerp1wsNXmFqUt4Fa38aKd4qbagVRsDxkDm4Ij2KKT0FakpuYGUKdPWi
y8mCSfoT34/CV4sZPZ5HzuW8/p9GQxphW3O0Uy8q0bDZv5VlCzge57/qWTk7v027hdr3oF4Qqz57
X4MC+BecczLItmvj3aQJMoRk4kYY685zyhSEAYeT/4wqjz0GY+/sbCVMyWDi07h4oLzAuRlYXFij
ZHbks+maA3y6QQwsZS6p04GIVMFb+agSQ9RefVktRPDLSzfuwAul/eBeBcamO51vkLy7Ri9FGqT8
NWe1fKbJBxWufwaIIDeL1DSunMNURuj4meULDeI0R7Poqw3LXSPDS40twwy/xwdM53srCVw/+SvB
KOgO0EmIBaEox44px0CHHtvcCJyOoSKPlhTl/o3dAxNGkNllmZKEvDr3WSECQ93Vr/kvFtM54gWh
YFVIAVJDFAVlnTNVt8cD2ZT5TdiOBnWAqrwvx9+WtAp3t59UslzE6cmhWdbMk1+8F/LvKJam6fTQ
cWFZCDG9Gd9n9/mQVMcgySL5F571Vs73DOTpnhZGqxbDf9vo0Ac3mO01tbWx3/OmfigWgrZ0GiUV
36Y9u/EBuF+gnwOSvdkI3R/fZw32B0sYnwlkc+OaZDZxLSSkpBCngsH+5iz3uOW1ttR8tENamASG
URQw0bJc9f/tH6OdRbgIY9ER99B24ihov2QPKTMrMBxa4c0Z8UDBsNnPMpkPjoXiGgo4Lr4gwviC
mWM2y+wKj9BJL65b5MnFY8kTnKiZDhtIzVtQX+DNei9mkc9ksPw2cFc+Z1tZOupT/LgshJJ7PbQa
R432x7oK6OKziBcM513z79QCcECUGELYTb+TmaTQo1p5kzMzfT/7Ht9NOlHl9WM5TeO9cQ+Xh2ek
jtHDjGCaN236C20tq+bR+oVBcYbfle/EYo3/a0VegsQ7BTu4zMOUlRPf309c+wGteGaFCzlOgMzD
AX0seWXV+SuRpuGMJhYbGoDIPP7L+zO/XvPJp9wCvHPY3835kQDvI4jtHOynxtm4ayG4DgVwvbIC
TQNMi9q1nF1WQiuGCg8Xw9vV9r5ibe7lVZD0qRrB/Ji6rZrI4ikmb105gbmKDHUQ9xFBs6AvO1Dh
MSpghl7fW4CKJedbC9KJ824d//AaehC1/4ZESMz7HZGBVW2mJGxUoBDVwjkkT6T8UPI/eSzGX0QT
qbAA5MEPfWLy9AzZfuCFqmuNXvkSj9t8d3ayLKbTkti991YzbRnH+rnuHep/pnm4dT9Sf0mWLblx
PwnOOUM14loQF5ZPSB+kiS2LuXLsgwKOjQnPBUcSZM+MLcEnAv4y2IGWCVJfAlH6b33rbmPYQlae
alUTAqwvxedbGPZ7ZxenYSgCjEJ05DqNe19jaNvJm5sVSe6/UC26OhI9v9k7AJ70PaNWpIA2nVr0
SU9wLftYPbXLxfXdytyvvWzKJ4RJvxJy6NegLEpqfySaMxDM0lEHJPdyDY2mvvfIjlkaChYBgBmE
BkOcrxED3tBSKa89ryakvsoWmwKX4WVM499yXzv3JyNGj/no5dwxnZ64RU38r6z9vyFAKxrEQ65f
lHJmruN/06TnyQTUa8udHLwtk0DT9N1VNPU6Xs5ysY8SToFsxpaxRj1dcgnhm4s2BA1pk4uW0Jut
sJQiVBubI0mFIcA9kl7oC9GewexedZDbj7UBOZpUOTdzi7M5Gp6Mr+IZfVJs/Lrp4qbj8+Kf68Eg
C1ShWi3fZ2lluBQBeNTHK60l6UJc/4cR4eArRAKUIhf+JgS+4w2/g90VT1wKxRf3muGe0QsBYeRZ
OoqJoiafo4JKgT2OlyU6v0q2F3/CsNO4ih3dr6CYZPpV5frIXPuyZGqu7vRJ33IeVGlGAkDZ+EA1
qEy5H1wbnKlhDFFdKSPueDsGH4Gols+YZr+L0KjvMmmU3xnK1ShIXWDKkFRfeNvQ3ee+cFdkk/67
32RDANjDu865ARopNnYRu1Dfpa5HlW8SR0A8Ohb7TSrqWJ4tzQssa0MAmagMqrAvRf6+UgkGDlWg
PpT6oLoN7opFgrN+xJBl3kDNFxazc5kHXzCg2NpXEd8pdOQT5ofdgcL1nCvhSWLbuAJ9BbcmaT26
nj+kpY1bpapwF5IefO/LkNCUi6ZE4OqAg7MtXg/DRDP/SwkF+10BzlAv3oWBa8MDP/sYARto53bM
GDkHWQ0EjuaFzpHHsA3fcWb1KTbth1aNHijZ5Pkxsf6914GNUSwY2UVm8K/DBpeD9hIPCzYVmlpl
0W1hnodr1QXj1Q+jcFQJ/Q5Uyj9VR5lDgWCOwFGEI9oQK3Ctj/SyXxxF1nOH/WHqYU1dd8Qa4iYb
Lp/eE6i2ulmZwvST+gkbDmjDLnoFKBBXGhOgh2ENPCEnmAEKFU3aN7r61L/nwufFe+dy52OwrFff
nGtBTi9aesg1N3JmGej2TTQc9clWdjZnGCTAPlDpkxzzsmqBG2NeGjrABd5fEGFCJO8aYv68H0ze
d6IAFkhnDK8ezf+2jmKQ+zDg2CNBuu3Q84vdlUjcFSIh3bX6p58j290byNRMm3lqdKKMCHlfbvtU
RQvyz1qtX3kulNbjbTN8REEf4DAUV5EWaPZmEsUuFj2GsVyP2KrdFUiq7BdhPc6MY9AJpldxwiHG
rAoT6HPBfJF9QGUREQ9W+0XUcEVDx8EBp4HAhWtt3Oqjp2tQQp8F5xzdy+og09M2ftuR2kvP+Amq
+qPPot2VtWsGGREjXAcx3AC14XXm2qCqCebUVhVFgR9LHBbEJsQlqubHLJrN03rsa7eATawgoX5X
Hz+Eb9NZeudeJtvVCD9Qk5j0P6034sBzmCx9I7u3rTnyxQF1so8m74g3QKu3Bdly1CZJRl/f4s22
fOlVtoICDSvQvRiDfENH/045AHDnQcEkcTVS6p6kzXswlnPuQEGSX0M0AVzmB+mk+F6t/vbl8AQh
NCVEQMSN4Cyg95GXn9s8HBHeLYgoOD9eSU2X5LI3RIbTVyvVkAi2gHS8GWbmMWy8jEBIHuJ8C+4l
c/JEhct61+D7hkUfHX43XdxYex7A1LHDAMigSHPDZxYWHp8TIoQ7dJQ0IF6TebJeSJCavF34non+
NXlHKunPPqSUSdLDxOD5/EKeaNPb+KIv1jfgNyAWfDOTbdmcsVNn/HV5cbJJ/NOkls6Dos0Q7qeS
V0XGLKo7j5PLXndqO3fsh31FJgjDGnt61pFS22/qp7DL3cvg0zaowHlcdrh0AvLa74DOVi8uyE42
v1jKbJwDuZ01UTxsfkJcwZDG6Z+rOBWugJrH8bGDu6osc5eIleftcnRXKWm2xrVOX3GJxLrxHhFH
EyVQ1HZrpSXCbd/BYMzP8Eyub/xhcaoGEKbtg9FL3exV+ddos0GAVK729a/t8Pw0z5lyoEMVwCxW
fx8K3M2ADEnAzoWS4rK1lTcHH0ArG8E1RY3FrO3V1c6xG2GTARblKRQi074Qz/oWhD2b/o0mYQqT
+BG7DL+MUdhBeTNyDbr04KFPYwL5dBz5A3ZPbt5Uh1JocT3vesR8FfASiAMtYu613k3QQrhz5nxH
FsaYSo0TPQLrBKbWDl2acc1+tz7dcF5eeTFxKYOffj7XPtHPS+Xr7oRmCLx2puIij3kRrhA2rBHM
Hh4jkFuiAJL8FGv7woir9D+3EHFW0U0derVLmubnuDdvT7vROR3i5nRbdRvEBObOGk0SNEl2vk+X
inAWZuzZKMijLY63oHYVH28r4Od8hBMgv9NWwoDT1zVsfNdf89eNjBNm+FRCo8eZ0SnMnv+60Luc
QfZ0cooLfe2WhX8ua7TojsbFQv6dZpWW6CUx02O77uT8vKelYgpELANPpgI8yVOtYJyrT40rQ01Z
WgHNPGNKxGLFMmbh5AM4Doy/S3WrJnwXXLcfsClZ/r+LtqNsvM9jIoL32v0ICeCQXge/Y6oFSi2u
Rv2lMcCc84frbudBmQ0KMmvdszhxSDmaQe+yggo8h7IMmQM+RvUOqHDtGGTRbDPk+4QCGeqxUkW6
VdHrYcGfwEZqw0pU2/QtDfHkVR5R1O2nijXn1HRBvGdpllopvT6eqT5tGsquKzGtKX6fZSIA6BFL
g+nJ3JDPNfKFwdJxIP7ihvRXBigXdPScFcwXulISM2zlE8ojxqTGPT5ikz0Hwq+tjuy1hPT6kfjG
T6fMZ7UkA3mkxLho+P+eHUbw4Iq9Vbkxw6p9eBNHSFJyamLbRn6x8eKhKOKg00C6/6gm1rjT4KB4
o6DqhXUEi+oA+atb0aW9W/3bykZC/jLQRCv7LAVSQWzwgddTNeucqeVRkKzN31hQLba6/3YCig/J
UcLvQlbK04HFVBMj0C/OW6enF/x26tty5badeYAnj0wjw44hsptXrW3NRTQOiNVJtGDPr0S2QDe/
AxaKy9MiX3dbf/JmEyMCfo+97jrIVXYEg+GI5PdxU1OHGTGl/r6gJeRBvFBHiGQGH+c7Z4bkHhHu
F6u8LJOTd2LgacLPA6AKPuyPreocdt11KZTF4NdNHVRhzaDkRtJLsiq4W1hyF1h7L5KJxgh3D1wI
Hbfp7Oxv7l4/iBocFhrhU+SQ6xUnGmR/f9K+sgLvQHNyXLMRPnE0FTxTkxGzutvfedbzhl8gcLcX
6N4APWoKy6zfOGWFMKBPWpbwxwZS5xBBZTuyj8qiSg7KaIrnEeyJE6U/hEb+M5H2VLTqO9naPU5Q
+rP0CcmyEJhT0pvzRikxsUM3FzCy+gQojuf+fUxzzDFL3HFU0vJbF+qxw9iOH2u2z4e4wfxUgrF0
rIrU9FVAvUSRWOExvZI2lt2vFS+qbzrZdIG9Xu1LkOxA/IXRUoK2IqPB+P4piDZaaQtFDZ3abvRn
HRo9m+o3FJUgE3WaxXpMMm74YEQOOkfaKE5PWtIZ/CpjSxNUh1ddW97m1jUkWB7cBLWga+cWLSAC
Kw796yDxd0qFjGdJFg9Ct9ERKcRm27Mf2VAyqfYPZXohKxuVym6uBBa7tLNVYPZn87A+MJeA+SfI
rW7BEMLr83YKHBhnDPZwXwIa2MFwYdiKeLeUiW8pSz92GYzYIXlpb+HLu9J/j6vGecyNHFhZfl4a
UQLDD67m4JcvBj4aFKgSqxFxOpO65TCmDdIikahg+twkMCDv1I6wF+OZr5uGGzGPtiN/qgASibhS
8M80jEoEOhBd7owdPl7BW6VkIj8P3wU4EacsOG2qpcZ26zXzihrhSHS7elWLOXO4NV1pCjTSA8Mh
klZ+SGpdyFkzSZJowjd0QAjWotyeCIVdhBOzMsH59PXUi73/MV7AaFZeeH23J2VY6HHRuZ3vJXLP
bp/F0i8I578C7dh5H0Dq2PFW+WZP6ZMO3QwwogvXEzZ5O9DlUzyLvlm9KoexUOyY/9fI6T+GK4ZQ
YmwgAEAboH8JHesKBAgRtc4LUn0zgvJFJvofrVt3USiRD0cg71Uh1uVzqyYkcQX80fZ9EaOrymuf
ZH1H2/oKsSZMObLGO2UNAQduPZ9l6oBLBs2ePm47/xZ0/LfZh43wTU9wfa+VXb1jkXEQRwVw27Ho
vMm07pO5Wx1xjanPp/3AURFYnfvtxV4syKU/7PA+ph2zZj1LbAk2jq6I6kJCn/JGMjRel3NM7Wdu
8H1pTfkwOUAKILBI7oaRoQKnt5hgdbMCtQoUBCpw7v4HmEZ1Qq4Y87/8IY4fMn8LF/RyAXKOywpU
u03R5L1LIHVHVI9W2leufUm3J+o4ndaOlC4gCpSmAAQqSUYgHpHUw2LjHHf4aVQ77HzkxFSk9e7s
OoJ5fC2JR6GqRNux8DZkruGIkDIc+KXLPBcZEfTGI4eHVPvv7SsTHoH7FP1CtBkGPDchrh71gNGG
kxRa36bBQRvJtz/bexBc7H1Jslu1137OyPRIqTDsyNCjm7KhTWNZNhX/dWr0kQ6n6/l8Er+m/ImO
0uUkdUxpBc/Nzyn/X9CgWVClBCjQFbGp/RZxwpJ99s7UCHS7cEH5nKHghqr7vdOZpVTgH9QD4dKT
jt5L6/k2kSjovuUgOgWvAeMcDlvaHjZmd4CvCXByN71zwjInTToiNQ4nz9TVBBmtjpj9osKvwiPI
u0frbY2aOEd2B9OmReJEc5x8esW8IJ04xJPiY8dNLYw9Uvz2dKi92QIb7b10ygHk0N0RCX3Qtkq0
5Sa9Pdrft7L89p2WN9nQoknBPSaSwXwc1swEQsgS9sRiT2QQcO/kNaz9l5G4F+22jG4/kgIXLfn6
J8B+8UTLFKuuyPPq6AoEYMRJgUKU3xzyuhdwwnAnWDpCHFU9+sUX4cOacHqAw9qCIviBEERztvBY
WxJ7M31kbZBqpQLSknaOWpEZTbsGuehkMyipMo3Xz1DwUBsn9Dcb9zfk3ySdLbL/Z3lTZVBhFRLR
In/zebj+qqntkJTTyvYalNPhiewE5ktYeytEN848BU+Fr5+szJJQQCjcLHLZ6FTL3Ni6gk9lG74K
ih6tQvkW1NuKOiaQfBGZCyZXS0GV6mjSkmUyT+4vDsPR4y0RM5CeljPTFiwYxWabIJe5gGrkhX5N
OcQmXAQ3PEPLAINjHMBEiLmqec1lnil4clNVaj24gQr+YFQFL27M/xqegxqAIRzZv2yY3I/fx46B
udkZfSX3sWChPvUD8bOPude67OFvnY3YYgOt5HrOhFWPPJnCNB4ToyIPH+K9sNQvsRenCNSbLIc4
lo62EUp+ryYYM+b3VMD9bx1VEeWNRsEDT1eJHJqwQLYN3nqVeXf0kEoI1JFHiiB/ZjBFN+6jubUp
YiC1dmh14BS37E4DpI9F4NTQPSHcC8L1nxtUzEWQSOyEZqp9ERsKeXVbgis17hLrVu12hNI0mJcn
BSDYWFg62KyNONgoO0Va1ln+znaJFRSJMuJa2YHybevnxtnefxexgka6cYvLY6gI2tJx9n931QqF
aP8VJ4IgVX5p/kPQcF8GZNsPb696Ur9h5Yv0D98hpKiKx0jYbh7akhJrxsv1w7mw35CtDG23nGYR
5DcDkP0VQWlEjOXjXgXo00G/ibD/6q3VfSJG8YW4+XBGrSVqWZlMPvzjkuLwFxzQIrw9KttYNrnz
ZodICODfI1Fpkfg4hc8qnmG0g8mD4jjtxXjtigAgMtIqdR0SINlyC7jqe4x0It68SxI9Xv7q28NR
MTd6NkisC6niKu6nY9h0pQSTgW1rMAZlRpP8T9lriWnKwToLmLE+xp0kVD9zMW9MIJfZIK+R9ELD
pX2Zi3BHO24vMdhnNTF7v0rQ4DkA11/IOC3bWL1ZKF8W7NVbk5fIB9BBBAdXnU4chka1gTLU6I9t
goF9evrHwjHvnL8qSA/s8DgAuAs+gR9L6w3wIqC+OQ2S/7wJZMdxQvvoJ0o2wMCFe3EwCR0nYhj8
f2BywyUkQsFMc+0MN5YElHmfueri1YhJI7NvmF/xvAkfcbAuIAiUJEHQxxlc3F38tzqGNdSK3Z9g
KCz9xFuTO0CD68aNoPUxAsCjiYAob1yBvuoKjIeOZ/pJCxNYFAJ/6YWYVkvbmS9fCbbL6b/JsPy7
W9QJ1M61oRoG12si6k1dgVcMI/FeavzzuKkvlHgGuRjIOUTjgBK4gcxIkJ9c0zcPDsoTjBgFS0S2
xMN07ggi9wfNeZmjGO/DERQRYVk1dmzEUUrES7lc4JxXdrOcdsMuCwRdpRV6iBE0S3N+gNTgObwn
Faj3APqIy//ijUy8mFfdVd8aQzZ+7S4CrJdpKEqwBLsfqdS28YpKaMo8wvAzYvjEVpwNoCOE/oiK
T1gFtPEObdeugxRUmfwNe2hlP4sURS+TwWBhuMmeZwxUUvGUhizlQvHEgIlUosa66rdHEGi3lIoN
f+XGHv+EXUn+h6xk3udHEvjnPeiXkTMgSSP2evPdVBleDz3e1SBOa4xwfO3lyA64/9mCVPOqbezV
qvlXMjSPYShcmS2OsowHnLWFfl3cNTyz6y7ShUR5MPs19fEFYa0wk+mq2YDhAZGmgWlK4u/bpof6
Ds+ZCxvA2g5Thc4yKNbqTL3/FA8zIFTh7lMxSKSPf7+d5Hla5X5sMpza0toHojVf1x29lYXMKmKk
ALzqMB4twkwX767Bd3yTb91TvMlj0PwKBHrwt1aDTKZpX/aFgibxtmlgAFcX0T8kQB2hkfXDbh9O
anBvFhDrt7o+/Wjxl+eDp1l6LOtHSg5K5uksMddTx9fEE87r/uZJrOXlLDzmW0V1QSPc0MhyKXrW
IaSrcNLF8Kexo21yP2OTgo05Y/lfNAIossEs9eS6SdSIqgp7jgiz6kFhlZFr2bFiJRI9VKwUMIMp
z0W1sufn7v1WCTyiMXE4c1Y7EcTplYcrhDTl3p10WlyrrsCpc0U59t1KTaHbernBc01CWBaMUKkV
l/f2kOz984QJOSKp7Natb0x25v6WpVJK9GN49ukoTwynvLupTi/zK4D9tGH97fzqZLf195XPxiiA
2StSqs/LfWWd2dQZiJbqnI8P+DyKOyCTL0FXd5Y1xwaVESL1YQeHDNJIdoWRGTVXARxvyPtnYEwR
2UFiKrmcWPtz5yHF2bRXszKUIlF+g1FhBZRIu7WwkDXG+DFteOrFvgC0aaWZ88NMtOXBMMpZDpLP
SunhepjhLAkw08S2hDdGIGS0mAKqpwRITz3JgFLCwxVpVpXbAeqLLT9eUN+zKyNfga6mdYMAlfXs
SmAQzlkkvat59nBfAFKrKtUfvjnZZo/MDO2g1qKH8YA2U/qozTx5MgFsqu/2zkHoQDycX83kTjdo
6LIScA7+zRlRi/xuUhDM8b17b15X+2cgzxZeN4JlatoDEtaC4W0vLbvozL8Zt/5B2G+ChRQ1tnXm
iU95PMqptsJdUoydsSNLxXpNj4drW0B88ui2h4cnclV/1aUIQM0KWhxWRMnewtZi/yLWvIidMWQK
dEw3KGoWtLEidTL8Wo8my9zUaee/paCas0wexv0g1DWOTMAzCOC4kEnGENbRjq0qTDX//kwihGVP
CaZXfywVAzcMtfeo9Q/OKllmT2yLXrQnrm1woFQoT2eFpZWV7TsC730RNXgqT+2JxO9wat7BV501
GSrZIEru426LOeeVsnIjW/4dlfQ/WmsJkm43OYb5SevwVT4KZ2N6iPHOXStgDs0H3MadLphMakEV
wyJLbNvicknLKnDgD7BjUMAu+S2kgOSY9VRjSyV3D19v9has4uJctZy5BaQDQgUy8T+Pe09iZ4gF
+06D5Cx1wJ/SeQH/zIYD3MB+Obh7+Okyyf8XuU5OEdlPmVdmhqHU5BywT8CSF0knSJkMycxc2tDD
RtwxyazqAwu2Bel6UQIuHjMROGYTd/ikPG8VoMV3yz4I8XlEzcuBmLNmD4YsaoUqiKiN7qwFucNz
rel0x5RmVu60TF+cfBjhPDQhc7ySRpXPVPIXdHCGM773uT/NEkh9HaMh3/jOqWNk6/VW1ipkpB3Q
mMSnQgJ6JF/73kGpOWN6UXUA9wi7TDNT519eYWyu1EAFO2Ws+gdedLqcTxuEBZYj0ULfkwMOi+XZ
RZyZRiPAtcnjKU5pPELumamYBJcRbPb9jkNbKHNQQCe0qflqMOSCAejLiXOyhKhbFG/SI5m455ge
EwkGEU7Q2un78TjWM0rnKNQYEuXUJQ13nrk/DU7WYAzyHQGCzZMzQmhbq5esLLiIhDOkMJn2loas
b7YrGGxvv44w2fYQzLljGQz2GifQUOejRBRgchaJ2otGmz53uwxU/LdJzyJa6FoVvf0nIduNJ37c
ZnIvgPQ5rwqJtn/5qa8izoycatneuDgws1SI7n99QmY+5hKPWvZj0EhgL5wa/YBL0tRosyd46pxZ
8o8fOQ0VHwOh0sYKmdwfkdptmPxI276s+aAT3QU7wYBw0Qd0ScRPiX9KzVEY7iyetzjlTknqoto0
XJzTVPTHFuo4qFshEvKrxjk5K6M1IRz7yHEZaqJc2F+UiegW190M/9m7U1MMR1Mr4IkLIS7jk2k0
L2F4lsOE4JRFLoSl/2SM+jRMWaeUi/owfmXnTr+ekZ0iHW6wZ+2cNv9C0LY+wfjHxd3fbjae+17+
L2Zlu9P1vadI8Wv8XuHXA4Xl25Bixgffg5wdanZiTHRvkdI1gYxS9/CVxhylPP+OB0t87vnt45CX
aG1BIboPSwhbOBsSdeweUR7UYtH7DZR3cDYV5KD0F9uBbK+s2worthCYE16gEUhDGd/81T7bVzmX
upyguGZYqVS26DYlt3NsHT+7x12S0yo9uXBJ7iP/QG5jlT188qHNysO4N56IOC3NR0KKhK76jvHA
ThXtgv7sjEi9aGIKv3a2xm7yt1qgNRNyhLYIWYPW6Q69VExx66DzqmYmmICzwxPDsOz9Oy3xfslW
LGxeRagSkeeCJ+4AVymMTzOb7r3ZZWc1DGcVG0XGEWZLQE1ZG6dwsJfMbKSSI9w24I4TuIm8CIsa
f3BmrXI2uWhbOFCwv/q9UHX/3O1NNVzxg/HuwuvYk3xDOo7P/z8l73TJnk0NLjT8rouWwozpiiCe
UJvCoJqgICcQfuLVWfd7BCaSPlg6sz5su1l6IAtCpzchpcpYibPRsNnZrqgpVsZ9WyM3j6PBwmSM
MtHKJ4F5Trc667tMDmnzEo+9CevR0cFEUE2zN+98il6mf6eWBuEVqtqPUMu6Lv0Hx2YVSDNMakwi
gpWHb1jQNzw8f8dflnISdK13neLCgtGd1Fw3BthhSIooh5XGxarSR2r8C1p3c+aeYWw5H4FD2LYW
UM0K/x/R9gVseU0W1kOOesjlkuSPjyMh1+uVj7INf4uTv+ylyPT5DJGNXLUn8W+Hy7Sxv12wXQ9J
epChOO7WO+QWjVSScfuWuOAzP8IiYAPrfCUbamd+/+q8t2TcJjcKKfpfEoPAgU43CIj06fFOBSHz
5UvZmfg+xi319ioO6UdFpYsYzwCvM5gwlMOG6XuC7eWO2VBP69VOuo6clV/Rn2yzBI+ndVb4mMMp
cN4mdpnG5Xfysqy4ogREgQ/VhIcg9qx3gzeeN/DX9bmIpou4ouSlOwqlX6XT3ZTlrkkD2QJpqDJ9
cFbjK9nhWUThRcdDqpfI+Oq8TKeovZSrK4vj0jxsHNNbMVVeA2hcBpTHfEDn3mFwslgSuLQ1TFGU
T1BVrnUVN7SCjts5q1F5Wjmi+nExKMxnrtuYhMjUyBW4uMe52b1Bs6yzlpI1vyScGMb4Vee4rkUh
numc2WCaUe3vInYC9jsB1NarS1tB1YE9RRthsX7dVIAbR0pXLy6GtAgRVlow/oZ0FXag+NRTKp88
pzPv5Sr+ylfRXvj+46xDVm/QmBBu75U4UQe77HNjMi3wd6EmEGvZ6NYRrc3uLJkEHGBS4UpZ8jIq
xwZiO0IOfpJmH9fxQEHhy51YC4GdO9n2oPnABbinp+tIYUmAczfDSisaBTBmtwbINE6K6g6i9Rld
gOWyVd7dCbIPJo1lIH8Jx6oIcWQhCSz+fmYU9EIvSgm9qf+/0dTpysIJQuQuPYo9dqZL6vnCG60F
vEnPfygxt1FT2x+W+lVprHOZb1zjMyFVOnqf7IDM/XsoCLqHJzCGuvCvNtmD3m7X75Lr+Fkp3BOI
KtBfA22Md6N1izTa/luSRkK/x0c/xsx0nDEO+yG6kQ5G+dcEMku1tAlqkW8ZFA4Nk9fvwwIidJJ1
NOF1U+cbAtkQ9DbqTa6ogTVh9O9I2rzOYebwmfVsT/9CKcqWplq0vxxJI/PXdVjoHDHdwZtvnrkf
o4oKGZGzB0mI61NxmJd5yH/IKSj5n5YZodZnopojHy1syv7/JCBpbM7idNmyXxy+MB8E+bXmvTmE
UgkkQET+nowZ47DTECegQ9u2xl7UggHQixO3q8YH4DDhkR9dgWLSSnqkopVuBdhJERpnPqmDs2O3
4+k6APThs/k0wzM8Jcxyx5ITJn8EU0g1b4nNB8lIZQ4MCroO3At1Y/nUJwb0YEPWY7pysv5oTZHi
42uqt7ohb+BBsgSKlukDggIYjH1NqvUM+TGo/nyHjZhbrAbYDMqnIZU6C7mkEvGY20tg/Hyfw51x
kYRqbOdLIkK0uvfX700UGAEveReq9zijF86NSEPtbHkkneg/1b8dCWb2TdWRNYmQKfxqSVXQvQ1R
goVdKt5TUnIoFrg28yivegEXkUTZiOLQjZ/7BtFbxs/8N70ycRnpdjwR3Aa0bpBB0oHhJhTWXe4Q
LfE/W7QBsjJ7tD9P3N+vgXxHopqFQk9ilI7ogBhcZVRpwbO/VrTzVDzGzL7dpe7DASLMR2jgUvUt
X7t0HnjTchUwWMjhqf7D29jnX0JP35xaMQIQSWlu8hPvsQ0yz9a0vNrX8N4j1si2CtVGDCawTWsN
5UEwSwpx9IiWyBHWuXfCCTle2Wtp9WW0NAEG5X2qiS53jL7Q8bfK4/V8zI9xXUjk1eKouj/tNNi0
6FkrYAph6F2qE+Vansd4ru7Tn9HhlWaCbCKGFfQshIcXE7fGEMN7aqvE1bvxzYN4PdBSOt4rhNfu
Gi/TxBuQfJa9+Y4oxryTigkMEam8n89y6ye5D+Lq9wXu2fN79uWiGTydw/aRDom0+ExzNKwQfcih
zJ1px9cFt4UFzcfS4236Bcv0joG3HEDstCcrml4eN6hz4/4+4PsNnJKDpmbUb4+rXQ7gspGC229/
TMMCCt2F7pvHl3e73bl3JacPgk8tOZMXFvKTjy7Pxt/rtYJinf8I+8GECeNYwRz/oK8z0kr8yNxb
LRkIfmafnXuu3NrjTSsCkeqNDJBWEPIJrXh0eonXYnyti7AZBFzRuh6542Pa+Wom5GTk/T2qzA8p
jzUagqRQ4YhuW+8wj5Ohtv6DzF8hD+MWJP2lTqw6F3JMOjUn1VrdcTE8P/LhLDrrYTiinTmBfe5L
uhA4Tg+Pt9c88X6stQgmeDSguK9bkG9ubESFXYmBgfLf2W+WY7W4OdWTZsfolu1VmAVDBPOFYC2Y
k38br+wKEt8xnwwh6pUfQtUgeWS2r7oNP/MhPyMCHG4+pkMTOAmTd7+Qg/OanTvp/lM2Ckguhw9E
FJGQdAaSAIvhU/M8flrW47MdyrizdBkn6KHUmcPenKxKHOxgBrADrhHwAjfQjpE6pm8M7+XEn+MU
gjxVkqWCNKChCyqxvBg31umNKwgXrrJr9trILrT7wbPTp/thO2sm6NJ13XmIkHtQc0sm2j4qxXfW
uds6xSLDa3eS57X493i5DR9pNne01ed+lidBCaPJjTnywmdTvXQp9vPAmG1j5pb3Q9vuO3UCD3lz
8eIRS34Ci1QR7X5DosyRRM00jlzJZouv2ar9u0vDkiA47qMt4wAKPOTXJDNYI+zCgaVXy1FojfZ+
LLaUkllcm2mbM54Ue7l+JhOuDqbK/N4JTVGrVgKepq+6VroVMRqbweUCKrgCyG0Mt2v7PLo+Tefs
O+dHcJgTb4DHcXxstIi1l6Pf59/P3xlwHFBxYr1dvudXefdiDD3lddDsf18NPCv2oNIWCr2cuOoT
ePZaB5mdvNr0kLrL6avO0Fy+NsdxtCNt/REJMsLmKrcgFh9iGKFFgk4q3sVa7XsV7HXSxfigec40
mD13HFrztX4gMt3NwlukalDWwR21NWwmue1hkNvN+LvYgKmEYzglxjCrUr9pDUtQh3xIFPKVEPn+
Gx+Z+QTJzFJJ60Xo2ZIMgV6+iqfqTEKF/d+0NYFLPfQn6lOd158/Dv8tlIMu0+2H7+gCxAUrw/oS
ViFTZUYX04X3q+vu4W86lOaN687A9hbjNDgksQFSLczJXuXrjzerzUWwshPLbKOlP67QjyElUX1D
N58bVfE8uObhja2J1LY9sncYXFcHf3T1BvH930Ku54LvjKtQ4mVPq0MBloFeACR8tShzEVfPSq2S
q1MdsXvGgdtrrX/mlKHJ26KKEjnCRLFtO9d2svBFkczJVvbvs//iSLDtAoPcXQbLIzFuDx+O3Gtl
priD+1BZ2mslbTz49VlWmZR/vkJgXFL+HZqK3LXTcPakOjITxTM81CtbNH+fmeQf2UvqhW/I+GPh
OSV/PoOLQHZMz09yCtoEOMOEZNJozbPN37XmdOABMTUz4OQnrMkJ9j36x7kib8mOF/wY8Y8Ylsay
VqBkAkDltOdqGzyeCi/9MgFYwVjLK+Cw2S1vo3IE5Tf6iE6BQJXqaNHhaB7jkq3PtDBeoKX09cbE
R9l/jqxk8P1X21AYjpLQBa2lWklFjldjgLNyoCirV0B75BHtNT2gLbspDd/RfB7r3rTHkfvcD1Iu
bK+QwJ+WTL4H6OUgyyaU3jQvXYVRYlpTkDCtCKd832eGhx0yer5LsjJcthqIu0KJ5kvWoA2rn019
yn9eGbRRfDKhuPPTkqOi1fukK/co6TfItNDWjil9530081UO863o3uz4bjZjJK6riFuN5emw5U/R
KRppuxfXjjJBN6JAQoxGMMcHUVMJ8sepV6G1UDNUenRcUYhGLHrQK+qE2zzc000wpm77BpskMU9o
QI6oAjAd3Lptx0wCKdV8+IEoTlKv1kiHNFsSFdtisJmxGwHB97CskU9zt0HqlW3b1vRs47Dh5E80
wAHvzKIe2BVcoeF2I1OvmJQ46Oy1QrMzPdEYGeUSl1HOKvSB+iUEeaJawRs/3Usil8vy2fWl3oNt
0ETag4xsoFkF09i0kfVqtZB2Y4RgkCdX/T9GbLLEfJ6Mqn+NSC0guP2Fqn5bfpK34YUFxCISDj/3
M4Y28vb1gpokqdKLtJiq3ckp4mUZZoTQlinB6LK/yG6phCS7aluxAuz9M5Qv81Z2zivSGa9pFZ6E
NZHlP0iZIQod9ZuNOqJ3KFI3XC2a4jDRUX6klkqyyYXIbbZPvVgusHf2CIQ8ALSLMPlNcY7Rn0CN
j51ad5FdQd5FZGPBYXjlQa98g3r4zaMwg7NxKVi2pjDPPfW3H6sU0eISB6tAnWDp2dwjksnqIQL8
yYUOdKBD0JPgqFkdwBhL6fir+omjPeVGTLTTVIXR9T20gYxUp1pv6MU+8OJy+BQXX3/RkwqT4JUc
xy8Qyw+vyNjhIhqeFxIrUGLiGa4krvGjK1XDvMAgAepoZOWxzh9rAxoKYuFEfTv9WHajQy2lf4/4
QNzcv7yAB7J4ZbaCeRG6QSSZqNAEZLfd8W46r06mGFlj/WWqyqwVwxheqAGkaI40qp1A/NPsyOo/
IrJDsVODXDwpICp0zS+Zz/SUcUZXnLd+VGP+h3GkEFkKp7QkcterCC9av7+3PHT3+EZ7gutVex7j
WpwjExGH6QQarBy4qVHJ1Pjy35yHBwXIA1+9hC9t3lILP+G47UGqHvkCJEQAzujBTG1K2vhljZQc
3sMZHre9o0D0qgFJ9BkQPU+Ty59TTZhq+Nv+0WUipYIwxQiQdubs8CWxamjMbo97xCjfRWp4lKiG
8Ua4Kx3TOJLK7ropwSVxICr71VZESMPBbQeo5oSGKARMCN2xFrBltRj7qTFAJ8P0qKv8DkkgxbQl
OntC40B+oH5yJ9djGMOSpcmsusp1WFF1zXtyDLya/t8Htg5c5o96T7H5N6I6Ti5mKF6+cH8jTGEL
poibOf25d41o6XOqwVyztE9+gAMgr4C/wJ8frFeQLGeiSSXZ0n7YtTavTlhBgSAt+WQa/YiuNrv/
ogB+rAQ4L8xNxiZmQkSkGKJvvRL7jpmUxj5UfwqmhjbMeIH2j6Sd4VonXVbY45xV/4v878L2SLTF
86GiaRqCsDnvq/yUw0uZLZvv+FCCXoCJHnuEj4VM0OYQjocVzvOk7v3wBTBi3KySDDla04hPttdT
SVL0iyIN4Sjq3MRpNt35RGF2GvW6QrSvSqNjRrKjp6UsIzM/up34Ow8YVQyGicWvLR571aDS/vKT
jn1FM/U6ZeM/hON1qsRDHfD7Oi35ZaWms/MqmXU/xCmPyHMUyYEm4zKBbqIKJkgagTI2wKAKD3tI
d1DRZB6gcbJEmnNvnMCOqWoyXEMJZ0iqyRbsTTmj0wQ7zWpWYnZFBpuxZUd44rZ5yX/5wZ8tBPD4
hZjg1/a9iOXHpRUAenAou5cww2shvJXXv3hMsl/v6319lqi1QDq7lB2xn0z98u1P3U/AzK6oKcga
SepoVKK1y3hhd9FrP+J0pWDIoVMYB+7AlaUgu1Y6FYX9Jcj2q+eApIQSLD350iqd1DIUd+oZ+OzJ
EswAmHdpZ8Pk3mix0EkTyGhmCR64YEIE8RUniSL8megO8utLpfjRjRNsbNbZIQlHpWcMvpjzh8/2
ll0AW5BB5rr77aXHzzW906/aMoYAbNEs3aot1S8Cv/ugSujxXlI5+vmraF+OwNP4sPnQJMn5G7rM
yrDRJrMAADT4/8vhz5oAPr+lJrDLS5QAgFW2jL8zenxyHUtGlhUY2ED5JK/i5tU8Xnms3/PxohHi
pTq6/CgKT9tX98UeKZBGuqjOJ4Cz/WvDV4MOiFMAeDFvjCHQQ6HE6Aqe2+YYC4sXjbwzX0vE+qy5
rCUNMNx+ijhIvYXmFKuzj17QSm1UpOjDuBSaOLZbnHnZqna32vUj+DXwhT3loDDhUPvhgjJMC8SI
PBfWP+wA3VMQqz0aJ//N/osrT1cq3UM40UJGRUza2zZC+6OF6RHt2wpkmA8BiNe5/sZXfc0GWrW8
uv+LrdlrrO9BKJZZTKiV+wvpAV8ixlH1QlpbDb027slp4j9Mf1YBhv5y1R3cn6jePR31pvw69Iro
m4oiaEKNp6tSJU1Zg5qpUw3dxkkWE4yNI8lTh3VCE5qHieCtXaDGTEGD2CLTqfpqBpuaNNHp9Xq3
vY1BLXhE1Pvn6jr/P7u6PBwxhSiGBWVEgkcYigdvtemkbYihfCxfrn37uohe8ald2kO+1JsRFceV
ySbco97j1kRto/4Tz/zmzXP4geiSMTYqPhs36PCIxXkBu/HR6fPULk5UbSsFSwi6jR0a3ooq9Ebg
lG2dPXOh9TMe0ssVXVEPsoAK+FlhSCqChVdwSuyfs0m6WzRDnFd6oEFVXN8Jy9wO4uIaXeBr8GoB
BcsvqfAoUjCZGCDEyEa0sfKMUs5VM3tg1yb+LP0EaZ16yPE0bJ7blD442NYJTDGpjFLRkzYExTWS
RuYi5+cApKfcM3SobpHxI2Xt6dGf4fFDN7romC4CizyKPssQDDUdzZ9paNWSo6VzwuP2VgS7AgLK
c4ToKuFW/NvKTubO4fopX+WqP1stdQ4Dac7u2Cn5tgqd0xEnpqaApx0b97bhas1EpNAj4+GP+uNn
zKZW3id8UcbTKQaaQSJX2PnZYNB2sx4ycugttq19oF+0oxk7PWlPygxDfAa1DM7V/Za0E3nf3G+M
/FXjZUTtv0cTAny2SRyObB822UzcLI2Q1m8ijOxpzxo+7G/ifuViSGinahUFEKCVNqWbL2faij7I
34Dii5pC/KQ/zdL4e0+KrChBlGg8KsIPvXqdFVUCRsYH2PpLzUfkqT4vwXOGOWFd/v+BQg7pn3xp
sSrMJ2M5yZMK+tp//mzXWLfjZDFxpzHaOdENJQ7fXJmZINULynInMBfYMhGmgz0xLFJal2Q+hSvR
QNSgofDeTguEBcQ4DyymZ2zgxSaSlmS4YtvJUwY2biTL8HeMcDeQPnE2GuZuXGvjixcuW0FhOBQs
CjsuUZd6tT+6czVMevr/M9IbBfL8d2GXOZ4DTK+vzKpVRqSSYRfthtN4h5uv0GsJlf1/Ad9DTj8l
EVGC7cR3DZxRz2p91rUnV+XeN/A3bB4pK/E/0VzBdoHw4IN9q8RQK9CPg6MtVSbdPwLklfI10uD/
ybtavHrkh2mp0f3//26srvCNnpVpsCbKL+tr2XoZRCo9ro4j5RLtQejsfejb2KM77gjbQH0aML2F
nxXy5z47ZILj9C2qmQpa5Bu+Z9w05efU24V6CvZUNCCCnoTHeQ0SK6ZHJJRjaHD6KCUNxsblmaty
/AjrsTNmOUj6fGaRjoXu7vdUJ/fBw1h1H8rSMj0t/N0jsENHqsIe3hphNR2Ni+9y6OW05SeEpkGR
ACVZOm4sb0Z+Cr+ma9VzEvCXDRHwRZPXqKbtrqAxlKTlpdkQKWelkq3fNvjSDVcrJhZBtDZiLMI7
iEVAoH13SR8PVxz/p6dSpnPuruRxSvRkDbisgbWreOtMGXuqpJQVTLhIzEMRl2AHQVvZ9o/5F6Ps
0WHVHZxjenAuvbGfxmxsBkWNw74H42dFWgRbts32crMmGSMc99vX+UCvmKazRreMxoI3Bto8jJFK
N8g87zhSqMSWoKCb07OVTJWQDrhSDig1OkHuntbNddoEm8QAFmKU0F9nAUIUTMhfyh4T+dompnmg
QkmOLevLx+RdPteSjUwWJJhr4R16pc4gI2YntVpTnmlqRQpe796ZIkQWXk9fPwu+kidpTG000pfH
jIvZHlGq5BYEeO9uwkLURzBWEZJ0vQv882D317zxJGTQmfGICmlenkzvKDjk6RCer278iyRZMm8W
bziqoO2dHsKZpSfyLj8Y9eWSCyckAccD6CjvzxPfbjpZsyWyyBe/IwPNoFO9+i87P7j+F2dQoxJQ
4YI4lWp4sJf5vJyFwKdF2Q+vMyp4obt4MQIk8F2kyB3n+BIqGiOP9T/I/7a7FjDoghAUSdegfbXo
xYJnO/CeIDAFt7Fn7KscO7swuFB7T7/qdSuks5gsbP2p+Pnp+EVZfgVurvyP0GZ2TuxL5RZsWlFs
kL6iYjU5mIrb3LEBNm3PSXSF3TZkAkp3+W9+rSe7e7pa9BAm6F0eFhd1eemm8rUKVMubFHfnzTzm
Gx0mYHNxfPWk3Cd1GYFqU2ziS1aJSWv9U9caH4qvonpGAt7wjvw8RJup+ghhP0DFAym+TWGhZJJ2
4RMIZIUPfXrkg2jvP+3AmISRNUAw/rNktZVI162n4+EUpG2hjmy+eoT9LWKdQ9Z0OWnzvZ0iqYwf
K8GMy+DOTIs61KVvwBHI0GkbjhTrnjHXFnTrAl3Qh4ltTp9fBd7V0c8GgetYEjj7zcwDK8cIIq62
3HE07ZSSf4/O5OU5Z5rKKVPJrfwZxYjXuSDalDKZH2oNVK14IP8IHO2ngZrQrLix9JBxlelcniWz
xOw6xoSe0L7WXS1KWn2MmE9AuO+t6uWg18xgUmmN9sHWHKQTVwxx3XqDJmSiqOOxbiPn015OQX3K
epuCnPBHgSQpe37AcolV+OEdZfReIt2DGE8eLoDp6lG/zjhTDVGq0FSQC614H1It0td8HT52VNWs
lwsHr/GzGow7qUkhlPX8QThwwffZVP949/7mmmnoJhuiDOKZNdjJWWxlqsc1NQLkXkMST2ZYtmFK
OXmmktAyz6TivSvLv3SXQYN4VsoIYikHls3+JRSRX3raDDoNqogHMDGBy044Upn+EFyrSlvF9765
YQkI2wrWe7YvrUHQ6vxBMglJa11Z9pi17WOdqKYzg9c6hH+Lq978B6wr6VMSbzlunGyFuje3H0Kr
lAj5zZi477W87kAezKoJO0/wsj8wJQLI4ZScx9IEnOUiPO9fanpsoecEzy1NfJZv/AsJ2P2n9vYT
1Ss9HtWIwMJqELJBM+mum/NCO3swopNY7uy3hQuXVX59Sy/h3+v4U95N0O+wpTOryb0XhEEGBNRF
YqtC5L/6JCKy7mLP8xIkEnb9zdfVeFfWf9nz6UuJlz7oh9nYC1tXtdyXHpljfzlJ5ZQ8fLPt5Ger
ijng+cA+237PX8fn+4q5Ro6weDwgtKOWKNrqh9s+qQqFTAK4tHOiKFdp5oNAT+XwI6PTU62+NDqU
TaXRGJBlRs+2g3nNSbFbmCZ+KuwXFjzBvxtcl+m60CSo9AHFJWJQsAiogeW1B12Vw6kQDuvb4TP1
X8fsm0Uz4jk8qDGj0ji5PTQacSi8pjTYLG85k+ZrhvT8pE7GEGQO+yfFt38lplNjCKfRfdht91zV
zQA+0+9xUr5iHYSuV1BBMOpawCcxQtWhbvVN/lAPY29FJ+RYUsZQXItQF9YO1V2btle5E4GQqJ8H
x+G2T0tH0hG2mPDqepSzqmWjvgPWaO8trhqrfgfd3w8UL1ekiM4U5enG95TMpJn/3KKRiXKtimo9
c0XHy8y0ZGpd7P58nQd/Nub2uJ9qEb1OuRql7e3POhNgJ/J8w1NSpzjHXgOmAoMbh5rc19w5U1x8
yX/Jqds4LLXu8lnPApFSotJkWmGcxx5/r278QwA9aOiL29d89K9Qgu+DXn0d4hlZ/tTfn+W0VDJs
xN9ZlXc+xjVEPHGU7Kn3dxWPq0yCwsyyzktm5bmUti36hGbuHnxflK8gOBMV00VjrkN8Vs3NFB3K
X1q2AIwSIT2EQWImMl1mUibHgL6B927BSCqAWNtY0vozE6O9VtXgBMwYlRVgr/mE64+2axNx1vTJ
McvjdQiI7YRpk3tkvUjOWqif3ZMr4Iu49/pKm/TQ11sCLZC7esE4zo3mwgdBoqAhzy4Yn+KBVvh+
96eE/Ta8G9LQZxY+SS0YDDxrIzvHN+CUEkkcZTu7L+Wno2MlxTk3wd0gh2WJnDPWNsUYiOxfXfmO
5t4fvJ8RwqBroMz9+xqXyLOWqUsON5dKubow9EKVhfUtPjLkkh+7YhkVDj/nPX43IKpLAcLsDjsV
lerWp/erlFBLaySjy+gjgxCFF+L0g0Ds1BDwpCN4Br6Tnr22PX7X38id80ryjGvdHz7R0S+Er2ps
U/ITSl3X/Ego59DmhscnQvSsu5l8+4d6vexB8UCZ2xNJUMYs0TFbS2dOG1zpYwRT3eYP8kfVdd6b
mQnUTEtKprrt+jzE2ELO8V3r1RZmONoki+2b2IgMagtzawCYWhDBVUsLXuI4rrbWft/khWQVcn8g
1eGtYbWlMzuXaDDP4Fl25qniVTOGhrW4RarVB5iSSOHJVumgzWdEHUPytUAF3fEoEfaygs4T5dz0
WeSZ+moqO0ml2Vu5rn4G3raLx913ZDB/XBR0aEXLqB7tseQdORTGhIaD24IK6n8vn4ykqcqZ6uAt
IVhqCkYQjXKy9pkDCif3i1lFhpIRyWirRCze+DwWp1AEmFgviuJHij2g0NvN5oGKKAzcq2sB/2zT
LE22q5BDPmePXgf006+3TAD3z6dsC5mfqYFbjKn8Lw365Jw7vQ3ORmh9bwovo2NcpxkXKVAw6n96
vWXcFJFCkZQP9cD51/r48g586/6FX9S/A8SQ/b4BWgICeTwPL7q9nHegY9w5MOOwrhMunhFyHHf2
qHIdtKFhiyI7nxH74fCrg/dsfLUBd43t7PS+ar9o7Isrb9IpxSNoXDim8lVj/HOcSEBVz7o4cF2e
w2mkGItS/zHBAEKGiXP1KZQ6ZyN7fH4Abt+xOiTUmvrw/udzrIZ4rKnySVrndGSDfQTDe+jjCmPi
ru1KNd3t2D4Sb7sq7Jr7H99XcqaSZU2Ug5sHAE/L8ycVt3rBuk3WAeVAEZ10Vym3LelNh/uhtvgq
mJeVxrvfpr4q0B7iEHDA6snAyEqaYk7ttxCLiCdsaxHmnphm3QDwFftRldK7tndZMeLJDVL+qFlx
16CrsoO+JzOdL/EtH6+bIqA/+RxsL3kZRtAigPuT1TEBlRAVNUeTU4yTzAgA1Mq1yLXExtDfpOH2
GzcYpH/ZOqDPPG/WYYrHG01Om3YnwSoaEBalFthZoFer3hk509UXh5a8wVuYV6fNVZnPMDcxLI/C
9nBBqUfWzqW2tNHByBnMs7iGzQYRrUZc6TfwduIBNN5zmmD4bGRyESPoGezSkKJBNn2HmlHOyZoL
nOo1Y2Q5XRJ5gvmgZrnH6n1TAo0RB9cKaLQiht8CAAYSRD/g8dscGLIdEBiOu3sXiBGSo33fJhLv
9wMIIbE0CkcDRqYNmFFUqb3Q0cTayCkL2shAgyjatQs6CAK1wH7oFJfmM+b1gR1/uB1EA307avFv
aZsUIySNwFv7RUl1l1ij4DbAUC5dNhyV9Y37YXS8Iqz6GgZCTw+FNpK6GunZFhpWRg4OpfPLbIlu
iiCWCfImVvCq4Y3EDxxrCz3cQ25Gu6WP8U/rusheHsKH0hEdHgAmrYmB/qG46m7C4mGr99jCMCTA
VPlBs0/DLfhSGXTYSftKvb2s4H38F+ykosYqwsSplG7NvlS4B3rb+KKN3fx71dbxf6HoJByue4rT
3/CbPq+mndupE2VT7QzHJcvSm54irGAvSt8C/QYTq4Y0gWMwZm8C+5NjpUx45fejWx2qYSZO9arC
GD0q0US4QxoIi99rGscO2JVY6baj5aGdiWVomr0a7h1pEaivSYl76S7c0kSvL27vDj8yP/sxeo4b
/ELtEETjOLYe2eHh6JMwb2owY9gW4iimj8pV5zVfZUhT9sl14/wkBlVVYcABO8RsrIA42CTczuzy
CxEkn/+t4/zbl+RhjMybx+5eQ63XiKrT9dcqvnz4YpF7sVv1+AT/h3A0WFT+I2ngmZQ9Ss4N7Yao
wzDr4YgfMXUTjf0J1q9fNoL0vR2yoONUVsak0wJ3UC0/+VPq4Yq0on13TcdFCFTJ5I6R1BNyQLBY
tZdmD/u5Ekdgsgzs8yU1t5NiRvEfbQXnUkZ4nzUJtnoQjxfMJcOk4iz0RSBUlKUxIASsvUCY5nzt
Ehewab2m1UZHBk6MJQUPMa221Q5N1gK3/zBhVG0UpQdO7b1670g+KwIBTaRUYjfWpAfwVZuKZ3hr
WOHpcPdzFSJO7kPjVwCRm3UnWWlg31I85tUwxyXAA39iLZd83IpvG+mHOV5PMowjlvXQeEdZ8RcK
dlM3QUnXO31wWfZRWvN/RVaAMxXYKKNQskwFa//gkVHUc5TTUhLqmHd4Qj+DbTYAs1xmfwn5NMLh
4W669wKy8DkU0Vh6auzhObGdXSt3kgi/aozWuyKsB41femLwHYO3Jdg9vcHhuuLSssjCQsO80XX4
C5JGTrT5UX/4ofKwgIvGeToQYGDjtITChZuMJjWw5JRqfIlhfO2/z3etNpSzYsF55kWz5OTwzk67
s807DFE0UneLXpkgHqkRwcm0aflOsrcHGnZ9Q3vVl9wQbfwtumiE68HLxfoZ1dFeROobXmxId+Lv
E5doGa0tM9cexxjhOmBP4RpJQsAryXXFDf7hogO7ObBvp/WrEDki53SmJu1FKZFIhbL9GfgL3txd
Ubjvmy84PnJmTs/N7trwQ20cYdeu+D3vtISv+o8YHQJFdcdhIGmIs9rb3BabpxoPppzGLUA1ofUZ
1QVNaPL7dEelIGxxMZ5glFl5hyM40xjAUYKuIEbQEnRGufofzJj+JHHgvJiZMLQJAkcCb1m2FLUq
SIcuW4GEmV9OMD9Z25kOT+OBnae0QPoCW+IezMi1Q9KUZ2cypFqFbDsMpRHm3ixVKKaemMXUBUVH
kfoCho25NOF456ARqoiE3NgAhvNWRXJ5VUz/p+oe32J2ZN7c4itd0jUJu61rB6/af5DUncM4zsV+
/ZzjeK6SOGPSHP6a9pX2YjmKoWplExKKvrRVua3w1+Q9PGlxE0R9J3pxG6AiT2LPaNETvJ4VtFW1
b7zWuSqGQQSaASScg6nXxubJYzXDhOqH5s5ybxKGR65QJa3Z+N7VmAYXBOjEpAHigqV2pnlcok38
QK0ZxpDocJMcB44wVVbN4kv+J5BtVpZLuOPPtYuebUc2qKVZ8D5xhJfx4pMRkKcXXwFHjHsIezKK
J8aEilW2kaz0CHAqrIigH9/7AmQ9w4dtwmM8KDmEhIzE2EhB4I20MPis/Ut7ncnEy/KfmsciWHzd
6tadocSJ7vEHFcw9z6/1fjn5SDvZSR/j6JBSO8a/aS4ehrfjUlj4vkInUoQM3ZmCo/syn+QEe+XR
cdfEWJ1Ul0tId/XTWCk3eJ5uhjdQl9ptJk+BdFvfHePHDqXAjFBV4EjbmSLYssqFRXSsd+hcjUDj
3A97/14XikxxgmpBsLSKFfJ2hN8UlD5LFi9WhDVmW2H77yk+rZM+g1hA/0i2arNf77lj+C8QTCVb
PDmIjGCKny4Nc6yGuCFXSTpb2Xs0Svn0Uv8aUJpgbSg6otlCt5V66JP95PXSOE7q3MrjS/damTuQ
OTELo4Jou8ep0N0CE6MrUTKBR7/HbzLtRfwbVd1tERl7QDmOtIj97qiKqzuPomOtSS5ChN0SJQcR
zEVQEvWw37LHuPfPIvPIgOQ168rJkOh0y+aq5xOUHkrqQfbNCIS19sZJBqHNr+X2FcgxacNnQUHZ
wx7HFAst8MUXWWLMQN5ZQ+WfNCrhEXhAFC/JIjd5Tnrtgm7mNzDptIfMWv+Z1HUl73s2A71FS2a2
CC2iZam0nbK/Ucbo0QzrdvuTKHCCQRohbM3zzB/FbvRpRR+xGcsOCBhD1Y1E31a14ELvhmM9D3FB
necW5AaCwDc5stBjHQ99dMmZf3jxhNQIr+ge9J4hqiKOCqPhsSjk/s2GVtH+qmAU0v6pmDVSgPme
pLwc9lu9nmLC8/cJPMHaArjhJY/yeqDYzp/X3F72srUip67AzBXQr5lInjrF550AmTo43+igLJsU
r8Wx/8zQ5syiLq2vvGbxZ6Y2VCWGJHlmrhGv+w/JJUdKZ6DQDsFiTa8oKEPFF702va2HBWx0L5ee
NGe80ttjKvsWB1suLVIZtPkyIl/hExO4vuV5H/2ZiFM/WtpE7oy4BnkD2K5MBA9TExJi4/tjetYa
b6JKq516YZU//dHGTVlDOnHKTVwYUEG+15HGIPirLgGlqzkvbQ6vp9y4wYpWpq5TuzqoLHmsLeaq
Ygm+Lf3a2G8cJbjLsrWg2g4jPT0srn5HNx7BV3CxWuvF6RvAL44bmxr6Ud/k7PXqZPAa/TSnp1UI
sjHo3oWmXNlcW5s4OM9ZZ5+VTmn65AC/O68QePD7OQqAFzSo+fcp4bBhFyzr1aM4X33VEo0Jox45
oiYjITezaeSAt8kWvPJ+Y0A9yYy0NA9nesMM2N0qkG3ex2FLQecleBr8ZjngMGPVCI8HQGpzS63w
N4YHPlQk9uWv+d9LSv9txW0skVO0ektghuBdprp/PT3NsQgbVgZkh4PiBqakEb4H0c9v4GPx2p3Y
8buAqOZgHEoXyT2ebbAjn6Jxj1aVGZFMm/GvKZhImlne/ZsfNpQAKXrjlLIsfcDdqlTwCP7Z2mHS
MvucuXS5GrC9svlia9s+CA4UstoQK8EyPPaTkBAa8WUb+COriT8JYW2BsG5Du3OZxuj83nL2n2qo
WPdWWY4OBcTgCJVoqqH2a/EyPeQ8AbICbTaS0PHaCmrGDluxlSggR6mKaPug9KU6hnJ9r1X9lQUT
CQsazxxgnLCqZJQ+KhI8RvLfWHa44GjRLuOUPeDQFNwnPHpNq8Pa6hHx6W11h6JPFantYPSs9uBc
GpCI8JTGAlrEfNPg1MOgqasIfM1RkP5TrxV7ehg2M710OlLa6eHIo0pJA+FQKoatZ9bHfU0Ug6Nh
XzLvx5V5A4UrGnqSj4dvFR60M4ihqbdvtubbrks6ZB2Jqh8EOM9gpflmYLI48/yzEQMDsXfn6kZ+
jVNeyEf/0ETjGSwTx8UE2z/5V7oh7FyniLvJwqNzsgu4a1EAut5QNq+uGxfsvDOehc3RYKo+Rkgb
xMANUY0Rus+b8BuOM2aywC3TCcqBh2soL8ySE/48gW90aT86lMMScY1gLKg44dLx3YAMggkAoM0h
6e6f+9KB7MWDlkIVJ10QxOHrMGJssV/Ooqv9Cr0Sk/uYda/u7LSv/oriU3y33Qq6GtvTQxx9d9ey
e33Fw4V6RRn4OkLWv0dn0ntC2UPh/jEFZH7Euc+3AXi+9OMHOpU8JF3D1qJYKgbR+yyjxQm5GqkY
geXqneC4Hp7UhifbVKOirM73Xxwpbrkvda70s38uy9DvbqzpEfaAx4h/jjFTchxDegWWkOJz8tsm
3Q8LL7PVqf0jetRWb8ZzTt3ZtQuLchctUoDFAI/4B8ZVuGEY6bYNITPupYsYfm5ySU0XsVGl0AGV
b4h6ZumRv0OT6xT0THXrkzhmf7PcHpzwjTvyHeJ/+oShBDbFZHhjzju/IY2HV3bRtKDLwBBfA1FN
SJVx0zFShFAYu46OBl98ctfquV7GBTflzS+RVbRIj8X88+eHaFz0UuUgmJe8rlKJW6CgLgF1TLjv
Y6pigkbZOC+V1DloPmdESncjmHdo208bX1BJv6cTfj/SzIY1MCGqqtxIFekYrBN4ZoCay9loQs7P
xMROgdXpSCEK3KUR9qvvN+2Q3xFmT75ajaeGgIpu5mU/4P9BUdwslVZb0ruWVR5DcG1kBhxpucri
p6R/VBjQX86rLXhmo6XgQWa0J1+Zi1xqvoYSPtMm7Nn0MAT4KanViauMcivD71h3wwralKrgFQH+
AuWPd/bf8mE6s2Qllg0V52ySo9ZYQiMUcBAWryeXhds26vNF2+veqRrJO+/VMkBGDzIFxpFcII+S
pFtD9zWQ9C26F4pAi6Goe6YuuvCnmd+oeXDzCLTP9qM7Y8LKlYHLjQ3rAkfRAWolX/qijxYN4sb3
/tZj5ouWODZEVHYhyo0Lr8KtI0j5ARumSI3HMK8m8+IkaDexyDjPvlfSZsu5K1T9J2LMG4qg4Z4A
hNJ+eMYxQ8mmOoRp0IRVy+pBvwAyR3Nq8bZxkLQNYLYo8066y1BxhpdPTtwFyuvRToNDZoaNlBqb
FFldyM40ErwOjdx5GH6HLtdUyG7MrEMgh0lLe9syV5I97Ggkz+caT80x7v1gG9oxGJy0F45mspfp
uxdSQEsPZHCu5IqBLI7ib7p6N9JGZRORqsqaUbVb62bRUe/5qo+OpnmKWSp8Ks0OmMLtIPclPZoO
lBJxlg8KtheNl9AJ+XzUP2pRj0GbkzScKeNvV3kgSgU7Zmiz9dwrebQotVB0hr+41fJ79BqKHw4b
LLtw3l0RBb1FevotzEwRqomkHXXAhzrstaDSn0kC0hEGMxDaPIb537+MF80mTBOStgr8+87uROoH
uEMCpzDK4k1xawzaWYtmr/YQpNQ+6vTrd3EH48c0mSfTUXp/HcLFlQ9/LFCJX7NK7L3zoiOeyt2G
zg8MQmCLs17O3D6/s5PJDkKTA4tFpipkKqggnsA2KA4akjE00dNTCyK7yC995HeQyFhr9qwtvqLP
Y/7U+qgSxnnZjXH3nOc8aF0eV2VROYztEQN7FV3S5CfsB6YJbZi24PM+AQVBdIWgHfC6+WoKbBTf
oBAWPjB/T0m899y6mh0FYyKkXF09BMim+rL1DnjFtyIo+7d4J5yMu6kmjf2iGKnZClvRvMKVNKtQ
oP9qQVay4DZHjyse8pEToiZpulqsm5jIQ4ehcEYr3LZnGYxi8emGlkjgtlbFMLsbra2k/EIdmWe2
j3aR/qTV8osOfqGVYvQ8yHQIMAoHLeIv1tjwvz8hDS/wDusARuboWR1MsfQ22V+320NKzkOOHsuU
tM9scSszwV6rVLySLkBOpa42BP5Mg34EhLxLvXgu85CcDbhv1C2KkwL0iS15VXXU3XlcuakOQJmy
yrILIxMhN4pTWzHo1HxlUteMTjByBpNrNWwDy/XxsVjEPVmvxb/kHARdgAP0d4qAT8SukBcXoqlT
N3TeKK1Cule4hB2uQoWC8S3a4NVnlubAhodGqIbhEz/UnQDIHFf9tpoKf/RC+7C/Nr8au1c0tXfl
zUzeaiFzN9bJlRK7ZLL5FCd75iXUw60deMc3Utpf/OtL4dqEPdGEROUrWO97LE7PmP8iEZB9g16J
7xg94pYxj/Lqs+QbKlKTS2ahhbhq2sOqOijtXuxJ9BhPI+OfDWpiUAV/2coJHDncEKrI8tSHL1XE
GKYeALv2g/HlXUSj4gy2B4QCp/R/BBYxxU0xW8iRlWNhs/xpxMJE54F11AOruHXfnWuoIooq2Orx
xxkHEWzWXRcGqFAKKcbGpLVOD1IsPxo1a7HkUz9yLuBr6KqoUrY2lW+mvGw8kBYfpzUpyqlS7s/h
xp4QljDYPXnu+8dK7TktEBAjga+tsCj+K0cAoD8kqpRur9Jh0Dp2zga3Pk0G8SUNNB9vo/jh85bm
x9ug6Zn40NVugAszYGKZW8TkY/W3RDAIz6akMtwBgyBccKK6eMCAvyfh1z+M2q7hupo81O2thSsI
IqxzPavbor2AK0VRvVpzLxW6+hVoqsmz1DtdyPAn7W17bJkdlw3wsm2bzvp71wCDRDB8VRaLMbtD
7lLvKnhwAozLSORvq+3BXiTpNlvBYLfHoUNarTSOsGhPlt1ef/1kOEatmnNxSne7o/H+Y/qbz8sF
ONnvYurQkgT/VJdyNyxHvTiSihPZrHI5kc9XVtBZDjCJ9dTzvNjakhAvBN7h0Eb3m1kndX4+pmrq
jr7WAiVcwZWVeyj+JmUVyisBV9MR/Ozw12hLE0IaB3jeWkyMbm9YObWYzMdDYpOvdRZxqx2539GV
ON3j3fVxEBNqqXqGtZqwuUIcBFYelYwu/TYCjvszWYm1y6ar57ynA7vG25OZ+8HO1R52iJdA3JZJ
irnJVLoiBqYX4VSDCmkmgqf2XfNMLhrNqZVTYAoVcInEG6LIXdSayklvhwR5uDxR/jATjgd3KmGr
Fbfmf8yFLs1HBGRCLPiZXe7bEZEC6xtR+7TtXoN+b1BhwMqwsQo29zILQISRP5YIE0Ze5Nlpswhh
J8duW3bD4ZYZUvxia1p7C9pUvxW4JJglcyKTZZodDx3BrV3Bb9TqwsezDKJ3euGeFuF7AEEjYntM
NrrIH1whXjjyD+GeP5IBwbYlv5wCprrDoQhSJg+MGGyaGFOitUStrvvbf9G17Ix1TMLxdFkfUwtd
wIhX4TnQKL+alDPyvF+VcBbUAOMWuIp5DEqCZ4810qLbQJQ8GIlBKRJ4fsUq3rnQtb+mSXITaY3m
9sYuVb6ZzvmAox+ywIrxztlVur0+NffxwQsJK/kdzoRG4DoORpkMF6HNBOUkWx7fn8pqpUxSJxZk
34yQf1FwPpCKIeYcujy3pfR83jTV0aWUGiE/7O+TDEAeMRbtyFpJ1a/3JWeskeY9cq+0rvicsYst
99d0RFb9zjHu7UPvIx4XDICrdPyBB5dwCFAXVYdnRjci0dP4+RTPE53cgeKAyJHNKtWEhHseqqmO
pG3pge1/x1CCRDfYTl98mSRq/gZPlGedeaJ+QWz2l5DkzubVtPd+Fy4GnHY8HXxOga6TUNUuYY9P
kEgJuMeaE8LaJzcLRdKj3amC5N59dKH+RswYSYIyIC7EGpuSQJkqpzrmlbz+xd0IpqKc2AhK6Um0
DsNv3qSkzejTZGwQUED5wa2KdRELv5iBz2Qa0YzlIKBLTf7WTgGhR7oDcWFSB3/OgV75xqmgf4Ek
hDlkLSS6ilBN104txqr21qNC6Qw4NA3GkxgToL6hLxSYw/GZuOFLZBf6XyHWdAo6T00xgZ05Qjkw
ed0aX3yiJiksAoE/fLGk8I4fRn3OuIh+rwMlOH+INjI7/hE9XDHMdHUNKT/uLrhWPw1gvHpcUsuC
a1ztN+X9lG+Gjhc2XreMtWxQh3KUASGxyO1GjQUhDm3/OmsNCfkfIqjb+nR9h7bJXSydIhNF6mET
qTR+Uc45ulyWGyezUbAMovMClKy50osAEa+3GK0Yb+xaZVF6N7GenCpnAVJ/0SkmBvzgglk1Dr1w
5/o0BCCe18iZOCsCxeDH6UL2MBOiSFoFA3l/oT6k18+XqhvpaHye3m3g6DqZiwY2PgU3dlpUxFlF
q5FYmwdjqN061TiLJt/YiRPiSLQR5P8XQDJHWeApi9caLPE5xV23pwmIg5zGVA+7kQBkcIrlXLl3
0QERUKBS8eSz1Zwx6nZfr+3BT05Rgx4fOkyRAbpNkpz7dvVKXiEBFRJzpSHr2hy2we+EfXaj4UDO
yBVIkBcCYCOXyE0OWktAGV+ouTxOdnLgRTzE6x/I1LnDPBGrSDHB06aphG8rNOFvdRF9ibh/DroY
HbY+XzOmBckdduGJ0WSnhn+2LerNMv3V5HVNXz6rmNNEVtBAQyZPbcVrSBEDsbg6nFC196YpVyne
tcYLv1taV0GOFmNIoSnXNv/VSq7MiAljI3xlRjn9w1ogNPsM7OZ9KGe5PKy6M1QDg0u6AWK6JXuo
huu9fRVc+V8TecfOh+/UA7oNHLTBh1EZAh7YQ8zhgHGOExunEs2Jh+0MbSTwSycCZm0Z9cR2lsYp
DbDnF6UotIPhsSox5EoEK6V+UKPUmiVBP5YDMVOsIY9j1i+W97soDqWJ5IXVwCZquofExytxhpvT
LAToyMaFdHutKgHQ9Ftbbjxv4+EkTScMUGUbVXhZcy0Kyba2vtqlMp6GOUhueqTxdmB+gJ5FS+hP
dIO0k4Bl3xSrRnIfv0km2wgT4v4WezA3JJkJLtFgv7uWY/Jbmdf0csS9E7UIEyM2OMLLzpmlbdLf
U3eckrMpnVjB3BQPvOazE33wVEzazfzjm5RzBaGGv9AKPycNsmAIom2Fz+vjHnWVcb/0L/7fVNf/
n/tGvZi3JcoiZI+Knrc0xShnRblnxPRCx9a89bnGkOKe0MpySWgOb7Npc78PlJJDiRXQA+qo2fLB
HU8uneA2DJPsmZfS3OgaoRTj8BJbJTahpE3cMM1OhLvRoZIxm8kL8pcyM6eVBzI1+r09qbxps/St
IfaWFxz3rL3F511pyQbYIHxrfNRikUiGJ+7RuIHMZAMIM3mtKFS1/P1lL0i12J6XATnSpuYM2mj0
fT7KPprTnRl6HnPNrH0GsVGyaprLaL2lLv9BU832SVyw+UlRHBUSvqwXEl3ZnLuMeOjYHoOVby1b
M910x8z8CXwcaxoC63/EA0sJq4cG3FJcdwajTiZWM3YlcYpEg7L/kwwc8isf06q3MReGV2D5mloj
Iz3g4uXMxChwBXerIcpMrs035Ms2W67NTvd7ko6QXMMUqk31wRso8sc4PfIGUHnbdQM5TjEGAL9W
fCT0noyALfYunE1JyOND3IeDFJRQSrEsBRgdTafycVKYze73h9EbYvRilUxrwgqkAjRCi9EDexnM
UYs4H6S73LqUhu4xY6E7LOQrq+VxzF4e4a+b9MRAxHMY4w5IgTtey5Fa2Pxg4UeXMXWn+OJt/f58
xZiG8YtrPORL0QMiyqsgaZm1GwMIqA0N+lmfeGvfHkk5VBzGXR4zKoC6U0XgRnXcL9yXf1bdIzpX
G8V51iOrr6TzT+5VtJMtabQyT7oitBY61gXfmV56kypmTASkm/jXVIyjCEj8rTw925Mq/fRrnz69
ZY82AVp8INO1oTIsWJJvhrwvan/9GfUe3IjmScBixWPqAv/nhybQoHPyPQEV+xf5yu5y1LK6++86
lAsMA8mfUe8SP3c5C+tN6ZVyV4vBAJkX//SssThcJnpkFDJ5njFDv6F5fsNGIIIJzfq7lcyIqcT4
/8FSfbeNur7A9ekMid4jDUiwTCvKzu63PlVqa+D0AQOJviJozDUwZQHl4BsCTObO7JVG+i1TDMTB
9czALnTrdKbjA+DhaMgQYAmEg159Z5aUf6kDLEzG67+TsRaXwdUMuGeWNP9RgLZO6WgP76an3PFU
s/SqhVn881d/lpjWaAwbl1Ged0u41JtEYehOK8QT5x+9+G1eGTnoGk0y6dv8YKGvWOcuXzmvN55x
iqpYcW4jvI4NgVfUnvY5MSawCbuBGfEJedZOOss4YAUIkX9ZbcTqLftKZrKOZDeZh1skI5B6Jei3
/GLpnVdHM/fDaWTkZJrW0VWBTj8jXXKjDfZT+Wj3dCCHDZrwdAz8Qi1vr7c76U95Xw6zrkOR+rEJ
QutPfzA7w8vqRq3ez11vBKtykvoaUSzN5il+cSAmstuhvmhlGtxr3+jByrqwr91kkn+iy7EZiRCB
hNqoQfIav9zvOHVjwYpak7zP73x1a/zNAMNOiHQ8f/ZXjhdBmF3ZzmZ4xNXVFLEuaR0dJUI7vCA3
sWUB4DPCun2Pmxun1NUTLqXlVNGUIPpCtrpCDiPJOmwVH9REogNcsn2HQehyF0cA4fFIqtf0LXRv
kM2I8/V7cDE2HDv6+fyecMP11Kexqc2i5ZhMDHQttLISc6iklWzG8fnXDcbx4qRrB2EiQdT4tdrv
+Fy2gZmdmiRnZJ/U+89UoxTGAO0r383/0Epv1oerifdE9td5r2ljXnvuGEMuswcqddgqVfqmsMyK
L0cBhGa2c2w/cYINiBQj+HaOf/YWoxeEDAku+leHqKSUCy7QHVO5xAepGgvBARnLEAputYMc3qyu
b0Jp6PMC3tDsrZU8xgUFAr7jxt2PpngegVoLBgN7E4xvnrq8hg69DU9KwsfEm0PH3ZAbhKU5xRnw
X+k/gl23E9YqVd8yd1MsaboZv27BpMRncNbQmu3j2hXQu4inY26ptmFjIMUqeb7HHlHb1BsGhLWg
gMoFRsPW2wIjn2jRCQediGpC7rIgb+xKZ4oQBB14dHpfjQOs97DztEH6FLZ2RNXv9i+oOZBtC6hJ
h6Qn9AoASroe/ut1DpqHC94PkOmNsBX15rnFDef3JeXQM81Q7IZ3+fi8n2im3YH2sSXevbWZPuDP
gSumz0mpgejyMb+aUJi0mWDsYXOyJnm29Is4DrnQ0LYVuhISW9LYdGdDdqoaZ0C98PHi7m5FrcTk
sCmk/YU5h1m2+ytbMGY/B+76a7vUp7qg9uWTtLuEYGVv4X9wJdL0UulYa5p3kXEXB2s3gb0H5+dE
KblbdDaOa2X+ip/T+aKQZZrWnanOy+oWd6lfexJfNJ4prsl/1QRnu6FHhgiZddJ0Q2p+d3RBuEbt
HFJYDSs/nT89yVbPtybWaQEXky3wgtCvwcBT7RHPhj1D97yOkkWvjV/R/i8SSSdxyWqtNamgtsLE
mBeN2lkwSg79nH/iQzc0qGmy6hAT6YQJNg04C2uM7zxcOViyW3leCW2mHR11q+kJuqGiUOOw9d8u
FAfel9JGLS+kVsRh9RekExs0qhxcCcS9Kaox3FGNDisajpkWXsOA9vNRFnMUqnv0QEF8EfwSG3py
Q5jTLXx+AQHwF6dqeRHh/ctizoXQdZ6YVk2gUeKYBiiT1Ly3GzfjB0nyxO3TKQhEGLjEM3AxeEDU
rCa0uunwviua35oWTH07UZRvwXvp3F4ZubP8kpt+5uiwKPcRg4Q37tUY8DZ70Ii6yaj/XLTFL8WU
W3AwifxqRRzGkPKpzWUp5E14B1EdjrwsJt0G4Z2JXnPCA55bf+phNCaUf8ydxkgBRQOmh77oeVqR
KcXZ72GsXV/FCgAJJG63LJMe9iTxz1wCJ55pMxA1LyyJJV8/sPRAHvEKutVF4BenbxuM1dbXma54
EmMGUqzYZ83nUtxlsurs5NJnm/8kUkquy05mmXB1/XVd6p/uxMtbwTYKghdLN53UyQz3UDuFvzZ+
JbP2ymCK2idbE+9BFjxD1P9xbCIKaUL8ji8jgMK2mZDqjC2UMtv3NVgIkVMbEBQHIpY/o3ylmuhO
/ZVID8ag2Laijs5CQTo7gIyLlAunuxuCbVxQr6KsmUkwggpXj4HA3MMOAmV3dETwAGomzyuJXTkf
f5R9NU/K3vA0sZ6bO3n/su+uv2NyyJzK1g5QGjwDjQK0hM8ACHybMg77QcJmVBE7txMGndPAMvxk
eCH8er4rRgZGkFjgM15lAFZr+Z8BVUvUU52dmE258wEq8+JAhI0Z1z4XruGjTVFD80GrgF4KimWx
QMqUK+ZpXxg3OK37QFqqjzNfpCfZ+Hflc/i5ZwraPjiFoJgXq1RxxHtRI9jecQoEZrVY98wq+avv
KEnwKIHjBONi1mzQiR4fT9vvZGk3zea3PHgoCXv8O8p2jTJBrGFTH/y7QL4giP4bTyvsWkakS5n5
QP5VMdFMD0M1BKBHidXtTzhRAqZCfnUlNK4k8eCvunv/zssw5TWGD69GhPYvoJJJqF1/U5qy2ToQ
0SGbQP4yujIaQ6z+3nQ3hz15m2XS/l7PYa7Dddwvc1ictRa27CiONLmDDpRUhZWF01bACsL6UrAq
AueW7jU7Jq81kpOZkZSO+sqI8dFVMelJp+QDCbxg0/71oI5CJ7McUN+38eAsXAxOIIFKLiOyXy2z
hlo787gxUfmpxvTRmWJxk2lceMhiP+z8lgoS5+VvosTFKeOrLd8TobANPaEYB4CxpMO85aJGBbT/
eutcwr2JiO0rj87tcUFRJc2PsuzjOZRPGIXM6tJK0A3pwQJ2DS29USEOvf5IQD7k2Nwskd2bH6zu
ljlef9IYYbPkAHgIpbKrV9vnk0jBAZiaZqNI3FuBxw6kAJN0JlS8AIn5IKD3OAXv1W93xnIzg9z6
zseg2URB6AWm1i2cY8xJRzR5n14BuQZE0Lj7bAzSdFdApLYS4K3kSB0QRoB6K6E6m1mfQkycmigc
CVr255/KcJ6fRKidznDxdGpGk4qafcpe4nAvxfUXa+btdCX3ra5J9kav8MID/XPA8wPejooBqI1W
IqcsQAz0BJ2Y+BUw4iPmak3RYIFO79HlyhVsWAHUTuNeHdUD3dmKlkcmnhGb1egKRUrskSmYq6q+
OCyinQXNxM0sK10ZSShNpSj7wOdiZI+Lf7CA0SN8TK/eywG9zfyMNMmUFpOKIrIGyvUWHpEtnJ1/
0X5QNEC2RcxXhh+InpYXgvaGFXputRUELL0eITdx+y8EkmQFknr1FnYoOhH+ODUf9z2cjdHvTXmG
AogfNvZ0RIfLsRD8vB1H6pMTal2KKEvGJhKWwRuMF+lRgLDCNoXvElBLPgBKGvH4s0kvII39b913
5BqMdncu7XveX7F3lYvr7ClVI+8TvUmvvGKDGTgi4P9VR8JXgt//jS2WxzbHtUtdUQ4p/G5TUyAc
9JGTB1bQYo1lq0ANE//oMJU6VChejazdzn6nfGOuXD82zr3OLc9vKr80ve1y7kzub4PRk57no+z0
t811yjibkR5j/+aCNY7dEnolGFDr9CLzhAicJG8OkgPgRl8Sw8QO93FxMtTfeQi1RCzP4esmVdez
VCtR4OBtWH1zMyibhYgdJrg8PFyVk333BY2e0q2wXLdtoElzqRYbNWvcna2kyOZP9T6Gu6ugaw2+
BZgqp/RseeN94GI1omAlbcm5f7IN5ggciKQ9Ly8zZdMLjxrJLWWfIuQYr5K8qMrRx2ly8C0tJmDC
/PsD8Z4pB164pqM7p6WfDVbAwD4jOItmJr/aoAKPu0NdK/zUXK4IAA4wqEVpnHOxHfWdJ0/4JBEL
Ua1GRUNOhOOr0ZAWzHJ6iIYmHNX01LG03Q/f7IgD4aV2rfPlDEmqDzNy65jmQ5X8bDjv6s4DgBuK
t+VCIMfxpoXLp3cV+UlhhguM0HiqfHLffubP4U8Rf0N0OKxWANjbDilLUWJ9O0t9dc5vtmn7Gzx3
W1dBWKEH5b18pH9+TnvLfvbSSxR5q+0Q24JCX2tDATnhzB36LIcYq1s7TEwZ94sQ2fegrIaTjP/8
ZcD6G0By5VmsakWSp2XoAwLtZuEQbIoeeN2oxIyHEl8NQvSrBEF8KRZv36zx9GA1ZGnFX4TYacnx
qfRHO1Ca3s/HBIZFOQma1EmLixNaUFMGQknjga1M8NEylKE3CYzR4vC6A+iLoQ8ijv7HEQFrYxV6
VlqYC5CpHERErHYXjy0G9U8GHb35bnUr08JbBzkOmjsBZf/5hxPfeDFjYHT/KCcXpVL0okrNXkmO
mlnsy8TmMAkMxay43xGP9pyivMC6xyWx/c6W0PzYcxorYNrIa4IpJlp+77XuU2iubNzFmyOI+m2M
JaYeYFJGxbyM2QacvFmbS7vMGdiag3rzVSlsAMw7DZvOPdgFlDKA7Rdh+7kfSycAiVfrevE0i8by
F4m0YszRkvuTeWs0xaHUJB/xzFvbBretweAGfv+hGk7JIXVUpnY4oR+JErBt0WrgoRBQsIar977P
G00SWZU+jwpmexZnt+qJ+ym2QyOYQd+OuWFQ22810Ch9j3oI9fOpsqZX0IgyOND0Zg0Rba461aaX
ZZkKnGT8dWM+6q5oAzg5/Gz+hMrJtkVqQdNn869rXseUZZSrgFUZO3jLbp0rjUuzyY/czetFmNK0
nSLPVsscgHk0aP1MdFGlvXTWsLSZ6SEr/f2mtwH8yKQuvt3ArhNLu3cODdA8OGpXF2yySh74fcZ9
M6m+3kFWtvkB/ZhspCwXDiqDeeNrwnR+8AJuxy/4lybxyZR+fDHFulavzLOg0EK+kxmbx0qfbI2u
8SVblv5vxOtSjTr8nDCw1jmeczRLD1qBw9ZhYgqRzf0Z1cuBqOJuueCE/VS4F1u+c8CWenBXw7Ig
UTY/im4SM588X/k9ye2KB7BcG9E8+N07WS37nSdeO/GvD3Qcvo05+NL1ZKPDSpSgKdTbM4gBSlLu
p70MqcztQOAWW38ReUmkRjgsyGbz5qLUSNPVpP8XyuTxTv/sVl6q0jRFPV1X+OpU3XZnXe6v/ubH
FxjoElDxxB5nVyJu8Rbu4owtkKK4aXf5b9TXTjgm4vyahIhjurysZefEq6sjiaO9/4R4Zg9Wf1HR
eEe5RX+uaTyoukgvTHugcMz5J6HhGcQMwFqNt8NlU0bEet5kIV9IMFpQy+pA1j2pTXQD2guPZ+Tb
vljBMepkyDCalmwXJttzFk4DCmg1PuIC5k4rklWk3T+J/9b///A7J5ol7E4QG5KNs9B92Q5ZYr88
0tZHTTpJK9JxgLexnvfHUIh3LL4Z5WW0Us/ObDIyYPDvpVO1hl9chQov8khn79s/1AXJpDHcWhTu
s2C1BcpAFrL2A6RudCStV3Xw0JmePAPRz3jRYvrcs/hQ7OU8ncwL8iBECzzx7I3kgev6iU0Qfubr
9y5KkeDtlZnUrCsqxdcvvEfKn0FZ3BYa5sS4Ab/MLQ3MXQgf8IX8lyr3TQFHVLOrLtnkaElycdOB
JGydZ+MFeG+0ombmxOwK7HbSETTbgTx307op8XhxxM/jM4rtYa/v5O1nJDBvTnUCjFvfVxOgDF1A
lS1aDCEuWl20StwE/5Js1T+7GCoeWutDHIyJwBgEQNKH1KGH3zs+IHOOclrPfTAaddJj29noYgIn
0sgx5UqeY1EUDxPecBAJG9nhvyP/ya6zSfHzINRepKzExz71Q6r7O7YHP3gyfTNovGhSdkh71R51
O03G8C7NYXb2+JpsSZCjCj6g3iuD5qCQdV79CUlYRN9ea+ZncHbCnA+pIxpTy1nO1N0nHmgG0USc
4AjeKx0AcfRVXei0FVl/KgY66tpxb/Rh06GGu/NGqtA3xjQtqx5oCDehz8O+nA+/IsAmeqBK+O5S
Y+GnnLh314ZYTzuEqEuwCt1qU7N/fnjGVGvf8NZjRpbD7ARt+NeKW7X9kBOXGjsU3rRg0gsvOcw3
46fg2jT00OyUFxi6lqD2mb0cz1KxYc8JsM1Pgk1XlE5b9MHKWrqpo0cixObvZ86J1bXIfzSriN8d
GD4A1AdsFT+QHRX6kxlO4ToyfcAg4McqzDDYBk3iBLCMQ9gvlUxNNvZTI431y4q4NjUBHZyO8niD
D+Khm8RGJYTYXzZh5nUkB80W7UN7WnqaueIdgQrjl+D/mlF3VMkQN+nFLuf08b7O0IWXtOGDotuB
/awoUQbsYYoGXZSKHHyMEQMswOYKJ13Nh+PmuSFy+rsrHfxghCFbC88aI22Un9xkMIHYu2TYIiZd
vCaA2hlo3FOZGRZdpUV34yvuLMA9YNhG2DEgh5MBe0oAjeGJmmBaF+AS2A8pzTnutJAIju1n7j0k
foivr/lZamfXQvTwoStFGPozUp6yHOulObKj0tH2zhK3se96/LPNgK2eCedR7ysTEIYcfhzcHwVV
m3sJYY+PQFAwHAepEfx597/qHoBU3wk+iRBSCxbVmcq+7nqGNjCM01VtElFfNkDJshgOvY9W7e3F
H08MvuyBypwbFLxcWnEsZHNk0Ztpl0pelTZvmG1LouucgM4qMRCvuDTK3svlRg5dY4fyWpUYCY3e
G3+HElMe5LskEgE/SioNmvYu3tVVtXHfmLKZwtZL5Rtb8tGM8NBuHsTVeLxRXN+MqFnhUuvaN48W
ghIxAa/ztw+XKZV+LkKA2zsfrWJEzD8UIqLg5dNd3SvtkDQyomXBRvCPMfA28+Os9atOKzoGlPZO
D1wuXggio4RE64UvMlRBzJgyLb62SbZTogQhGzLzCNz7TT0eVGV8llPWh7tnn2Qknruz58BM7xhD
JHwbeeLOrWivH8Y7NiXNg9nzRa+ie+G8kW/tsaWXgeQHOensIwyf4EjEjprbhOU8iieV5PnOQUsr
Z7lY35K9Yt1sTmR76Qpcbx311hn5N9ykLt65XTF5OgInGOvcVIEIhQ0lzB1dRqa6t0dlUw1iEfkR
djFC1QJVFqzR/vxHfOZ/jhUen5oNn6GgBaRyUB0gpjiy0pfwS48GvsqSpE5cqEyE896tjasCS5wU
mKH0hwqFPWMIWFztNK481Lo5CM1+vnfgqAKbK7h9WqivGaK8INwlO8aSoJKQXCAv4jsXocFrinsU
oCFCDAmgM8/RcFKAEHGx2cQz3aZb/zsiINbz79H2r5glMESK4v/ONrZ3i97vJLtXGhkWcU0uCTcG
vMH6x0uEiEGJZ7p5dN/JBtkmD1uT0eRUabOD2U/Tc3ZQzQMa4t/mL3r7yBRoeNo2EXzYJ4m6gx50
SdjlPCAfQPXzVLPD4Qyi41O7fTSpVsiALfW2zxLBvHPnUnLI/20XTCYC2R/+e/tlYQ2Uwg9eks1J
xFvDPD6EgLkb+z9lqLXdd1zkr6HI0XtQOJrZAiv3LGcCBhuBTkX0AD1nE+deD4ogKgUgo+No5Iyf
NxdnAjm6+4fx+0xP13QfKvxIn8QAp3gOlDXXNXKAaXGVxYtk1DQiuLiBXOfL1g3fm1vh6LsxZUYb
cjnbCEFer8Q+O0AEyUIGpuFxSFJKTCv70Ahq+YmjT5h7WBAkLgYpCg4XQNzoYhoUAZQC7modcnoO
hNhjEcvVT97Lg4MF1iRCVAggcF/J4DC/LyrztJsuAlzCIhzgX9VUdw5LHKvzqO5zHwyRxWCIj5p8
tjaV1u9pEh2xneJxlaSpS2CfqBHiQCmeIafDQ/mia4dcEv7RH5zqBVKorMzQSVXkhjkZgKJdxiMj
X5FQz+6bmIj37538glHw9bd3PjcMpp/LmHR6tNuEgS0ty/klOzJmxUuxgnmQP5PKEK1+qlcZeHaS
3FhYWsc23XsxAn8Uu9Vo3okdNy2C+rThLCVbul7M3Je0qlTlMeJlU94EekU1K7iXYs38LV9RCm8S
unpiB8agFzm2K2wKgWXD7fZdTuGa393++1eGFqvvE6OFoyQqEl/PCVogkLlO0lJ5Pky3L9V2PjC6
/z/M9APIpSwuhMJUKreqCKYT7kILoskzD1619ABLjKdFrV661VSEVFQWibYcnO4ZMSmv4a11vsgX
yUijU6gUBm7/tcMwsKMlfdE8TkReyhpDayXaN4ts2f/nhwiSofGStHSu2uwPINWjfEjCgrFMl1dM
XGds90JEx97V7Rif1nvteDYms4fYOZsUahPzmTwgY/xmHz1i7K+xpDi1/8Rw5pTRo2ZqZnQw8Qsw
/ULvfHfcrqYzm8YiJ6OMwNk5ZaJSlSZGo2Xlz2LCpVZHRQBmfenbWsQwTiIF8qiNV1gEUbHgopDs
9tAinip15WxzlvZQrNYWXKJDDuM87odeSqFhVvzR2aTbxvF/0+jYKVwGGcmjmLE1u/K+nqlUmsin
q/wIxPje3NAeH1LKmEjoaXxruwJPD41ZVemIY4drlrRNba5q24qZW0D08+Hs8k4FNme4htN9dOPt
1v2iiD79jR++G4Z1eXEZv7amHWTfNbS/MJhJyJ5vWQpCx4JoCcF4qHCrMCoiYjaMVHAjkxLm7PDc
XN2r2Fgu+19b8LHj7RmtiAa71u7ZnIBP7WTxidRYSSsJzECnhVwGZxBD9L191Zqa3z+w6oCI5W41
bP6+lndJqRoz0zxx8y8tEAJgyRw6zP07swCSLzdoAf5SPtcesz7Pv1FOnJNO1JJX1MvvFZW1JAve
jaAlhyRoUk03OiBjf9PDBpwDYL4MkKTTtJB8qwOAhnsxt/4w8w1otEU9NUAzHfKVpjjGayIrms+W
8Yyhcaia6YIdjb2sXWPn3rjRDtR4LnMrCh2HVTVhMNKFzhmAWPorRPlzEN2yrM6wIDxbkG3+OkXJ
n+wTSZYfrBjCdAsqzU4qqBEAKyZ3OB/bc6IxixY4xxSRC1fvH79hbZWAFg8O6ZNMI0MQ34MEAD8R
WFppRQKfO11gNqhpqw9Pgt6PDCGHRlPDgSNnghZIMRm6foSPAM6wgmZF1KYm6EXZySVcam/7WoOT
PxNwoeeChS6AERmbbl4InJL+4X0nNnXf3JkdDCnQ5+CkdAtT62pberwkGXl1qf0pm1+5WMJBCSwL
V0NVML+NHLV5Qpv3M5XyE15lSC18T6LpbvObHv9nQ6s7xjySyWRXzizL5xVLWuTjOQl+j6shgkcM
LquJcDMtnUwElB7uILgcZRf8eABpuzwdtIgaNZpQoGxiFO3lZGu7vMGPVayXiMkZkC8ixbcipXsT
Y5VvQOPd/aWtL1J6Z2OflY3VEcUspLCvUX3+9B/ktkw+ODFVqUSAHchbMC0kguDPx0i3V8otOlaU
7dsbpLuoJ9ObPahbtTOAOW3JwDt0QXsuM3ABUhmeE4J1cnrknzKxFgdJX+ddc6A3Crr2UEA8W32F
Fk/L/tiDwmycmCv5dN6HGUOl7/Sdd2VXfPWPuhp3zzjOk4HgNGPXH7SSw1Y5Czs6o24CmKiXBYES
fbzt8Czc5f/LbHYJnJy0lSdAjlmD6aF+ZeCTYrOKigQ2bCzxe/nIjo8W84uJJC6VRG6nqQ39Cvpd
GIkEqYfD7S3rU0S5fPN1/z2ua7Ke1ZxM2+39atdQHgpIKPSqZoTd3faoVUZPMTkXMkyNT7rVxG2Q
ikXC6yGCYuaLV4x+YMDFNeV3pJqMrOoG4TGoT9vGIcQeRk+nfyzOwxPBLEQ+mATF/bXbZFejrgys
sTuLN/9eMkFOOW7s/nBMN7FIVwNF+sjUyapWiueAfRk7OHdJAtO1p2wBG2WabZFNsJQV5CjLbdZD
OA03jkSzZqJCg3mkGPfCSQq4VW58CWqcrolmbjvQGDfx/gd0ZZMqHsEEbm24+86Yc0G7DpG6G8gh
PgIj5zpwOzTKs4bjLs0r1mxc8jfJVTBCZOaa2sm9mcKFFKb1oPWaU487zKwMoXoSlByueGCi0d9k
sEyfV7nWWAT32ka+PyOziq4CgqDePFvLISvB9ibun0FiYdUjvq5mv2wfvQLltSiugCyrrrslyN1M
ZJVAp3Cbt+jgaTNYf4EDtNe8TUtmYnP3b8NAASO/qXVPJwkFLBBnAwgnyUG34p7+B2QGk4UV53iY
LBEWfJf68X+o3PKEUqK5UdnY/uIT64M1SfRfeh/AmZE1sDfyLhpiUkzLzRAsoj7TTkT2PCzp7xfn
xEREs9VxC4Ub9qAGqYNQhUbAqo/Bg6K29GaO/60Xlb10xctdq1OGpvRSV+SgU15xClNLD6hhzDGm
CZE+pRJvmtbmInp+yhe5rMOptmXBqtstx3MXDTOkQc6gVuwUtFdoHcBDcG0oDsGccCSDFG0fpzpL
4Lskmdx3CIn4a3mZ98l+3IoVX6vjG948PlkJdb5vl+URQCP6pViGeqMZiYuPpHSu3XFLnhC3na3u
RCGCkBZz+9cac2KyF+UuMLGUIuAKeokZ9WM8hHPLQDMmLvhma5LxqaSGR0mNyP5lxPwHq32y6NR8
VZC8zG9xk20HXb4FhRhonthMD6P/+5H3Tg+U9DEi9T/v8FZ7AseagwFnJbtMZuyb/afyaAhqjBN+
mF6kwxStFcX2C+abfLiG5IiF4BAoEknz4TsSFSJhRUwktOffvZK2FKtw5vj9jk/cawByTd/TpXVY
p4EXY36O5dG4gz0lQsFQGGWsX4BCKqHiunhkQa7iryRXUrqKAL0FqdnveEdsqUV/0kpPOr7ar1Bv
YJC7grFvWceNP124DhWJOwsULEkMfRZpXxJxAOjRQ0odUw9SpjClH+gp02BVEGv08ec2Mk2iwV7E
fxjaqZ1OzWq0QTyvoIXXQdBePRouJBiRYIdeJvf2UMromS0DskOJOX9u8C1KdSwYKdi2qOGTiHMb
KF6Tw07/5vEBKRECpmn2I4g5YTVAMSrQxqe4S3z0qEMrzu9Xk3HYtVddXJ3Vak4cIMW7wPlfjynK
UBNDdd+wcf+CNNqfc8Cd0NrWQ9JbJEvJSwimcLPhDBuxB8OK/r1bSBPqK0Vru6Y6cqOcuRfQ4i0e
Y+m04z0h/VMfqwX2i9kRX8440/q31PhB+2gh+Mu4jv2aFQJJrCoN3VFuPRpSXnmJEfuJ+DBG5S67
6dRapWMCq87jsFesOSIFPim/V0mHdtsDvo3Nl8jtFPGch8FQJtmA0Ygjlib7nrUjpAYPFh0MX5+l
gKwfL7HLn224k0mA9LxArT58bNyq5DINU60IqMevqNFouMbgn9ndkbaPtQFEAakBfY1NdOYnNVpv
yREcsla6l8hO6LW6pNOJ6CkzDqs7/hiMZLIVUi07URqYsflwXBXFSbyC80jK/FIzNygQD3Bgt0Rv
LWgsewPBt/vd87vJnXRNdDwdu/SWKubk7I7LHLAf8doTQYmsfdB/yiTn9Z0rNRfuV1sYwFNmsyTA
yphtRb7iODr9NEBdRsRkxWJtC+hmPsj8xmKb01jc/LfnV7x4qVZNmo+SFftVkcf39JmWjE/k/R1W
PzPI4cswK/zI1mOKpORtI5/8GFAg3FYnp789vc9ex1YmSa4zL5w0mafzou0jNDyTmN+d+l4Kq4L8
yN0giXtJb5KWQZYiVP5p4MTNgEzXiQVxd45yE4w9NJj1mqqNjm0CF1tODzR/zwEvtLet3bqflaWg
jUHh9tsSHFMa1IWJcSiHDlrI+QW79dvfaVm0Y2fxegagO9l8GVoMuIwEe559rsuBGIE+1FQTPZJu
zUK6WP50sMPX09BxUP40URQ4g3+JEZ+JV0PylcJboZNNoQsuGU88G0EKvIk/YyczOaoVtud8dg9E
CeETqAqeHZSXjhlvW3K7OJE9Olh+mS0iXPDf/hFAAHIH0p8cx4TiG76T2Z0+0HOIpcGEMPPuwnHi
mz73DfFbGzqgq3RgCRG5+C9OdNAJisyiAWRNqYj3k20fyMjdTunA8Wn2WY7EgP2YHRj2AIPNimSD
1eUA+R6s5v7/qW2XMDkBkeVBg2appHuvg4FnVPUDowXDHcrFK316TKgbBj/nPlEfHubsWYtBM6UV
Df8A2ecizZsGevE454kC5iN6TRAaQpguIwKf5+NULoLmheBtOHZuqCZKKYzvosZqhKfBsJ02P+0y
GN6l3LU0DQdABHrzQT7CAbhHqgg9pc4dspSXp/HH6QQxknTtil7ZbzUAjz1bylj2+Qh4SsZZtmen
aeB75RNjpqqeSijzBm3RaAP/v4Fnu2iDYj4ET5W2FexwD2drvSbqxU2fvgUChUh1OxkFEiLyd7dj
4WAhygiuVsqZN2qexxHWjMvsWr8zejkZk5wGVSYlti63+bxiJgYp3R0gKsz1HS9kc5BeETYgWsVq
6dBx1aFzZRI06C5Mrh0Xg5tx9Gb/zuZCwTAb6Szu7jGnlHXDc9bsbLrJCvhQfsN9paIiimQfD1Rd
Uo6feHx5U8SStPZvcjcCv7BxwiORy4qF2fHmLpG85+tW+OnGnqjp0pgXO1hqei/DDlrWU5Sor89O
ZAPmxjG4kL77KBO2HQOPnNqgnHxgXtkxlBmkiL6FTqtkrSLlOXwKw05pnN0cQSVxzFMVxueZW04U
xUBKVy8MyEHnq2F4bHGBi/dh4NKbW3M2J+UInqILOYXdtEuQ5C55hfn2s8JaDkTfkPYM6sNUfb8u
18Q3UW2Sd128P/zuunN6D8P4O2v/d+0NtPsJR+RPQ6Oanw0g61jD0KcY20HAJpczUhM79PK7u7cu
mvJZP0fb3KHOE6dceS3rLdCSLl612MT6lN12SrGiuZ3E8BK8uADeOrl+2kBlqamqthcmal3+/K9s
oQD6YLRlPVTXNii9X7s/XIqg3be4qSMYe1qybfMY2EQ5pJ0ITf4x0RrwZwNH+VPGo5a4RDMZ9lZr
ke9zH5rgGXq22HXaKBM5dgLmBfIe7L0PfiPKrY4N5gBOmIp5PirOaSiw/NWkTCLUGau+K/j2HfxB
SVl+vKJLTFCkE1c0axawlGDTF3mVa2w7q3bnbYBFTnNCY7UwnrIm1hR3DTNC60MYFJ5jEd+oqeNh
iTso3Av5f47K4Pcvnf4/IFksZWeSmwFqgwNBt2UBwQaVgRVR/GxYaaIVBFykDyq+py3C9ehGmMgH
CLn4TcYHDMsSfhMfDJ/uu7TBpmJnLiOcIkh1raCfov4bNAwejKrUeWzBgYDDKUq5R96nDG61qFnG
Yp5ZP5v8XjDvUl0JPOEkLlv6RtNtDn/Fnguad7FLkdhxOODf2pGPs8+I2+cB6T6wvgR1DelhZQ06
wEcVAZpO0NO1DUVj76QapnmuzdludDtEJiF6umWHy6qSpwGCok/b0UoffvFyHJNWAKznzXa5twUl
wbblL5DxwKSNSC1604iRqbacQiIlYsUX4bQYzuMwVNTTjhJvwgglq7eeZ/xtLvhyWG+RTPgh2EpK
GYZSjYD4+E98i86CGTY8Peqv2bxHo65aD/OppHv0RX83p+e7vv8zS6LQuDDXsgtLl6dzqqEd24fi
q2sNLWH2qAzGgY0o2q11IcJ5WmEz5XrLvy1rzSBznkDeD+9mI1i0EPMirOd1qSpDh/miNA+sXc3E
MFAdT+mpSwk7OBtRAYSk7e231p1Ho26yKbpWuKKrBwjQjndFQSauIerRNP7wL2bKT1vR1pRvVyxv
UXniOw0SO/hLpsy+gE08dB7gcn80g1T4Gx6lF/sDSxnXub5MujRyrvNhmpNJJ4s0TsdboKL0sodB
PV7gjLCLg1FbTvl3EjUOPAFFqgmSfQNJa1Zw+jkBpbzfLjH1sbfFFyWaTl0peeivntP4D8wXPdus
LDz8Sskb/NlVJLX0mvcPJ4RkHHmloYK3ymtGJHY1k6/CLjg3esi/T6iju7w43oc1M9Gw9zDF37hr
EGjCUHlrt5B1cf7VaXnB4S7ZbqXM4ajyS5MJMI3Yu99jlvCGGU5vK/V9v9yamqQr0xtSzbIqFY6S
iHAlY5imwgHPzOiXrrf8v70OwPH95A8zaVSUXgjUWnUF4StvmvcXjSwP1j88dsj/Opw93/rCuCyE
eyNEpjR0bg4Z/Y373qvsgeCtsLKCFKRVaPzrvMWR1U+2QEjUIFZ+qxNtntke+F4OTdhBwkxyb5Mr
vXqDSUxdvfHWscpc4DMwhl5pxVBKteV6mSUsrUCA6vrJFVIQUcXKHUYiBifD84oPUgu9ELV49Ii3
Ux2OrYnFbJIhL6/+/z3Hg7HX9bbLHDK+SNsm837Pw0ibvqsaOxVSAYVlBaRAhtmaA5G9Zj/3ix0L
67AkXGTHeYYkRoTtdmJvYpDWHuXdyA1YUVS8UBNoD38wUe0iKW2mGAilPO7iyMMa9fs5focTYS1p
PfvoBDC2l7Jm+/GG1PWmM4AOt0dzK0GGqslqs13LemAwcFaHbqfzJ2Lf0DZ3rKT+9wuBAfRb45z5
Xu2WgyuF9LbUM8QwxFVDhqteKoHLmzQZcCA0EiCtGO2UKK/HbU3ehm1vVXsl7g4vWIxIE7iMuX3f
53OgfZwuF0NTzgoW7Ga0HGGmS+NwTrjxZPvspOOb57L6dTS7b03L6FsVn+YQ86UXBA4GZYkAwkHL
YBOjpBBVm5vMQlbRxWA7aDLDBxaTrf5RvQb5W6v3FPaVRoz4MMF5uGvX8xWZOuilHpQF04kPDfcb
hrx8QCwx3Yp25mU2i+yyAoJ45NSh18rRLJmkEm0xEYM6xO7yUPEZ6Te99ehuvQ4ra9bCWXNut1A5
qUYaqPMo44uOqalD6lPxh9HFqLaBVreaALeu2wZVNstUKadadiIGeotySB2LtBdBGO/odyC0dnZ9
v19V3YzeopTjmRvHh6I+y0JnZKUuCZg5njO4tFgNgGRWXme86iiTGdyrLB1dFM2iGphdmVA30TRX
/tVgwEK6ZDHeuB9kFN24rzvuPOWtBWPJ1NJ64KDb0/mwbyfzL+EIwoIwwYzdS9rnMiV2JlOj60pL
F6IKBBV/wA7TkLp6OXgy8uNKzgIs7mWd1tjDpswOffTmaw09+dvGtMj0y+aiO8QMDvo7c1TdEmxv
U4phhY/OVfn7fj2XhZydFb/oUiENEfHRgXNB+AA8JL1wDbuAyzou1Oc9m12f7fKGWdtWrchyCGEi
SzIdORo5OEG6dTE14shGGEJegZIdaxXZxrFsKiKliMr/CY/7XEfnagWBmKRX6dBnp7LfE5DIQe8e
SK4/GS4Jik5+E0QQOVvmdcqWQ7dtjD278RKJDzQMjWqBZyjpBS9wH+NG+eQZWfXmds5/fa6nBujE
7r5shJ/IDbh4GkYVmdAzWjBO76eLjV2khFUtQg1O9JSpe51zpjBHBvoKYB02+uYw0OvCvjbAgDC5
xfUEVkOaXxCbMJmB2+HdT8k/u3DbHGJ3KxlbbK5n//u7ZZ6Aa1sEqywIeNhb0l1X+w6s4jeiTru0
sDESHaP8YMUX5cH9nuCb4U8lEwWNC6AO4DJrzfwBfvpHTys8NMB6gxplGSVIMmQI347sQN+OS9zZ
F+2ZqStBuquXv6hLMjP67tcDDc+HAKZAr+ZJKfg9v2DBWQO3Ek5rxtE+Pkzg5lA1k1UupfbHzefh
MrmWWNNP2hlmyZw/ODzvPS65r1CPBQUd4uz9NTJ075yd2iuur9gzHB/p4NW5ILB15QwE7z4bmHZ5
zMmtcZKMd1LE/rbj1nH7ntWFoMUTkMvsPWT6pXMCgh1VLWqma5JfKhGJRvStnMSpGjhhO587Dlo8
HmmzZNhJEEEMmBRBYsA2l61SqXm57nDuppc2OWik/Nb3YtXpVprcQ8IS1OSGvMRXcd6aWAhIV9JZ
tCWaWYeQxCul1pJ28mrhHEqFkQsA5ZC+QCczo/ME8uIxbIFKhEqT/xS7HUESoEIurHX29X9ywHJc
hHy5chs6mQCDq5jLlSVFjiTm26aRWWThRlfFPfIbZc2LX1C+JvZuhA3jqcJ5HkTZvKkRQow2xXWx
XK2iZooiGG7ZtLFFBu+him2wI4UJp1flkgnXyivPu1wgx4piuyCAk1H6bnoG6yXmjoMbLXmlTBqU
8+lvocBMcjWWIjqXx22lwsUq91SuOub6r0roTjMtdT5R4uU9nvmFdouZ+P2iJWQfNbt0SOmKunWS
pgekOs27iQP8g7cpobVs4NNJBWceG3U/dzkA+FstTCd+9lm+r3QXlfoON5VwhCUdwjXPfOmBdRs+
+EWl8PgpsKJMF2fDz1eO2dsdbMRRjCuYGUE65egJAiiI36FMVbRZ/TRxh4PMMKe92DBIlSbwcnSL
Jl1JGhg0qfqFMAU+nGD/P3huVHCrl70UBsr84bvgNCjsae92FTNFet0Uf7eQ88jKJGQhTQmQvNVZ
IOddWot6YpOCw7aRP7yvGmt7wAvsmww9KgEILPf2FrWTeV6Y6PG7Kh4XeqmF9yGOBtR7vDXFkU4e
UU4oHVDgLhtoOI6qqj6BuaZ5yy+amnZcPI//mwagiNhFmCukHeQOZTmUOdIS8O5DnpYAxnfUDqOI
DUsjPIpDXoZs8zB5G3jhFbd0tUA0wRPpDTlZPcMJXLMtOIAhnrMDcWjrz5hxvALRnzb5WqYMYkaZ
9xQHgRsHgo5PrqBjpS07OwLnWbT/ngRHuHghoe3qd9PO7VkYlgkBVJttVgmWBEEt/o2SKgT1GQBh
oVD9MFPiJjJPAjJ7Fhlpyqc22Z2S3gQMuma+iKgVZIYbx8fHwrvOdLBIyTu3sKZGyzXUdY3bmGDv
llH82N05vJOXs4IqKYjXA3Mpne5HtEALC0Aiza0eJwvwhW4eV5SCOzF+J5Vu9kFnoVlSBzbu3gSd
WkLbnQjqeyHwXWs1ECoUBwFkp6tE9gYpU8RJBzpHb97e6xcGmUl+TKsl0ynLokcOyKkdUdguxQYg
M9bssKnr61l3IPXMK7/k/StsGN1L9Yl2oVQGJhuolZOvkcZ3lHQMezEA3GFUYK6qZUSnOQ37JAT3
6+kiM2aQxWE41XxxlHQS8GgYwIHD9IETwpZzdK35MjHYVvZGW6pqU403uEQ+u5NoN8cW33KbfsNI
ml/Po2euGAKLCpj8/OP10vdkuzCfG/af5AMkIJW5pRjl5fCwGcBgBqkG8vKrOrBSMoh5CqhMmn0f
ug2Ggtyo78AxX+cjMzuapWooa51wq4Wj0cjvuySRg2L6bGTBkts2KbuZAJ05tFdlPLY5jk8THh5I
ATkgf7lgdu3MQ63pAr5ov6XlZE2tHaRPHyd5ZML0bfl2iKqHYrjnMgLiRPB5mQ5DifR5H7vfiokM
ADPbAqFuJEwEHgJ476aaob7BR6lL5F48NL18tAGXzdJ6h49c3dzRIIh3K4+6iK0NAIUFFQvCnsHy
7dbhHSGu7e3Tm02BAxjmZiSxVmvF3GejCiufisglkQkrjMLFn3Dj3FvfniDx805ai+TktTH8l92a
L0pPGpsWGiXdH/oKsZYHqCHNDCDVw++7bI9HpW7iXTW+Gnzid7FI+tA5eo5Fpy1TX9N8vDSaa9KZ
aAOy5g2QYYoNWEvOmaU+jh5tmHk2WTwB0wSU/dfcfMU9WrCsCVoOIfPjYoLCzL1ee4+L1jUQ3O3U
/fR/J/pHB8NDaaz3Fr2gkSFVTsHk2E3NrZyNvXAw3/tVR+T3EN0DYrppzITc9wAUEnaTcv6e8oEM
tpZYUwSYpkV+w+NSxXuRIiOIqqJhZX4zogsmWXdfMmSjRvcYEfq6BLAlMyPMex301oNq8CIX1zHg
y5mkr0WU3uYnph08Th/EpxZaKPyvuFD1PxBDy5KilLhUxu2MDPgJH8sV0TFP+wLaIy6P+xtozr5m
t3MmUSl0W3tFxLw4ZYUgYeLyyyNGAC6zmGDNMfe1C1R97w/M9aiiLbSJqn2YzkB+rR2XHUVXFpNA
7fhpD8/zJNxyMgRd+AOUxdCNE9RpVGf6/+WTpqSVgiIQsUjFlxk9cA5aHW9co1FRcLsNh0gwWQDq
e2ISx3lUCRNDMHfgslQ62SbMn9LNxsO4M5dBRGyjnHphdDPR4cYFmDWVkwebuVusaErh9HG00Vch
Db1eFY8ZlVjXeKKqLttyblKWfqMLy/HMjYm4bvnGddcLwKdLXi77qUtdgiwXu4z1/Jr8Wwup20fC
iZwcLD/LypAr9f6YAqucYwA1nH68b/7CTN6ygiKkMmCSemRUxY6Tq/rb0P7Oupppv9/lPYzqrzE8
dxoZ5g3pmO3q1/UfJBQ50UKFctS9vSXiKpZGlCF+4UgbdYetCyZU0ebNCkTU18Kc5LqWE0e0J7fx
sYU/BG6oJbmXdnPswFwUeBjQCsrUeTcVz8sPuLz5OFE0/Uj6v4NWnMoHf1lNW1RGgQDYxQnpxuyy
LSwBvgXanSKuXJCP9YpXDw/kfBuQMb+ZsTAK8N7MKDChozDiJe8LgvLBSizOfO35Bu/1/Zw4ifDg
nk3hONNvlJfZP7+Lg5Pal63SpSvNQtJUcVbijVPahRSTFGnhJo3UJxg6bQLK8qxrxsSQ/D3+J9cm
vEdBtmihfQ27ub4nRTggzydkTIfAQMo2KPPO1K/s0/lhlCOlDCRinXQo8Xc/+uaAceRX/qv2quTQ
4d1OgYDmkCD99leHN62bLuQJoMFIJ1umjfl7QJ5urqiOyh5LLAK5CvfvS0DoKiJ/i+bLSxELJx8j
PtjFxgN+5U3LRMDkKG59HtuiVrWDJGeamjZvY50hvmBYhjbcz6rwjL25Y9axfFLnEOVIV+GsLSSg
0jaWcJ8r65pIznxYOneG4E+VirekyJeJ3qbnIZ+EW1nIfpVXblMk0fRFbjWxVnd7Q49C4H3gP3LX
wngeU2dsVoHqkvU06t+JTA0L68iWMM1AeT3zvfExO5I6LLRnIjNvVgnRULo2FtYoJ3iLCSvMdhHk
BNPU7+mClXzy/II9gZm28Wv7QCd8Ojd5fLQfVofyMhLK7hcgTw28a+ef7C+aGf07IyXXAxZL2N/Z
U2Nq/y9sGnF4NsBtLfSyhNOB6PlkDwQExG8H6hWO0QQHLc2RF2GiR/AVskByAUCEIbLJc1uyBMoJ
wTG2x2CtHsdnZKGO8LyEqgJFqOgaGYOS/tlYp3Q1boTLZqbKjDvDTaY+sDAwP8UtH9GRu8S2v/RW
u+w7VEgvqU+CHYJiuvq/F3YIxI/j0kZ5SE/2+/v9jxe0T25bd0ZuhR5LL2Mg/Xka0V1GcL7YBSBE
2EkMbklFegv4NdWs88cW8JSQEJoXEwgaMetlout68MPhmYQDPSXGhLwVyHXsTzhOyVcDA9UZAsh6
IZ/qJAieGHyduY6ZMS9hMnqMUIvruETDlpc8DykhBe1pbzvr/LW9iNxfrdoe4hg/qjBMR5F6Vzlb
aTTwUE3Tw3E2T474V4qGAncq0CpRwLUBv9SoP4SjFHSYk2q25f73I3SPSFuj6UHgl167lqokBI1I
U/RGw/RBoLs8vsHR8ZR8UNrC0Htr5JXox+plZuftcYUfmsdu/FBB4gWMlfjf1uRMQAK6QAT7USjF
coSjwlRVHKxr6OdJExxVKblkD73yWjPNlp11yyNxodARZd06h42QFSgC3FwHRNwQJg6Uj2i1+98/
onakftO9swuKCkR+nc5fL9MnW8K0KntWN3Xsx0fj3kdaKNb0AkFHA6HbIviGbJ8b/jgJ1vVhcr9V
xxCVRv58BxjkYVWMxqeySsOkGEUhbZEtgMhE3iC/QsnoJ/AwViGdHodZTz44IPuwJ/+glefDqAMA
KitkeS0MWRbuhflGQtEjQ6Wwktq13MHnKxCnQWku3c2nWfo3fP8tf+IZxO36elw92syycv5XnNpZ
O4njvCftjXca/g6t5jmQmBjHm026OqI1di7VD0YSP6Eq+xb5sptDgT3kv1aO3Vp4e6qy+l5/2lYd
kf8/QUO/vmfJx5RIfQhwzqkmEJfzh3h1wM6zTGc39W8tTd4V+uKI1uJ69TGf3G74Y+PcwcN9rO3D
+0DhUhe/jvflyLN9i1+lmq1wyQR85tjyWX7c7DoGkhyYE2Ed9NzIa51nI8umRcO4Ez3QKQnGGhav
3xmefUSS4b9TZGgX6BHsYA+f4rUDZhxCBzEcEsXZP8CHWf+qwiWCg9i4hMzFoIysi/KXBQvuK3ra
NccLbY2yUD+EnEVHqoI4xYOoCFArOG6o15i1sgV9GyZgDXRTdakra3f6JE1+ZMuck46bQBKuGHJv
WGm85s9TRSf4EHJE3qCQmRK1AMshNFtgwKlonUDGmPFDcy9PN3Vxw4yzU53wTT0F3H4uDN09oATs
WhybVCDSsTkFJWBY7kzwiZBqWm2guWCafjfVyV2QMJwPqXe0w5N68NtzzFrE+hZKK3wz3iOhAva6
CLiaTAKYy4HcW7JpBRpHPSTjNheNl9OdA7M8FpbzAiy3jgXT5L+ZQ0cWHLdDn8dLGyBjjnNUu7Fn
XUJdQgY+L4/NX38T8JlspmGgW3X5fEhojD07UVMepR3gGZrQmPm4j85pjRvs5pUDkHHr0Wrsd8r3
3zVidRkd5UDfP1qm5G3uJCh9jNYY6ZVPp4En0EekQkm5XAHbqIQMbMSSAd1q9dT3C4Bz4jBcYL5A
6KpLV6k9TRGzTKSxJRyEZ/ggylawcFZW8oDkG/ao1hT4PsPMlOHGChvOZ6G0g9+a0rJUyqJrDtEI
RmLJ1XC5h9+rlo9dSA0RodvVC5DXx2T0jDNI3oxK1cBRx5K3YpBhZUufsj0BmqTXfnz61NwsPDw/
PVR1fjehjknc40KW/qhbyVbajtxpGdqOHqTI/QsrMP4amz/I9Zd0slqgI4+aF5rQTasIXhuuTCfm
Ddsbw496vV5QW87HaA2HvQij4cNnN4h4YEBMJlBRprrkCvLeFPQn3TlgIFsjFswspzrn6sFGMUtf
Xos98Tl0qXFw2C5bohi1pSYuw/uHwyzph4OZdxzkte3WEPuo3VVJeQeEV8Q2/v6FCS0N4iyT/pvl
fshkFaXbHUpgorLUIfLLHNrilpVtIW1Ju+hBocrCyeP6FVgufaY8CzLMJyqE73bX+PbRUvKStjJh
teoVTjyl/YvacMiOv3ASwFu6K7XuLgbDmrsNzaUrdIvPX4XIcImRV+5tO8xFjq8QvHSx2tMDKWac
l10M0KfZ2dqguGvXJNGgRHM7VHh7UkpEGCvJY8HEcFKDt4lfU7smD45yft8GDN496srlWPqSdJeS
L8cayO5rnC9/m3qlA5ChUfpDDa1Vq/0lZKyWyzZreViuRecqOnveEkgg3FtNGDD2Tazug+44nGT0
43XGv0PxjVPr1bs514VOwrZlk4IWQIAzn4WDOuNnFKICrfO7Z0BCpK0fkP2auQXgPzyFlFjRyqQS
SxAM00oA9rxUexueFM+gFvwC5SGFaLxl6+Ci/rqOEzrxdAMeoBGY8tJPGR+CcaLYLIS1w6y73n18
YXDroeCJnKxkaHFosciPrG3cFEIjt/towX/oKCR30d1eh/+Ic9mKSnaPr03PdG82Lx4bFHx5n8p+
TDy0T+u1zSg7rxiLsNb/2QcVMpLzv3rKhKGJNDuE8Z85FBmnb+LkGNcc9buoPtpnQ2FHaTo0/P6g
/Zo12RUFbqzVdYY3PX+yU3x+IvWEAGEiCI+a2xKrC7sxVT3wJHDd73+qOeVYJhwHJWyoJBxnNIqp
MN4bxp0W1qCYPEKloYj1OOeHEpUexuWaf9dXhlS3pN0itnYLCD0ivJVy+gugqQkReXu1Sh002Hhb
CcAvOGLvShmfrF/abcSUZpgf7PAjFmudepGO75T1/y4R+VOVkJurN0VB3mODpFt/1ZJvp7fGeCg5
8sJaNhghSTk3Z/0Vpok/lM9fJo9gpSD0x1zM5CpWtL71HMqXo8XSBCASX7HFmiRmvllH8RZlMACo
MuL6682KcxZsRSOYbSql2SA0swF9tOAcBlMC7tNoSFVUeGJe0Q2JbL+iLuOc1foVroQkxnlcVsUH
6Zwt1gpfwu2HtwsCGuO5kN6857rPjCj2R8EYpQiEVFDn599NR+HLzRXSYYiBDDnkmqRhnsmQY6OM
VLRbrZjOPtPUCM5ewfRg/IKW6QsidbzE6YAFEaBJHZH7+i8OMJRLHn4obXiMSEmVLqjdoWGXL+CK
o94dAKc7y47PcwIeOJ8iVMyUk4+/N91Qzab0Ex/ur9wqGrwpgwwD4Xwj7B/r9djyL/gHiTywi6B/
1r4V+mcqh6Viff0S5UFphSA1WUdsFOz6q9cW2ZglQ2V04atjcNXbNZAm0JmAtqO/qV1BmLaFW+on
6ba4m0mrA0MUBmH2NDzK4I7Uc13H2FPH8+i8Isq/Sce/vdYH0mD2TvvAYiBIuhj55lxkZzqtVjlt
KZGJXcddCmNNKbe8b+bU5r+fsQA0Bg0ngdidDauxUcCAjM7Fy5gG/ccORVDZlLxWIcRgTFlEPtBO
bDs0hpiwMw8RhJ1uwo+3Iw8D5WSgGWQ9OazLSSDhhsZ5nWSa1AJYmPEfFLiyQXtzUeCd7hqO74jh
ewc4uDtDrA9fxF9IZnJlsC2+I2uJIf/BdttT/x4h4lmYywDdO4+yqY5apRSZTziUOw3zB3qqLuM1
gxi6ojPQG7fPsLBAneT+w04sGdR8cSL2sZukTAtj9pYAMJ/jmeDloue42/9ErNjCYhgRNFFtvmYi
n9Ehzgi+fHyh2Nq0W54yhf3dzjTKVnQ1JnYTHhV3D7P+jDmH+BMvEVCPSeM7t+CkbZcR9h0Hd+Hy
/k9hKRI+e0GQwbBor+3E5rnura6ykQfr64FpBkDfWvqOzV+BV+/djBh9BvqIOPkX5ANOc2BLGHRy
S5Al5f+rdT0qTRgreN8LRLhiVqhBOPizLbiRqYZJfJr6kpQxtTmvtDb9bI7sBGQpnLk08L3GqymF
I3Mc5aBKbc4eZFjapHBPKukIoM92zBIxiZo8VL19NMPXqiNIEg8DjAYSs7HVq1YrHMuiVYNFtfsG
xjSMh2m4RCBBeBoChZy+w/vXDa7K6OI51uSeErY1tDRLxo1kbo8iudMU++WlopfsYAFvCkFgsd6n
8IssTeSJoLhUPappspeg27WjMan+XdTIHf2r52lyeIDs2Q+p/ZAsLMA5EKqiPZm+lFqOEB/vBzpx
/nzwbcRHbD2vkq9+X9n5O4vkG7CyhEgPt3isDF2jF/TeDfk8qZzR2vSE0b0f0ejLhRo4KvE2XkNI
PLTxcd+H66mc1DmMjuj+TBY6ruBV1pEGcYWt+q6Gbx1J0RRzCLGg0SAwCbU/P4ywHkWHH51HGFoT
X1OxH2dB5M/yCkNRQTjlVr7Gy3Tvu3Mv1tgjm/2rQ7+3FuJ0/ieSnIaJ5xq29KWj3KQGUyVUFhaP
K0AOWRyOv7iOlZk8clxVpuVWlJ+7QoVeLeKK3NtSM993apKANVjk5lTtJdAxeDmdRXSksbAravOZ
BsOl9aqkKOaPAteMFG1sAyaoeJTviSicsLvo9z+eE7QKXGMmd0b7rkFh58YjL0tdFOXRqoTCGbU6
vAC+76cLAxs1L45EHbI1wNPLuRd1AqSQ3rePHp+JkqTf9FNDRsF8JF+9k1H+zptCdZgs86WxnFBD
6PLjtFcEIYKbhJ8qUsTGoePKAK4jQqWBwtYa6OxzYFzA1uK9p17LClj1QjccawzKVZ4UnNvSpU5g
+BHGD6twyZ9vUjNEG9lrYi0+sS18g+DHe7Wk1cRyeHPKtyo0N5gtWKQVXV+3Q5HrFajIqCmkIWI5
P3y8UmtXpI43WbaTZGzvTg7dCFmELmPsPOfkt77lWlIcrUnxVjGQFHaG3daDpaSCjQ7lnLzM90zA
t/br3M3Cy3t276VxNzLIzU+LigLOs3Z5k6bfLS08jt9fXyJBJsDeSxVSJC3ZkiMWNvvqR9cDKd2N
vLl3Kpdl4QXC2JWngqpIWujScOC7v3fSoPSP3W0MS/M8WpWnwh2fp9g/m5Ru6pLCNpDKGxCNbIHc
zhDjSDEQMC2ueJoyHrwdMjGfdTAbL+AbfKU/0UmFqYTCQnFJsx+K5xofV0UKHQXHj8SHXv04RErP
nuQMIvvFXbId7MJuZA4OmucYe99JAhoj25dc0S3HArxO7KwyjMtjwIE8dk8/EElTszOdPplbCzkI
KEnBhPBqO2olZPH1KHXgFJJrL6GWBwb/CQpmOIJGD9jKXdiZH1a+FOH2N0OXArrtac0SOnEzalWD
KYlUoREG5xohHmZBqyjzoJSchxw36DHiJFXMF83A7lTeaachu35+I+WD7QDQQBhTLCysHvlgA5ts
ZxYcsP5ddHPr/F+6F5IEDFp9O1LBgbz8Ys4R8+BvjFC8DWcQz2E3eAyZQqPVukn339sNSzpuTzJp
n4NSloEKfxiqa/LBYtmBWc1aw2Iusrmwv+I4SdgVMTjyANNos3ibjFPq/3IdrjdhrI1EWWAQVfLj
FLyq3DOeuA7CgvovQdh67ZZ9/tU3eaW6rtOfG7yfKaNKPDETdQ5clevYaEVCY4uEjbVoZFtuqQDN
Zc1aYWVv3jxLYZT3vGeRXAxwoARG1x4AKvNlHM+60y/kQhZWSwkHt15fiyknB1299ExEs+/R0Z57
3occ6FwGWO3PPEJAet5zgZG/XIHzEDVroRYpBNP+QMxoEGtLrwc/oyHWt84Vo8Ehe0p5Rx060V3a
GZBKPKY20C5oHkFbBIFQFUP8UbRoZhbUjvxtlKX+OysOHvVsxGkYOrIX7ebzLR2HXJTMVuE2UzhB
3O9oKtxw6p+4Mu3q/hQH5ZiUm9WqxKwO1K7gHscNMMEAPi/Lzl5cCKuNPtn48FU7ejX9tnxdsDQR
hpV/kxDZEqdnXh75UXAPENBXud88Zw/MBfB/FCDN6q1b2YJQy5kOxF12Jhtbc8cO38rmGjZCheZP
sOAm6hbbumYlKAnGIRi3g4UemiNn2BFSuoKWHSRQba7cjFAkH+uZFlwquAZDzs57uRz+OINo9T6j
dvVYqs9+Ybh/N617+8V468A6hQrB3yZILD9oEmOu7Tzn7S1ge33GrTY6vIXuhNYOa3FQMygqh3YR
a2BgqY8h/5HHUCyT+0IwlDU9bKJ5breCgnk19kxkr6V5kf4OiiNHo2mBX8kkJSInHWoba9ZAE30Q
oUP1AXOCZpNGln5f4kwfZDcqfYom7ktZsueEvH+bNOhacRjaUIqHdfj8XQGwlmWfYpCeBRaqsCq1
980HbNWeejSP4et5w0uSRMius81n88jFVFLFMjTIpqvNudedoGoSTYl6cQWhywMJPBpJtk2iZmut
w4ZRdo8cngAGT6yRf4cnTq5EJQvoBBNXhWv1MJGuTprCQSDfjOvHa7qYnufrtH3bcs+SH7IIgxgy
M7HAo910RVcMSYdX+1nVI9goZJDn30ZmRDwd69XUSMzZyDlLpZXb3ThKsxjypMIB/cqLHRKYk3tT
loPtuOT8Gssx8ea5hQus5a2SYszNW8xx+3a6cLhDi0qmz8x5sgV2+66EdeXtWt/AFBU9spcM0sCC
SDUprotU/BPQganQDC/8O7eOZqHPtrdN60kXt0HIYV2R76c1509Qom9MhwiVav9uK1oMusBGjNJs
GLuMlzFMTgfpCYansieZyf62fpTN6mGELN12Y2GbEyRWyv9a+GPRia+vRVkDlG1YOp8csielIN+W
A0H+JA1dhODumMAMCPPJFV/psj4mKZZvc38ImVBsGZA4AwMxT3F46cTZvUTDAxPrgs9+9w8xF2Ec
JvMIAAIBT6Iog2LFQgUu4z3Oa80Put9cLGVlOQvN9g4scJMedceOUydMezcymwpGk0W2i2jzoXff
mhHUhdgr0ybPiocqwXvnzaGvegiMeAl2zuR36RqK+0zUx145BqTALwuEtkzpSys9Y/usTMs4kkcS
odnAcNQm3Bz2G6SAVYTU3mA0Uh4NVUcxGhDtPxVL4PRIcMvzB81dY4ht1IbnPxE5EIPxh100H7Tc
SGl1lWpuEXvKKSp+EIYXE0ZVfvQL+F2y3NTEv+76hisGUnfcN4vaVm8OroYe/c4W86LOjrjrX/5u
webQMRCgfEJcCb0INpXi0Wx43UMbGBEMgNavNRwpvanyxZryndyy3veBDqzW7zzh3kPrO72wJ7y4
xk947wdBX8t8PFrOogzRaLyFdcVjwTulHh1B6jgG/PJ6dKvlb3syXIv7EAbiTSF+6BZ5aqdOq7dl
26iafMP9qoU1emE19FBg1IU9cv9bWRoVWoo509BWmV4jcrt7PhokcOdOng8YmeoS5v89Fe0KLlbS
f3sdRIbvbWV1xzmvKHWZphp6tCwbgdbOWym+/ChxYJTPP1PAcW63y8KV3oQJg1oeRasSTchDt1YD
jkSYXrKQfLsqaNv5utlFZYasBpVPwzshMt53Do/9H30UwSKazXQzrSnKB8x1KtzJWiVQM/O0a7aa
VgoTbYioqYt/xXi4KSS8aKHBBCVgs1RkbldB0z+nYAipVJE9bJLSt4JQQR0gVVaL3ezq07DEyDoG
rq8ZLkGSQkJ8BhjouAc3MTUWij7aPsCZJ42r8NApPfWNWix7/paExI80QXjTPcXHpVqKGG3xCumA
3EVgrHjNfRzhwZgqI1nTvnYmzAB4mPt4OWOiY/Pa1V1PTwmTKkjFvBM8C3Xz/p+PoH4hILxtevAA
EN5zY76f6kYYENbhorU2yftk+Gf5cL+ROTbGFMyRL+UoquLGtyZ/Eyv2/ORAQKyfNeCj6zAAFIv5
zvb++9pa8NbHq7+G32vaewZRHzMY6c3ls0VWbYj5r9Zs5BDljO7TGAphMmHH0M8ql5dz7Gin/LF7
Dq1i48j/dA5qMzvQzvO7Viaz8ePOAnIUB3/zo3sEjxxF//QvFIDvsFHZdDh6VBCF2AjmltFwKxkE
ErNnSDwjOtt0N0Rsy1GuWc4NnclQYGXlHoPB7B5SzLbcm38WxZ0qEKLPimu6LbRozbashKMSiKGn
iHDcVkPPrM++/2LJDqzwn+Pe3zLludSGXZD5/wq+yeTKBQAKyNsBPjjYP39uDJLPigRIFEpvGHq8
kk+z4bPHGN1EIGmujJFHihCmOoZBsveCLVjylAGoyMwc4ym2Kw201qNjPdRzXwuuFFpql6buGKix
0hVQ/eGwlTKP8BbOBvYW9o9/W7eRQ+I31oZ4V7ZkZKQDEca7BAI0N6Ek+uUhx2ui+eOrG9PqrRqR
CDhvsy5iDHzjuIjr5t/K7ubyGp5+cS2/xSN/0lTYjkyKsrJmGWvcxDV99E4j+u9NCI+2z/s//QHJ
MTojmB55DeJcNBpCTpCrOehC1W8WoiAf9STi2XyOqmHVG8XX9VCfP0gJ0CyztXbpkFjOnwY0w7tY
7/ZLfysJvKXsBluRxy/4yJBB/2FFNWQiRQre8jp2nHu3NQG7Z36AuFKmxj1ApOt2Q2B/zk6S1bfM
ts+vCD3NTxhLnqKhGOCYIKiifU7aEfxIiDY4Aai5Z1KExd+0A90GXi/7pt7N0NCgwt6V7UaKHUjN
D3DiXDnZY0DksHPaDAzFCTJNncRg2Wn+aOJ13YaT0xnbY2XHt+dsG/7LRJbKr4m8sck0uOrje+z/
SYiEMKxoLCExGSAauPgVXZWTJFO5IljxIr3KcorV3O0lrpE9NlgqvPJXygZhdqd/YwIFTK3lV1O8
V3EMztseYoMnIYvD+cnrrNWXopNMDZfMvuZSecHqHhkYuMAA2a9GvHucNdbI7YrDy/Iy16CniZnj
IkikdhcgHtseI+G+Xcyvmrs1Pw0B/1WgKtz8lQQJ0eCeVG8h12aFF0Ltmg24opf/Xxoj852CGHY3
Wtsz0p/Oh4xto7SPXLVqYXBDtqLk3p6kkjjjMqF6rxkGVRpuZw3q81TRPfBTd4x/kot1lopfWS76
2HshCVePQuUly+fBpX3s3ejsMbtUJK2bn3eAtCiYIGHVdNJANEIaSmowxKCiiTjoAazjQTMLIeva
JGB9A9S0xm6OSdZ3IA48nbydJ94bthXYa+9Xn/W1dQshsDDCi17GYpxH5Yjoy0YCAsXDtLvMotoa
way2VyCRgzuAxetdMgvRLhtJaA/zBURQ234xtHRtnEJyDJQenDoORUZFqKXmDOAoNp7M4gIgkT+J
CXCm0S4BX2OeRfu7scEJRKPcNufmgUR5OQb/FR9VTHI74ysHwTCsZcJ9B5f9TwmWkMfV/QNC7xLP
ZH3fCjbPyVCugGWXj217RyVBmbDTX+oQwOFGYOHA0gPvC70g4gzOclSZAINbE3x0Vv0oCAQ2UN+3
ekP53Zbed6I/k+m3+XR+nvtplI2j91+wYxzKCEuCGUMt1pi9qWANmYcdG+sJAf1LO5D+G/9324hB
XC1GR93RY1ro9iP4+MLhlJH5wNRaVN+p7sxB+eZsT3wBhAEALrMQ3t8+hEFSWYGESwHj/auWXZGy
zl9m4Z1t2D262ba94lTew4AUnnutXYPzVJ47zO/unpX8inPUoMBqyyj5wjJlK6T3zR2ssnE6IziC
OJVn1Isv57jbmDAunKbj5yP0ezmOrNSrDtNdt2RQLMfTZneCepbbeStFSBdp+f5Z+amIN2TdosTX
FV/OV/zwS3jv1MvYcN3wP+UvfIlYgxbudx7OqToQg9PV9Dpy8g8rSmk3nbtN7lyxk88cxdXTdHE5
AfcX6El4Bnvse1dBo4PmAMrA5PQ/72GIt6aWRHCc44lw3CxIF1QFKncexNACct0CNywL9PFxNzUK
a84X8rNnTNQEnfJ1hWiOKnobtpD1oIJaf/MMeWEObvrqNHpkoBK7CoS9kFkCL0mqg2a9+znLdS8E
slRqIKJ/a8FEiu0GPFF/4rdwSlkZCQDyCqr3LFlZEsz03iQA6Y84HEPnyvmYWxP07aWfebPZIpX4
1zS3kXIKYg5jfzIBVpltHCywK53yyD8CPqrLSbxzzTKSki7QsWlV9T0wzjSLJHEiCg/7pfF56UUT
rI248nDS5ILeoBGAdCNJynKb+qfrgJL402V09z+xHry78sKpikGq/dx2smJzC/iOnAt4Dh347kfX
YsXhVthy4jZpUTMpwg/OaMvMvHFeO+iuC95CzCfycWlkVC5Lvy+2hA1hY199MREGgodKyDSK49ff
9UfdJ2W2aoKnfFTGtM6OcJP3XbR3/7nXyeb8IIQTBpmLINHuilGQ0DwoN+GBZZhCWV7Buf2STdYy
BvuBZCSkQnG9YhLBWV21V001NKXzN0CE/6YhBTwdPRRJ+d2XW6SfCbXwgJRse9kkqYgRWegLGOpS
WU5E6jbplvTfs5TlS1QDO88Mudhbb22tQQ12cChHU/c+jal+vmJGHbVys9bsObqhp9JGkwdFwR+0
6bq/SeKondIuQ9VQQlk0+abVO/yD+MWD5myZjNEWPPHvqo0/NeadQMstaE0jy82iyl6I6VplnM1m
wXgMOdch0sOsNOirkKm2cWPOusnGpDgkD5r+Fq8BOCmrwYcF8/otcVWmIqVKum493XmefAuGCRbn
qkrVw/75jZPjy4Un5iUWt1saNjQ6NezSmwcp7h4hhZl61lMEDAeg3MZ0GiT1HCUT3fUYDDXjJgFc
edUT2R/gNcFUroJ+2+kzxuEVncqdoGw+rVZnlym6V34shFUm7Dk9LG+9iZtGTAwykriOZWxYGlBO
MLWkN3nC/TLQbCqjNq8s/EvJEtcx1rubBjO5+cGgZZYFdQgGVg2LIffWEORu4Vrf5Y+xK9TD2Cx3
9jdaOfL1ax99i5aP3R1VB0ITCbBvlWzrrF9EDgt9rQZI0ZhscT6zdyMy7KBv16eX8x6gUXaKLjx8
6FdzEczIBvBvwtMdCk2HQ9XVVmZ8LRd5Ygjknx7ayxKjHaAhLMirRdKnKJnVdF6ze7q/2kJbMDJ9
3S/HqsfsCbRrn79YnO/QYrLpsP1JmrdLKjMPxH0uhCMNyNAdLcJSlCns6csAewUu46H1mzy16m9c
Q/wkRYXJTKyvaLeFkO4pgSpO8FEl+bSSEZv9jANXwtCBAKVAgsFHdiFJVZ1NelKBItqz3MH8vApS
WLxOxZDPNAn6LK2t2G5mwPc2tNivSCCyrkVHmEP9gGL/ddSSkHiAonZEv6MfNU16bWUqFwAV27p3
KwXI18A1Qgz5wFB9xCJsNjaK0ICimgAAJc7cd9kcUto8aQ1U+MClViCQDQJiiX2e8odphkKQqZ60
9nHJ3A906/MgJUfNgP4md/v+Pg8SwWA/gqEo6Uoj1zI+lDMU76F9TkOAhNa18Enerw0gEDr3y6Te
YYqn9Eb8LT5m4u4NAUZeWfVN+oGbQ7UTFeHDV9F9JwRsf6v5DpKSaCM2W5SXrVilv1cNhXJ8Lw3o
fur/iFiVWAVJNI6OZkbGH2ez+d6MdNc0zF9guhz1ihure9wm7GTtJkm4OU9l5TYYJColYm0AkwR0
o78o3k2GSLmgW4kLTqt7CiCcx5ddjukDmyAidPmwOUElIzE9O1MISj2nUc0hB8k608PqzMVgxg00
KmwT/6tHQvth4yrfJuybVaiMS7SGRbhqa368Vuc1p97TamBOuLNFtC3LXwqA2tJ5rZAG/Zx1MIf/
e0HfSYZaI1QoxD59SF7+qyUyVxzWbvMcEzb9uCWun934UMAK8/Uzk1+/Thl/9es8/y5I6Za/Qeo9
Dz3pcKds1v4S4orhhpWIP/B5BlbxBjhD/qA/QfoSSI0R2E/ElTj51re4Otf6+WrTY1dN4VAg9FFN
m4v+zIJcXNfCBVL73S70u3rH5jfrQIArw9VdZSYpL+RdUI8U0VV/ys6Xhk1d9W6vmfss8J/sb43J
xsfFgTWdNEvSQCCCPE5N6tr3fLLSzFtoMm4uF9kI8i1IwL8VrdBhf0LCpzUe44F0vQYQJRTdtGK1
1/8ISwXWu+9dXnZWuxB8pkK6ftKRtYq6uOWWBzJm8p9fyR9grr0lU+dJnSH1S1FSgL2+igJEgLBj
fnqz8EBqcBtRPPYonOIJGBFF7pZWxE0ONwRfGpJYK7/mmVR0AdVoodN3dOf5bkD+nl8LePJQlyK7
vuI6sOcFczzgMu2Hp9igwBA/gZ3EXF3MD/8YSv+Yzq0jvsYWHEIChP3YFhh3q8TpfwmXUF3hvi3B
YqIGQJj+pbU9BmQFX7lFvPYJ2PrYPC0DPRf22U0iheAUg01GS2ucHkQKXpGAT6OsFiqOI4nyna+Y
1YDR6qU2AfVSB6foLaCFNCarbFWTir/S3usMJAFf/x/+m0v+coIMQKn0+/K/sb6I/BMlClU5hyow
jAKqaXydvK8FBlRDe446vvrkkRjvLzD8DE3Cb2iaxTDrCAD9zapQNqJRMrD/7FZHDPkxgTvtwY5F
wQK8YtrTo+ay8nQ1bmr/y8+n2xwqfjSDDe8Q2cRZoRodV6e7o/gO6GLd7UACy3JZngvQ80XDQ61a
gkAaFLz3+UW+3x/42EIzSOZtXSRp7xZp9hd+J0olbLVnGyKR2GWnyFaCKOZa6ox/GPLdZcJx1/up
JMEy/fpdMpkdGjYCz5y1BmwxMCZbTWyRDEfjIxxrdp+Ia+wJijy/1KdCVigTJWL+kgJX9onX+dw/
HGY48PIw5o5rwJ0C6Mhi483lvN6WGVhmA1DD4aPiIt5hh9oju8dGZQF7XBPCdwkwiPTc+8bdw+8c
eAlecvso1NsSv5rXlnG59DwCtUOL1J9js5F73jq7piKRDKqGESKOMup/TFrCUuyNWUse8+3GxzPz
Ad+IqH+HMNIbCAaf11R0sI8ah+AGVwAeVQ79V2jN1EQ1sfuoYfcmbi+mWSKm+KexqeRpysaNQZSh
I3FU2QPYtSCDdfFBthp25CxnW6cA5RsPgfTZC6rujDaka3yLiVW4rCzhdBOPJaISV6VSapqdkKWj
04ZMn67nCzx+2aIbd1zaoiJPqaxMy0lkJTA3AeVdOMr7OYpi+aI8WIwU5hMldbJ7X7Z/Id/ku1kG
AfOU3mziyB8pt8+XdDr5briicd5Db2HsFJ9xu268NwzOG/F+BqGo73FfKsbBlt1z0Md7kLBwHenx
yR3icMGIgTXnzmhA0+SwNUW78j2UL6gzimdvXTzPkY6bnS6dMLhkxf7BQKSFwIR8nBnrbBApcD/T
F78OhF2ftOeLAR71aBiF5hKi4K1GfQaYMAOfyFE1sEkuQKqyAPFXcSG6q4h3BYmjk7l8tjdJfmOb
M04SQt/CnxKnApJwnGwg4Dq39CZilA2gd0BNE+669KWrIYUGOEouRTAqfgDIE9Xv1wj33UuEHgfZ
puo90V15LIuQ8B/YesYve5jMB6F8qSBXRKcGmCKAjQKgcQhJtFBe2Ud87vy/rgGaoiq1RG2HWmVh
O038nWm42xzYeAMix3X1oXayOEAnWtmU84bLZAi/djnSmroyvSqefxh7cMuBOSsezQtLsNZKhld7
5QHUkEnbcAyQgIuP3whqx3bEb3hXhBNs4JCX/n/klwZ1Fq286m6wpL1hBSYW+M3zY1LqQ6b6VG3y
lXbxtBjZm30iqxrYj6JpOBYYuC1+TW0Y5bDz5LIYi9gAC5/nFMJFJ5OLfkoqcSh0J5HCjOB0QXMn
oyP/GbpZPepXamjN5u0ZLTl0Swn8TtIeyPHMyIKHd++xXdixTed80AjaaIqdfD3SY9ZI+LkMWLRC
1adL8+TnzFKitInH1rWA4jMdeCKm9dqB4+D3VUoEl7E2+DgLjvBgQ2RIh5sLZbxP9ozK3SDtgkHP
XVrBbSrB2PmmRFkL8UUVZnahtEIuWnQtxdKqOsf1evr5y1WQWFmjiTCiLSiOcqUkgvAlxwWOP7D/
ajqMGPD/vXpMxUgQJq3vtYqg+8/9IMX+EZeVzxvEBvIDHPVerarCijPYnaGULEgydbJg2ebeBZMe
a46TItVYccpPcn9hjx4zhFkbk3GUgeX2x66PV0NmnlZXrLemvuqQtriAwNw4YaBRYzkpd/gi7fzQ
b4JAqmNJf6hAb+dM+LtE0wMTGiV5Vr9MBEk52mpNC2Yp0Z4u53Luk7Z3jPn08fcYV8nD0ogv28ds
tkw5DQHNXOSdylMbT4Bjhbs3GYFMRhP1rQVDXw/ZstgDpyYHU3ZvoV7Z4vaMIx0Y7Cy2Kz0XRxwZ
mpjsRMe6qaBof87ZxwCtaqcKVi18TgVYogTeyDl/WFt2jlULA/vDFRuI2O1y9ivHX+olIienOTUy
LSAsmv3aCE4XuRLcFIuEF+7sWnnHEPqCDwQ6Z+MiP2nDSCYjTEZonlHdPkQ3bJk0U1HhiYUT3yqn
NZetBAzvAKEqafbK2kvDq/Z7ZeKamNfaFIlpqCfL/PaqFhYq5RDD320b/0ma/WEfpAGYc3c+xJ7u
GTUQoWfrTpJlvYOeAWZB1t6e3QFYDBtYOp0+65AmlEJXMX7Ob+NHYPW8yeHxS7ozir8fCQjtetBZ
aC00vlFJoRnOwhEJ4PXubyTu82Gsom2v5g2fnwKPtoirRREB6eeU6M/4Jh6w4qTpm6AcrZGdbjOV
sbYBh4NWN2IcpcdutmgMTtnKO5yL/okCTZvye3vtu7IKcshospWo7oI06HAW24DHOhDGTyHYrWbM
GwNdo7HehCoTFxtYfw9BSKU6A0LFuuqH5SNPJ4s+mClr5z3DVzrx8W1YdD7104XKioAS6BS1xPew
0CNr7AmCKGANbUWNNCzyTF3zOB0paYqgyTc+R2/h5U9COdYUgjy7VTf4zQYQeDtB1XMeW/hzoJBz
OqLKMvcVC1rbF/1g/a8n6+ZbB2zlTxHRdjW67dHM97UjchmDhWLXRrJ+HrfCGs6wZwMuhLr5Durd
Xkd8ROKtNeceeanj2rtJhefyImYCeDj+wg9EJ2fen7pqb6ubB3Oi9M2PX2bp+2bnWUmd8/8GNbKY
GQpI6w+HyGAGMpbrbVJJANy4/f78z4ZjlKjixBOprMe2LvyJ8gruJttjy5R5tqzqsatLCuBFc4P5
GLTcgvY+CxgCTd6cshNL6mXypzN48VHgx5qnj5s9bPBr4Sbbks6QR+E+fBswfvtqIdxcJV1u3Q+V
U1YlWcy883fs2NqzO2/WIMSNhCQEALlLzlsaQVeI0JSmvNJDlC4Ft6XprJzvUcvM8hv4OuZ5Tcet
sVmN2JQT7BKImVZXIwmRfoJGnYiTGZCBdjw4smX6u+6dBKPm6KYk1W/JBfaQDivsJydH3egHD3N1
a65r+p6RbAkLcoVuznx/IwNcQVJZGGh4uu3dndTwmIjOizQKp1/5CM4rp3LfcrMTZoBZeGq8IpM5
eHDeytYqVvZHjVN+5urVx97jupJhYMrAVJ93QbFEfFiPMExQzjx8JukWTqm6bPT01OOJ/F07vYEg
ZjW3XgAApgB0x9fcq+vn/p6JmpkrLCDykXiJ/VN83LMp6qI6DqZRSRBUrfcBTtUZ+jZVDq4EVTyE
pbYpVmr7/zeXhJBSLP0RvDapx9llMhN8mrOW6ADcAj2rs5rhi+Vt2oRf71OrpFEp5ewpGI2VTdew
oGHfT/oNNdZbniZZ/JI1N8kZn8bReU+ol/O5ZuAY9Dkxy4Q2tXd3AePUy0OWYjphkRU3Lnzv3/RB
gGKcM28yPK7hu6IbdKSxR3sHgh9TsrbtcBMVGf8YrO7PLigtXKYSJWFaOrq9DsOrFkQbkEm1kea3
Yo5uSb/J4pnRIrX/ajGMyKbl3NEvJyaoC39iVYJiHTl1TIKiBRKg4u0Kq04QJvreYXUzdPEv9HwY
tbyXOZQhK5J6yM81/antbrymZo+kh+8e0slX7RGwtGj3iMh1cCyHGdxQj/2XSV+B0hK01lrAzQ6d
HbEtzSdaH4OXNb4qHnwu7FCVxTr5I08NTnIRtYyYLM4e4syBdyMiJI/3632TgL3kNj1o89S4bjqt
ZcLYANFFhJ8v9f5CSQlYtLW1VFuSOroVyP+nR0g2xDtJg8n//0yrzdgRvBJvdNg5PBmRvAVOuDfz
3BHVtZnS04Pqkca8AhuH2Lc2AL/msqFVAfDqrou94uUJ8YIsnpDBLi4KT2kFdCsr7s9VbEksKKTb
o5FbdmybImueA4D6uidRyG5HPaLyFxCe+W+Lah1fLb/czIvi8Rr8Yq7YDTJXM0T0CENxnsPGCU4w
beX7TgnoiOJfwBgLr4bB0hF9JIvM+zF1fPQzicGMz77SRwu25hv31mId1oKVjyq0VSG9hBKkzanW
MLXgcvfCa08wgz4ZFjn8xgzTKONLAGU/v3D2U69CWEfH36NqeHUIev+qynxFdeBThdJp/XFmIndy
Ppzw9tVv3wbSflUR13HTSZ1kesndbkKJW3bAhoMxTXyc/f5GFWt5qGB+hUXOJmMMvG2A7zKUkOsB
Oxq2LGWy121Z+hIyESd+Dqd9NRiQcsR1N6Rn/EbVGf/LVUKknWYhxr+Mo8knbD4Xwas6qS7ZqraP
5erAjINYA+vHV87n6UpznX5oBfPSLOEnnTM8nXxEDEfWAQ/G40DMYpeb4tlhYAICDovCILc6F6OY
DO6gP0MgavooVoGp3Bl83jZRaO6asyonHkVGpckjkggqiTZa1BqW1NFPAUMxljbRXgz/Fqlv2zDA
tyt8s1J72UaxRD0ywVaD66Lygp3k1Mi+5B6d3jQherQa8uB4oJx+Q8xSGstZiQm0VuJEaofIWzFJ
Q3xkYlH7gyQgUVYu3+J7c6cqXdAh3G4cjGpp0OD81yNp+6WfuFuUvMe35p8IvZBYXwhyOMRb5Ky4
veax7oy3tgX7TTt83uPMHnVv5OL/mkqj3lyK627CJn/SUEqVDPI6qrHswdPjxxtO0u1u2LV9fqOd
aQpxsntdQVsx8+0zKen2pOXaD/mhBkH9fCsVaR2K5cSXWjlJ68z6hQRvPXPuZ35Z0fy44YsgOCtu
3FWVFlnrVpdmGv3fDWB7ZEMCNCIjQeX9eYwxcfW9v992GjFzqcoq20ar4Rm8k0nHgcl+rwUMI99S
AwRQY5h5uv5JHKzGfjua1sGSSluXpkDdZM3P9eCydFfLzcbxN1F8OTLU1NAVxOG7uSVtFbnjFJiS
qt4L2kDIh/nx/j15aEi42PhQg6ciPdXxhuiRzOBWM2hhpAWvz8x10JJUqn8ypEelKHUYvwBkCCIQ
OkoEe62aweRxgqIfpXJdNPqUYAkHZBT6derQFFLrriECIeCXvdTsElUEzyszizep7dMiPpvMMF+2
JcBDRANgBePh/b+0TWK6/WJA1Z6tc+451EBFu417rd+rxf5+9R5S9jG9oQwcairFzxiZ+CCXsOQh
bPZGmgUiv7LXa5ub/5VPK490Qn0x6SSUTKujKmlQzex3IcIY/+OE8yu6Dy0kYsig+xq8AujibF1q
+06YtX+YwWaeOWpZWjhk2ocQGF0+JiEMszt62enYALceEbMwc++jN7PoI1oBeoCBKicKLOsjvmAT
OCE2dFZ//I8AJ13hbKnEbJkvHIkqk1GMBuSO+rOS0aAQH7lc0DegpS1FsDFkvBR5/uXQzJhGgfX3
pa2jHFURogNZWDQeUo3i+Kl5VxOF1wmTsPW/Q1fS4PTfZvQNAYXuFRKQgIJDw1SKNDyvBd+TbSGz
mHbtiCUNRzuVSfiu86vXq9KhEeJZYmIyh9b/0WQvUe4IIic0X7uOZplHCKmHk7KwtkxmC+mheom+
fpPN3jFLKW5evRjvw/1Ri3cBk0v5dOjaYeCXrbhQaMOEpyyVss0CygQx5Si94RVqeSkRb+KNoLiG
XwUAaBdShnClsmrsub/A05Nd6/V8APeoukh+pWQy7b3FzvQ/YWn5n+wFFT6427LBLhel58vUTF6M
/9h8v2ndp7ms2jl2QBZUUy3merSVlYitbRQTohtcRHMkeEaADcLnx+EOGg2UmpzjN66O/XqJNtrB
3hhtHW6jnPBlIk5X2ZiAEt1z9a9kFCm4YTgtRbyCR77uI46bJ1gy/6o0Ysh+YrYzRJDsp209Yhll
GA5ynCk0vc0n+7bg+eCSwmqEu2eJppVJlt2GmrwBmWwED5yFEdp94rUaKaeYQxrVR0gxqEVbHPYc
tITCDLGamgknNc3G93VITfaLH12UPgKumOH2KM6Ze4ZoJqiLVftHcEieEWvXscsh/f8zlHGJHjZ0
xEst0V3Xbl6Bq3WoL6Hf2L4lihkeN48Ed5wYVNmp2K4+DID53gB+hd6NWnG3sRuNXd4MPXB3RBUV
oTNIo7PoV3UIsED8ejKJ4c3W6munlmCbv2d4ng50533K1NoyLerp5OMDO7JyGE91ULFa/7We/p5p
rWlZ2nDzaGAMgnbIj0LO6cYqjLlF/4TuwH5VOj9bcfdvyM0f/SafLYZab8ma0Ei5RezkjTWZvjN5
MJNH99Kbvqmuf8PosGP48y4L88tpqwqsn94zM4xlA3xESPPBFnyN6nVowoR+AJkIbMbAZZyXpWNl
ApTIQITDexHJMv8+v45PHbVeF4Enf0OZpxq2R4IR+JbWPHGvyblIhTv+VF+DvWy8J8KdtNLguLCn
7yzW0yd/CVAKK+1f8gpylRBHiWYjMgz3NC8vZotNI6tkM4LB914jQuKAkLoa211vAf9fl8/Xuk7o
CRUgDGdHn/v3w8UVtc2G+dNxJi7GDq25v8H53xnD0afFWNKg12xR8cuyBPSymf+2lkRY0S5wszrf
V+gtP6tvlrmii5wfszTJwjjdcERdTjeGxLduJfdFHl/qwnrnMw8HQH0VXu3mCiuwa2nYbw9W3nEa
6M3mGCTF6QBjO7VrHk/CvqjrgaJCPtnvkf0etIwr2ugXVlkw+8cJ8Y9I6/y3K0AEpMPBXBRnkNkv
YltVmhkPTRnZH701km58VY8o1xVcEsfXLUWUAhvJerkoq0kRF9GMzOjVBxlUeB1o0C5BX1bCjSMU
Rr0Kue6lZiyDNxIZDqRouyYTtvwCDOYOMA0KUG10Y9aEPkRqfZBEjCp2IUtSmiIXF71F83pkuZV8
JnGBFMn1HKbIxunvU4mGWdp/fZYt+ib5xf/z9wGh+qUiuBFTk4UK8MesEUj3L8XZVtvn/leBxZ5B
TyMVqnocHF5H6gkxZ+4geqswX8qkd+Zo4nQ5w43UnUEaHakxV8jSOhqyzdt0WGPZp9OANJvzm30D
PWoanHUuYT6QPkB3YjiiU/L9qtVO8o6mmhmqvEOti6BfBAwzsRnJETO8+Dh7ZJyLGF372cKoD4lo
lsw8ndgurg1HmekLK9S3G4dY1vrnxvgo6ySi+K1PzltJulbO+lQUfcjYOBYqdApYXPHzMIefkygN
iDuImo5sUpCi7hYSfKQrpNmWBp+DLOp7fJI56UzA4RbVrFk6qIbx7BGSl7jZ6lBl4AdjO4DyxrlQ
3C2I0MqNe3YXL/KYYzvdaMe9J4KI78eBXQirYVsz2V8fYBY0EfhWG+6TZ/Uh3jAFykt7M+WaiTio
olInNPhyKshJ+zbQL+xTy6pK5C2lk08OPXuCsX824QOYe1654Dryj/I2Mdgd2wc0DWTcx0f2Gya5
nRwYn4bSB6LQ4eHuj/gO+hNEjMR1VHTvmUZplplCAVe/Uvc2iWCxf/RusXdWZLsoDGeE3Fq2fwLI
n1YFKnhmm7GJQxIuC3/uS3DWab7yFW4ccQNpZRTNGcnJw5HeN0DSZyx2ED/JlV2MBXFr8ToGRgOb
VEjKzIT88S/Z9DlRS6CWN4C7WI5t37FurGyoE8WzuEUa5+VSoJ5YMyddGw3O6uyq6bBcIZtwdSB5
bKt5pmM8Fe/AfpfoiOYdcjl0O+HiZC3vCYcJAMPuYXUy5wdfa84isAsiDLtBdGEWSIj+c384FDOc
LJ89+NYWP4kFIZzDhiaaYEzMMQgp9P+tWWI+sYAd4pcf0Do3HpR8g2bIshg9hViAyV/Cs7l//XUm
wD10xTBtDH9GT2T+6IsKZW6Dg6iVGFfh+uv9TUt3JM2gMEl2zAshQb5SZzB+ZBFgM5O4Tx+X20pp
GBuo9kdzta8s5xDFxBzUc24bPDmqYsc2V/PNlHBXt14atucR4r1dgEYHG69gS7z9jvWXfTyfK9v0
d0w3sYOcUXMvrdzfn+CaNE41t/KHCaB8H/LCzZ6gkbOWFcd5reRzqakPV27APGQqdYyo9uoaAL6+
jwg83M1Yxw43hJNjiGwFxx6Sm2qPVDg6KCIwe1ijO1zvU3o6q6U5R/PFJH4t0MJ+0BE6NzLgt6ZH
jW8OdQMlGHSKLT9onjm/6iLDSNDD5qYJxExnAqmOj3ENt2XYkRJ/wwWU5phWVc9puR0CTYVK+Ot0
5o19qOotpJL8t9Z0u/kzOn5V9fOxUkXlQDQLT3hDAYKw8mVfRzlXG5Ri+KkpdsZShPPqZEhpksRz
ZSpgPcMSIgi1ZVz6J6hrtYRTsWAlAm27QwpnNLEsG41FPytbcCmgmx3oEykqdI/lnpVWzbAxbpN7
7y+txYLD6kvyzLkIrFqPkpXEPU4Hb7Gzcakx0KVsiz9xgfyYYnjhXzwbdtXfuOX1r3Y84ojCMYpI
kVanumVcsp0n72yNxLhPDuvXIiothDsSUrlBFdV78kbiruIMY3mzI5+ONScHyWgm4vvyh/l1R7Qm
yfe+mTm2EJgLusznuRGqs/1m3e0c7TmFJMzkQ+I9NUyjaSLJqeH3vMm03ffcThfH+GUlyp3pjzqR
1DaJd6E/40AUdMBVGfIKMRFlY8MknCiBh9Ze6kKhYGawj3t/E2d/KKbOAGQ9YgSiqY+wTRa7SI+I
ylVGeqZfGNzyVbEpLaz8ZRGV+zC4PM2Cr47Iy3zu5XZmwMKSszhzy+EGVrxWDhG+5LUm5sKl2RdL
DB94vZQAtX+a2/W2X3DArw1f6H0q90eUxI/b1FMgViNyREeM3mFTqMaFUp/N6xNvMC7O903zGbmP
mrZmiUGwKwipIujvlf6KHr9gKxGfJ+SVx74MVetWA4CC1SNM3g5/Nu5OuiTr5qHXObzFFOrI765G
RNYSYqkxbXaHYWylbMFxLWiwFEkjpPivlywdV+Ib80m4WKh4acm881xleOstXbq+D2yawU/SZ5D+
XalkORerO6o9MINlZGZ48VnqDkYyMoPZ/qoWOKDRQYweWldUy9VkxZQmF7Mj4nz0UjoK1nBspQuX
FnDlqZa+GtwMPz6LUHyNm1w9vRrOnh68hIoeIxK/v6OAIWT6nn8E3aAke6SvTizV22/XcfPyRSEK
6ONk36yhMHQ6Y6V8lkl8db2iB+cQURXvvRxOfIONrYSrf62F2VJo1zPnLxWrh5ORbz3m3Tj4rbZ6
UpqtYwxHHkZ+UyIi5LxgEP8HCWwf+tPSFQn17LAg1xhK4jxvjIsGz/F7ZTxu73W4tPLCKpBnWm18
T5M1Luazboz35Z6+tWN0RGgBxolOhLz1eX1yEu7yEv2GXQa4xxYfZqCls5CLhWmMyZ1wW45k/nZc
Uftuaa6fvMnpVF8aKQNcTeNGlBGH8Ia+xSmN3vHdlsZDToVeNaVsQz86ex71OuFovNkxTIz3KHa1
coxitnn3o2bLT50PX9uYDJKFymPzp8sYSlQ/Zo82A9AyPVzbeYHXQTq9J24RMV9dyfj5H05UksPv
vxcQdb5AaOxe+muN5Ix6D6mqzz41LUS+PAPRI0GZYsE6LgxZTS/FC4gzi6VdLYON2waoX1DNzUlS
fihaMPswFvMQccKCMt7gb108t1BzfUS84oDSiawYNl6FS4FMb4moapTgCe2mmXtKKjdpYWF9q64W
h86bI3sZNAa02IuN3V83Zaq8tbmPOub7KfQg5J3mtGofj4IhZlhrCcc9hALH+FnVX/1zw55BydXu
oe10nJ5mHI2h41OetzAva/4V3Mudr5YPrsy9eorxPtmerqJF4PcFlhFkUpAXtVt0QItu/yLCNcb9
r5X5QqeTDkcKYmMoutSybyocnWEkoydd2o79yTuPDqqpcJNEJ+Q4cfWfmxkFDzYs4BPdDAKmn+Cq
ngR6pqL3u5hY2M0d8EInv7n9LwAh45xwb0KY70NqPT7+5LMleDLQNpmtm8FhRBOgradzRHCTQ/G0
jBWPw4f9OlT9JYcwZq36QVcJfEPxIVDlJNhPZLhRUz93HXBcKwK0HF0twE7wvM45Cx/PLaqRBN9Y
FSGsR/SNXfTw+wc3R2AYtuRnH4Ik6pYLnA+q7v6IZQ0/7V9UPbf2LPKwujGCUv1PThQfowNyqQ2x
L3ChsNVIEnbQyhLdRFxkbrHZcE3xQ9eDhYsKBNWcvydNivcmSpPChRAScG6h4Q9V1au9N2iu8kGr
pwHBDwB/RN6D9ShvvxiYU147F82fAAYRas2mB//Ey6TsxiDLhYxnBe9fJQvCgE6fWeV3RQFdUrr+
V2DDOlNwLbuGEgzgfIVeNcF4xVCKzZrnVRd1rt8FSzhFMGaCdQml1rRpT0Tbcsx03GK/JvMGgKkL
z0psuCg5MNx37jz7+SdBMB6I764xWnQSJhzkNW8RL1MgyLvjfbtiu8zzLaP2dPc23i9W9f1Xx43w
EeXv9Ah+5E/44GTAGtJG53fO7gv6P96laICPiDlUHH8lJCWwxRvAjdznHcbllYquVqncYhBtDoaK
BWF5p4M3YetmcI97+EVmz0eiQjGAwknz0Oa8zUZJRYn/DhXj10PpcIZ+Ju/lsA6fpZx7H8lreGoB
J3lIJfPTsptZ7MrZ3MM+Y97+XFOZ0+ayfOliHH88isGWctv5Wsoc4fQaOdGj8dr5Cx5Qnf25/lcy
NBUasB9WKjIYLr8loISPcWurijlps6qmkhbv6L/fBipbuc9asyOztSTuKsC0XEjBbeG3o48YbBmB
g2isK5xP3Y4bloLWofF11bygyiu19oWXsZiE/yz/ayzz98wWPl7SI763+sQSEtkPRlP2W6FhZhJL
U5ujHQVwSebN56BV6v/sPqYZGMft3phNX5x9BEE8KuE1DkgAuKS5uTVsHyVzy59pZia41sWoOPyQ
8r8oKNlXW/Kd6GH4GpnUmxGp7SjfgjymhjLSi7Vhoq+L8vt4lfWK3LHYjKyIhcUxDw6WmnhHRiq0
neAkf/SNU5s/Lx7bcY6l/+4iRWDZiyRFmPnqPzMk8wS1bDN2KgfQGzxYsZjStcY4NWef6yrU7P7b
dnXHo7F4GYVYr60MhBrXjCOjh79KRzduLF+5As7h4CaaFs42O7EfhhKvQJtWhjvvwTimDOp82h5K
LA85PWY1SKFfUS1NwmwKAN1UCaB1vB6lR/PYhWI8fxyF1yohI/2ZEgMu67Pyv7268XrWmc2akslr
VC2hNJdgSBKv6BG29+WF4OA3OBNjUS04wm40yz6J8w2xuTrP3pDX1lx/duRIQeapo21iUrPRyD5d
VgBcDCssKm+Ak2/C9CJkOA/nsEux6fwIeVRqd546s0EYL1sogFC9nXn+LXi5ULOS7Ctq+wkY4TUm
nIghKsEyqKCfXldaeEop3kg1BkxGWBIfBAT0il5lCmGzilf4kWSX2XPiy4rSsEYgdbnua7GkYW/v
BYJyznii+4Sf3vk3rJXnxh4zpmdf7aHEjYTcGir89L3guJydWA5AEw4d2c7aP19mrtnSDKi6wghZ
jeAgRbNSBgFZRXLpVqLN8LebYgpWxqNzWFep9XSBiVw4NZBWI5Tji8QpzcCyNwUVqBmKmW+cPUaY
uCcNRwBdTBkwF0PytCgUK6S1TJivlgwEYmx7Jmm5yqLmFH3nlA+Zf3DA+/8dN/KifFQnK/01uUli
gykGWPl4gSe3NI/bRbWmmK802P2rtOYCrRX4uSylLzq7FVK11K764AuxgIzXdYmbXguhD+p6Kpy5
fWNrMgRhF29AdfDFs0LLeM+RfwFeKOnwFHuQUTKM0scXqjQnAPnrQRuytoRhFYf93uOsaf7hOp/K
PoAXbEyHJpxij7ZIKCrItsWGu6ibBOIGS1hDX/hOo6pAxv6G1VVIYfvoRlpjKYPazbjjCwgoVm6R
OJntkjZEwtzDYOvy5bQyxcPNMitoaXzpIVT2vWEuLaMRRFSiICjuCBqRVUoblJk3XNvk7tYtELsf
km0tbBUi26CgHMJx6n9ZeFLIrYB0CJQ70dLN+hORuU27dM+hpFAlBBN9X60GYw8ffurwr4XygfKY
MJxqlH7q6WilJq6OL7yad+icPqhwCCLNz0czTh7mRUVIgJB35VUlTKro7nGyvrNTGxrc8UgKD7Xf
huQouD11ne85Rvl5WpY/dxlG7KRlnI1a3lhRFCz+5kH2bSZFbZCtV2iLIYP8yeS1E+MbZUut82VB
nkQMSV+VemSVeCpssN4tozt9IDkn81d3hx3eI6T4Dn6iu0GDiV+iz2kQYmA+HyGbDGEvGd2kmELG
AjbT9RbMiCBwHct5oDUpf0NBCglG/TMW8pSYQQuZDGuTrfpE9hIG7W+IaHvpC+l8K8q+DImpIZFN
PnnUUvcGPpjZUl11juDvbGpcG4uN4twoiPuaUaL4HsKpuzBqyO17nlCA+RSO540xkXwYGlcU4jT2
3nqOilfw+Wv+02bw5vQgEiJtvZ+1WuXCPwDdi+zoT01OuivbsH514uck5eLPnph5KANsqSCeiJyO
E5M+ASB85TTu0YxuXQGu8gAojDeA6neBSUHGfplVmrmGqAYjlEx4c/RorqXu2tDnHPca7Gbtfnp1
1qLfGxvmigWe5s5GeMymPHeOraneI9/119twRpy7odUjEzvvHBntHU0wqPbrO+8GEHlu4ZrSfkdi
jIdpz6lNx9PcuhtKj0r8uiKVsIRfAVhORE6AlA7cD7EknMXNBeBLUXlAdLQT4nUEObjLOR6IgA46
f2ERbmAPqDIOE6CTUUbCdDJ1T+4aHjm5FAlLFubvRfcRwXIZ1mbRO3B9yYq3xNJF2oSzgT5v0jkC
CKFmmZXOXpGW5f0DHf+mepGwzjmBTgEIhYWZBMGlci0+uIB49TMh2IU5VhBi0kRGLrDBCF9Tfn8a
QZCYlWtwVKcgoeyJ/g/6+c0btvsLJ/+8cgyO9c2Ypqk0nmsf0kpmsHLccE4sf1U5fHIXVbIsmr/K
huEgcS2dP+oyEjVceKNZGLqSFc7xDk4BMRcSLF0XonojMEBji0q6uhOxt3WBKl4QvHRfZYFYwhqn
n9LftYzDDALbboKn/197cO45ZkcY+6NiXdHLRatrpsnOoah0YiB0sXQ2fngXk8W4hUNy8lJRG0U6
FEY1qVOopgKg1GaIAklhVab3a4DxAQAcsRwDcTalq155f8gaNLCUwgM87sfeICpQnC24otRhsv+g
TZCTM9LWEwBhuHC+ONbJYXj7fbxA4iyb7Q4hlW5/KxzOPGCdL7LYL0ZIt1miPlG1sCEGtiFTpvC3
6S3aOqHy3elOlhgljp9b5U6N2VZQ6e7Dk6jticLmHlYTs0uVeJrtitdp1sYzP0L/5BcBrimEY5Kr
U4hh4Odmj1aJ8KaDuwRzft8+mpMsSVa0V8yyS/uRHKsa9AqEQQ9+PlIIZVliFyoF/jtVcYS9VxNb
/kJt5PQiP9yVQqe/dg0xgAAD3AOq/7BPa0wg6VMffsM/oxsNNjKWki/3DvzKqimcNG1rHqdLMPiq
yMzUhnLWdBPqp4kije8kPMbD/SUuK2KQSB8fsd8QtJo5nXnu4emrICiMIlqQlgWq1AbD0rxbI8HO
wFgeDpDnYwVqnIwLHOu1ePPWayggChe0uxtcj0MoFoR8spfHt9r9tJP7URGadX0gZh9NrwJVEtJv
hD+hC6oFzn4jrGjQkCfap//ZEvW6lD5nOyvSbhweYV3cMjJO+jDzj2hF9BCmaxOKsGzTNSXiGTrt
wyjkq4EHw1XnKYYPLUQ8HJSKoug4bnEI+J1h3smjRhm19MasGZNIrBE568+1Ci8ppYzzXv5i33bP
nSsz26o20cFI2mmWDY/5oeKNdmdxpwPEc+Werd2P8ckOkEh2BvslioV0I370Y3zaHtYgsnGixVLr
m4kLNK0KsMdIf0uqIBaLfKqDgRHHd3kDZ3PXMV9WRH/61Gug9wwB/VHkOTfRr/jnbhDJ/Fxv2Jbh
SZW6ieFekUeIMXTr4zIq8lvN5KZ+6J1acIQK27J4WKxWT3m1d6wizRNTm2JBDFtKdS8ZDDpV7bFB
8HEl+MHyv53Vbo/MZ8GWRVo/ykAkpOSn29k8MAJouW03ZK/ISz5TwWdqojT+8AeWN7WPgHHZ2fr5
rrtzJEzgRrbO5daiNlNkmKbt0kklTxKJM1BOmlfWijFDbcFlhsuqmpD3kGpz/3vNUB4UU56er8a6
j8yLf7fwE+12OFDAP7tOg8+6dPzlAZWBoNC/kTqvHPsRkc+j/2F6nHw+MdYE2RKL5VJXpDBGv9Cg
3RttOaukYvQ0hQ0hkCuI3gSbwwMlLaZXJnCDOUyraHhnNrX/AXrO2lKNY7jGB6s7OF86lLNoiBZW
CtNPWOyXCcne7w4I03DzpvpqtAnVyEV1vJ+/2q78om7zuh9Zfi8UZThROkr9fR+UQwulish/koZl
ww+3z4nXQrSduajkbQ50hJQBl9uCY7BG3I1g7ffVErU//wQsR1IiVHur+iJAMVhd/PVAmGRUMGGk
MixtVVM7G1qLtSECvmQ8Wvf7MQMn5+1FlkiTbve9sfgXPdqNW1z1Cq1VQoKTMnvPFuu9n5uTWfg8
stIrXI1HFoPBQCCmvbwXk8D+Lw5h6Qxyz9XklDwOv0j5d2lF4TH3ZQs8dQDGWyClbz2jfDIYPRRm
5E9wj7NoshSwuFJsPoMK4fQgo4bSmJbvpWxKV0b6hoIdMpVjFzsEIO1+MxJ9wCFPd9NegY3yGF6r
eJ+rnUBwJdHMe4OGrT0xSBjBTOuC2l8zFv2acunLgZf2k9aD0E+u0WJnlBPChZKrhHKYX98eb9yA
zH6Ldpk7wJpafw/V/1fVnTo/EkCTh1I5UgvuPx+VKKXg4zbC9zGQ4eZK+cFtc3F59ctYUBFj02l8
gGEkXXbr92RlTV5PAJZhKYoC7xkfKYLUlilwKcf8xVnymEP3u5pW/V98/KqHxG1Y9eUeT7WLAh6F
dtiOMGkZFqLXCDmnr8C/+wLy8YnO+Cpay12RO4lnP9FvmZj3Nteer6soWstIOoJu3QZEpJPjMpI1
Mg6wDUbDRnuFekrgwKiTHqZFxCnPIst0kEaZQGnJZ1czkbMN+KiwXdYc4J5QynqEw2aUK/jAo6Dx
OII/r50hAjVIiyW7dqBxD5jg1jnXR5AzO+3Peb5KyWg3Uy9LLsPRQUw8GIq/cFcxVcqrSTNr0ozl
70oOlTQkcda6xGjR7axS/lxy1bYFtIdaXfSXjdeyWMSVXi7S8J9VYYWhIvBPRthkOCoOKBoHAt6Q
aDDvoK1PynAOEoUwWKgukww0WEd2kfBNrJ/kDh1rxxBkVj+NsFl9NnFCZ/y0no6y1e4TYHC+nz0Z
/NgnNVFHnY9/vgW34BqVNfGhW6iS7GzK+JVW2SitADY4MLz2gajdpQw/cHoiBuODHn/hncBbgVv2
bw/J/o6RB6skUUMTYN1L3hzYWUCqdTZV3v0eIw1vFzARK+lOQwMuDfCZBgmFY8ub1KJAJYog7N5Q
K3fxu6StDkyszM02fXq1XcMXjUeIWeYj8sMFKBcNBPn7RP1GnoCrZLPjQYpz2WO8r7V5ld6vGmXg
HoqriMvDxshAxcAuYa7maXBdAaJ/x9idVtRtgz4FXuMtsj6CggAQCDOcgafHk1vGp/t0B1F8CB1O
oGxAPl+dR8otLDBBE0D7l4nS5Y13ZkZby73rmoT24H7b4DSo6bQljoZ4xsFxaZziSGhC5hitQArb
smq5Ls4XTC3rWwgiZ1hRXMeoEfUVlWKN2Je5YQTHJJFmSyxGYj540FjUHfSKck3TIMP0UE15GS86
LfXlxonmjGrB8h1HqzqPKVYBksjNe+fsaoaLTEdf9SPpkaJkQoeG0dWbu5N8tqy0GocVV2z1BpfY
P2sI6MDsqkUIWpX7qjkycoJcMyhiZt+Dn1Qn8J6jOXEcI9fmfhNihXjOTV0W5Pc2NPfTsdhTXA2G
hVi/bD9CFmuKdWs9Y31uV7D2jzHzR2FWV3E7V6O5mngfrj3qIEma0AyYLz7pKnWmOeRp4qDOJGNb
aKAkqHKb5iH+40BSPoC1u1SLvpayFtyIjEgjoqmNM8sRIwDmovQRLsYrKZIdnICEp1OGBfQOnmRt
J+supp29yOjeUHOpo2tXD4dsLyXerKwi4+ZAQxhzV0lQdyGr9gn81AP2y9O4k8TYcT97UqpikpFk
05UxWLi+kkgk+LCvV+zKw902EjNNoAsOiK0r65/+cC13YNzDGqsxRSr+WJLXzroUaykvarScncEH
wuyxdot7y5EyBVOFgCqBt7Al3bfR4LuyFbpfpd1xJK6Dq/+WSoRWJIcFEBypXBUF2lyzu2RrZuAV
QK3c4KBrGOMVXkfb9NN1IW3havJConczZAuq2325x6NzVe+dkfsVY+xeyVXW4jDhNrx6nF9Rd1fY
uc3n7qeG+FCigEkenw==
`protect end_protected

