`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R/8klGaE4rNh9MmCYuX/Iy4tnSar9y/DvgV0TXyRlBt9IRZHelFA67K+DNrfMVt0hQWYPzDPDK/8
hhTYXcgdog==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZvVrjbQ7D8uRXx/5e1R0+OcxXV88iVdf0pqBD9Knitx91Tg//TSUXrypu3RlMAA5cHZRKupVzRG2
gLrg+FPEH/sgL2GFocpUgOVPO8fyhrOEbwc7uoI155NkBeTp5PWJozWpLh+Yr1Sgp2aJhVtSgpYj
YFDXa/dt9kjTALZaIf4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HMvoHCd6MwP8Zy2lgNIVJjb4pXIOo2sqTbNp4dDZKqJPCqlFYKs3n08l6Q+4mkHxf5U2LfKI+mRB
4Z07LcZ3n9SV8/0qRhR44llTnmXJEvdwDcaQAOKGaF2xLL3rG2Y4TG674zgBbyeA83xopNDaLNrC
w38QNySdL/pxlzAVYgaw1NJSAxE+mQDzcQX8IG3bM91yWjc3OkViU98nzlYDiPwWcDOhpYq5y30P
dywTnWePsX1WYsppCwDfIAAiJJfbJu/j4S20rWiudH5evf4IDn5iWnEQHB8pbLPwHZYkk8a8tz5F
WsGgL6AJXdxxuP6fUJorkAAOzB8zCi7Jv6njbA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D/iXIWDsgbYOLrw9tTn7AqkXSZS1S6X7c0WPnuuSvZZZszI4k2zv/uqXadj0ziTR0fRUMcBrTgW3
/0cqsCjfy2broeHqze9cef2iPy/xfTuuFeL4/1hyCegKvwG/ilIGXcFXcONfCIpNJTiiLemAHx+U
/zx7fhP1N584mSnXGsY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u/IvMvG2nCOkwNyaSTeTlfkSkdhWkrKtOOsnX/cnnmCpNqVaq+x5AgWSYo98Cl05zmiglhAsHKsh
FGaPM38pSULjSSkj8teY2eZJ6lIi7Ouc6Z6Nz8ERJHTGsXnW11HQOK1467Z1tlji7EM4INEJqMkv
x4BJc1l3L0KHl4DXDdOiMpPrUQGeEnetvsz7ahn1JZorG1yaVayzjyMUl21P8/wvrQLVUq2M/+Lm
x4+c7ChAlzlPBvXBei1gmwIj7L0Brc8O/MHp2LdIOvnhfbSAdr+j1PsWawlTi6124oEA/4rbmUqM
laQ6qzxFVDBWAdjND0PX4GfgU3VfLuMptGifDg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vkm2u6bKaw5cE1gJILxPQNDT/0Ayar9EVnKG4+nwarO2pVND1GaI7yYgOpErI2H7L2PxiF+T/lzA
m1ckuj7lnTN9/B0TJMG0hhSc609tITg+nRIhl1vC9o1Zp1/ikQcx/TqmHfAkdiGjmUAuvPi7H71q
1IYLAzE8L6PvTKIFvUwxzlD3whVgpk8QMqiFY5X5HNpQAkwX1Heip2jpHwctRixCED9YpguUg1UH
giBUYyTQ6BTCGM7DVPXx/2mRtHF9ZJ7+T27SDomiQRDeLNxaLGn+ij+vwDwzzNd8d5TBWMc52qvp
6c5HTxW6mh8KQEiDUxBXBarfDoLcLMAaP8IjGQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 168544)
`protect data_block
ng+hTw5QCzw6rCTGKSyFSKJvZN3PMMwbMlOoCHMWs+aTEF8WPQj2KmSkp1pstiMAhlxG0EUnGJ4j
vujD/hEQUPKC9yH5D94sf4iO/IrUzd6RhHeRdNCEdlzLiHyoqYkBOnEB5zyd/WLkUQRArhl6HisJ
+GZyNnuCquigmgn4QTCDCxh+e36xXmBlCo21D3AM04BxKpPdDHfPQMI4c74CHl+b31Bdk1qA6znl
/9fEG7AHznCGbOctntZFNvHOduGgV6/xFJ4KIwMyMPo7vRie07+sb5pq57+Z39jwVg+Jp6ykfQ1d
ZOQv/IHI/AzHRMYTASia+C7oX9M48CiFRDzEgr6DINWgZDlzCUcTdkb3ZDrZJkIKozEDvi0Oqx3Q
IL1hx2h73I7QodTqlOPO+Y9015LZiYLKTuoEciwNo935QZJXeh29uZ9Olv6PLcDGVF+Y1EedpWoV
2e5HO25nu/Z3QOlhGFx9n3Wkkl8yoOc0oz+I54tMH6Yl1/+91sKXn7WSHSUrGCH9BH7ldx1qil2y
MjErgpw3Nu/0MMtfYoySB3RheEB3rW0MhNhrVLyMZbejrZJYKlNx1CLUG6vKWCtjQZOB5p+LXtAR
ZQeI0rVAjjO4luujnEnT8QBB09XM5ggu4+vU9lLjS68n59bz360fVT57nMzG3zkMoGCwyNwcqhkD
8iyPUnjJm2bBqCFkNSQLnjmV1iVPDzqtMe1qp1xfVFP95rInSI74T7KMVRdKoqOZgg9CEFyt+T5H
lqkGEvLeuJmgLorNSl7g0JbRvOPPAs/vOZtU4B5cuKoTd8mBKItKxM+BGL+ofIZz0sCXV/iGDF03
g8xPLG5m/tOyYVOfR8m7kN1Ofy6PVSL67x1ZDF1sfdxkZWvnzOakJtoUUIR8nNojf+wGQtYXidaH
yQMAMFUHrGSZWBRYPFxkGp/6JnuJgn/oVsFwiyqsDXLecWFCL8IFGawchRiP9lbYOYYdO1ykMxUJ
j5frI5i9naBC/iVy4U5GXIt/YkwDE/iMmBwS+whokrAA3oAdLRQx46UoMRhObwOVvKl8XVyApmVc
8BJnDjRGsxnEDIiNz2gTkurxqCJz7crvtwXZ4K+fZiuocmsEO03shbLv5FYC6vF1i7Y3MgDdrem4
AG8XDiqTnUJsXROU3MpxYgAeFaEdlqk8TbnYGNh0z+B758sr2WEVzLFovTsanGfhsi6RfhotLPev
ckC7xzPZWns8TGi1/Z2NSuQDO++95+xP8GuGqMFNejQXQGg7W/sDTuPMiMpbrj2POPac1W78/49T
IpDcBbLF2JQGjsIutLnT3u+qvfAXyt7dOV7dWKG71fniGxksrsyY+WBNwYE6EUsA/u0LH7ZtOV09
LTtY3i6CBiASSFE2XMbnyQ8kmqDe0C5wmmfHUXUkS1jRYsjz/whiL3DiQgCd1CP7hDVc4fiZRhb5
TLjQa0V5iAydqqjcEPQUh5UrQBIOTHdnOCi1gpu0E2azsvXbUKylIMdC4pxB2/vUNzc6xtp1K1p2
M94BOuuUZpEbeCYFW41yQmJeIyyYSKpeGMp6J7OaCnMcmlt3uIaid937p4besW67Bn5mCDaCT21t
I0k/8b0K2jqggRrRM4RToxZN2ignwF/d/yQJak5NSUUX9hRjeIBJSxdWARGugbq/iu5a1qj53aGP
xtLpLbT73iVPA94x2vsf6tNpciCPHBKFJ20texnSLrSCmoqK/XYzH7awrnCB5yzLlFpQLZo4WzB2
OAhmf35pfYg5qI/4iuGPUU4h80ljqyhPaClyfN4k/Quy8nZzIdbNPx/G8l0PQJfO+3R+N18eGkj7
0ekNp2fify47VCIwwB5PKXv/7A1yu6frrCmYwtDPoWTPFqS4y5um06ig9qPWQ201W/Nu0AxkoWU2
BN1d5jwj2/sCYYlPA2Qh2Lu+y1eXs9D+JEYnkRU+jepdRxYkKgGAEn6FlCCrVtY3OCww3rbsfLgF
oWL6U4VYyopDmA0BRsNWep887hdoqWefju4fhPyICMUfi77lvbEwm4aKKXE44AcNbHXfm7ujRIhw
dYyD61Dt0llOu4/LbnoYm5bx51JRSNtx5scYOs9rbV4ak/QhnLsGuPlBWLmyTZhZm5AH+d93FTBD
HCin20McUKyVcPkAkF6zhNXWjf5YLlLdZFYuircN5pOealDdRcS5f/OpX7R7CgEIxkgKhfdaGZI9
TAfeNEpAFQaUHoevvz27WbmEvWV3Zgcf+GQebHaUZEc8nI/CrHODMIKlwnYo1AimvbalUtr3R6Mp
lZRgfOcWzNTr5T9b0KSg8U7MJu2Q6etXQZtjtKhnbPZyHK6RqCPAnurXSEWWhVjRv6uoRENJNcXv
ayRtoVNMo4CYxexARmTcsDXe5sFTYnZ8H9xnm4pzcf8JPD0k0nW8JDgtH4G9db6JyYCmkaZTrWjO
zzmlrKsXUVHugp2Uah0QaWTs+5S2xYedM25eTiBaZ15mZCu/4LFO6m7EUPaRcSHX7NN7CsbVLYZY
R9ZQBSSO7F+M5nlY+KDv6cak10s4OnGvEjHbjKlw63x5BzqcqIOZZwblHRbUP9PknY7ZovXnA3Mb
sPAes4BBawr+0QAykAZSIhnqmgdloMhbr/amLez+CVgIxxVO8e7KELD5TB8hcJDQoUHmF4AIxA3J
SkihZDwSe/0QAe2jzOXq6KO+oITxKAZgYuNHIomMk++xp06lLoPQOyRl0C5gQtBuYqT/ZJNq/6KY
HVrW2g2wVQd9LAOlshIKov/6Hco0k6/m8unpF99HUEEnm6/z0M1mWu+uJFvJYQroEthAVRrjhNV5
Y04AOnBgCYl1Kg95R58iIiQCppzKxsPVXM8kEdx+U98NnCfHHVISPQWloW4vxFGcKVbBFCAuY50V
KjI+DXYtVeAXoHUqz9yn5t/Lyuu8+Mz5dzedYXQLt8JqoY+wP3tu9QjcfPqijKClmdWYI6hG/KVc
H6qAVmAlx6GPEMqpzdGbc2xfrYBYQu6O8d3F3xL6eGoJH3PrVEpOXkdutvG2BPRZA0/Wdt//5rSA
5orwTHjUfgax/b5AXLtl6YAhQOgqE9DBSxttHQIqwleg1UvYtgGTLEgVPwbENH8ZWWDFP6aC0Nvb
LDhPar+o/3Br02WcVnl7ACYhzIPSpYaJEHv3ioNx22XmIyiHXHDSRJLW/c6waHxnQQdRH0d+aSur
O4i59BPh9WdQ/iAE0q84eA1uOTy9AHqu81XNDdjhqNQZadOJRIcdyA7hkfEMdthMlChw4dG1WfNQ
hJPhfSiP0EeZIHVIyzr6k8XesnGHHFnlusuygo5jaCCK7GzMq8hr7f40SZJdyScyr4mq2tAW4rwT
TWU/MNHrHxlc55pQ0/I+Ws5ODJn3zXsMM/jvNms9cdQpmafCPh6gVxNuj0qkpahgfDlV4Z1YnhRx
ouEbpYLIiiORyM7d9we5kLW35/j1WRu/RGOntR2U/U9LozlIDh2utegdVBWWj6sL7qxKZTFADvQK
xWZ8uqeb6zDGO3yladyUooqMNHzSL5pS6ZIPo8IcASJfEKdriQR9z9MNLwkmjKHKdoSWmFMXtvWD
ydrwkJaVjXcE9zknlE4nef+bC5uOgzZQNA4+ZZwT/qxkeI/tlOMpbUMiIghfD+FemXBnJy23EiMO
zSicFzdvri9V7twEjSSlJvtFaxMqxxOHolS9RbwYo0wyPCfUcWf+7YZaHr6A+L0rxDfQvdZi5Mv3
VdYmIV4uqrLKeAcgTO6gsKkij8uQBuycf9u15zJm/lKLtNNXW0TYlXNBqffi0nKcR42zTADE9c5K
QTmyEw8z6mFR/KfMQw7BLbMI6Oy2fyQ8p45D4xUCwCFpES4g+8X6mR3EoOrhBvndJ8aissxFpUVA
CdtFmJRah76ogy1E7MZxh98BkJzsBcuwvgKjvvgShyYRfc3WsJDk3LNt70UlbDjyhVQonlvXd6PW
Pkeu7GyULfNl9W3Ibeo6KuVBowEPFdhw+DvpGxq94WbAMcjigClmhWNhZTIXPsquPTlONn7UCh1l
eYFlOvvUg1pEYVSWdy1S5letHMFNU6PgAMSv9JqH0JlIU7VnHjKjNyzRM8WTkpLY3/muoDZl4W/q
VJ3oi1fbM/R7tdNGSwsd/qxpZ9dnG3f3c0BDd4QDKS59UPLzESPwak2se/T+w206HFTRP8i78nNG
+PHeQexkUnVkc929Q0tmcu0CTHAvkXO+dce7iDRyCpnH3ES2FWRX3uMiP18UJRUCUY0W4WQTw/n/
xp3GyYbk0O9x8zsA4FZ0GVKZ/o40NomDvlSq/gzH/3q9HPBqgCPmG0ub/x8BONquDLnlN3ew+qJN
PfmiXigVLZfmb6mDF6+GttqgiiaaWuOCEEvOIHovQ+QIBcG2mocqVZ7eI4Qm8a9WRKbBma3kPFUi
LI4w284C/V92Qfb0IN8HklQoYdZaKIqufGT4iWA34TebaVZctls1TYbZblNVKqVS2X+wchxJL2tv
pqH9/H83FEl/GIQ4jZT1uDxXHcnizCoJyoESjmhuRTJFh94pHYJ1MYRd1v6NVvXb3UDgHxQWHdmp
gao0eaeAtTSaQzb6u+d1eQH0kQcoLuDF5IVfm55F52Guh5478GKUKNsHhOW98s8FpOheSa3Txouc
y4sYrZZot6SSRLKw8dBP01r2sSCiCa33NduOOP5ax2TbLYal4D5vfQjis568fhmrqbZmV5rgrw+g
AOr/FKpF43zYcy+7aFS4tRwlfad5qDXErrph0EwvLaKTgmv6UNV+v4wLzEY4YGPt/XStr7t/qr49
xGHnOyrsrvIrpT3yDi2srmFqzKTipZwAKpVUbbfAh2FLcZUZ9Q+W7tZrvPGhwtgoPWsCc3C8VXt9
pAFDVb6uvtPogpSj+x+/Eq6Ozyd5BWiUhsqYSLo5KO3T4uhdVdVg9hVSOtmDBDEfj7PxChIp+Xcm
k8oO+qhG6nGCuyU7d3XPeSUjENDsnAny3+/6EfzoiRvTU5H1FfALw3uNYcegbqS1TryjtXa9UPmE
5qBuSi8vWDMIEByk6xIsKEcXTA4Xm+g4xHIFvZsZlU9jjbGDK3g20cVgrdmUmfpMZggvdJAJ0ywD
eHYQGSWrvgiXTcA1QkWJdV7F3Jr//WjzBpD2q4ypfI5IUxoKsABFYNrmndknuVWwafQ6toiDODT6
grEihQI09t7Me9+d1ibkYYwd0ytfTT2YRF/E7lrKSLMzhYgYByNMUIFod9wmHGLN4I/vI5KFeiD9
UoAJa0BsO7SrY2a5prsuxdM49QJO3K7OgQEIs2UmUcWoIJmcwQb0u5GPq1h/Bqi5X3nC4icJLH6j
oBMlEewgrGc4QbyXE9v2MwS/JeBf2EiKKMJAcXfGESOC+cS/7mPQMdJKiykBbtTgnLQksooqMuiH
WlgJOVsN0kNY6NFIkG67skiYiUPfAbc4QaLuLof9ZHpZiGy8rRn2qsJoJPEM+9GyNjVffgny0UFa
TmEhgvoxOQE5qrR68EhY83u/yrMHwPPrLQN6ugUeJ+UW7BJTFSWZceA8s7P+9NAyBUMfmu2Jlr7u
AMQDBP2oSfMGPbj31MN/gLXKFzTIqAcomkyrHg83Z08YWE+KPC4VQKI+aymCLUZnFdYMHVAk3fYx
GTVJjFvBaUmyc7tae5DlY8CHPuhnrjwN3HLT+IzpGnbatoMmrGYj6V7RkBJ8mB5zCz7l321nf4Ne
iFjuUbML3KwwsIR12iWGMdsJ4YKOMZccA99OnyvEq1ut+S3yzEfM6Lz2gnICe1Q6UIok42pSoA0s
8igW2a4Tz4nEIkiNJNZG2fT58nYCkxjrJWA/iIz8PIqS/OFQfancs4rE2dodgGmFGpaX1Se8cTbQ
GMNvRgpOTOlFBe8hFQFurJ3WByR/bWHxmon5NMibhX8TczAGJRGx9yQOVnAE6LksJP2Em0RNoShd
OOuoyVtj40bwZn8szcfgGopN9ad5AIdnW1lKL+LUDJcvL4za/smyAyd1CpXbUGQYK+SHx7RcQVxY
/faXkAMfzC9hdywy574eBD2uFUFZjvReYu5/fSxVxG2XTlSwwWu6PKPmIQOpPRo+081wt9WJS8EH
bD60jauDxPJKBTjN7rDNKEDPD+7MbsWmzQ8NbrFScdWzhmZRuiolFyT2qyIlqsAR6jb7JDDbu63w
+RrJnR3vglLz9+Yipa8wXzwSlnNpVwrZjDkw8/Vnh9ZGr1UfLbv4X574cPSLg3xiWvdG2fGz9un3
lXojf40pu6adSJwAbyfJTPT5TL/q17sm0U/u5hdeRfg6Q4Ehyq7dWu8g59EcYYeIfeZ8stAzQMFm
epNZjMPoOO3GYaUzzHkLfOdYpJF6/UTpYwRpsW81zbg+M9hxZ1h6BQoczm5fSKbwP8eSj2rN/5j0
LsuhawCfim8U1bX1Yv5BgbuDz7H+xspfH/sqeNuOeAYTSq2ph94wUJ98pFkcITuIk04KUiobM/zT
9tyX/7e8JPmEAOa8faOCgvLLbCsG/Kj9oWugQexX/dzXAHe2n6PMWMx5wG9JRdqFOMpjEdq3+9vy
dVxZ1C4NtFR9sM7fivhmXSzZKvO4jl/XZkrHzbwgeYmLXN3W28pUuqjjU2uT3GOJgOotcZ7Qhyz1
u1xdz8n3kOg3rY1VSgmOPjIbjvsJgKZbldpPf/Scj7K5mWorCTu2zV6BoDhpNbQbS7Sv7V5oJodu
jzMcDJYKtmpf1Dj8dOX/7q+tsfUN5umggqnnKsA0q176XRgiUdlGpA2UhhLlmNyqt8z4xllupzNJ
zFYWYPUukAV0WRbyqO+aW3qA2SC5J774Zlsg03EOzgKHSL5exQuQh4PizlSkBP67fkJpTmdSmBbX
X42xxwOXTvE468XYFlve/f204Yde+FNzWZQWRpmvNWAGNhAP0Fe5Rrm32rll+2mDhfHjDYEX5rQ0
n++MizZHpdHxtASirRRpvJ30RUdaaleSzUBFsNNbqKP2KfJDOT3drmeFlHdpuzvIzvcY88A8AgtH
y00ii2sxRJM70L/B9z8wuos8GKCepMKyRto/9Tn98+ZbPpv2DB9v7D5V6dXz9BwUlU/zj1xxHQ+y
R/5EBAePOtrz0ulWh2zg4hr7HksTLJmIZkqBpl9FK9ldaeuY9A6Y4YcW69cWVbhx8JyNmb+9c1Lt
yV/isLo6w1bri1gopqQmO5t/hizCV8Oijw33xPa06SJuK34qiV44tVcirYW4e+I+qlBrcm8zt8GK
YiySntgtczLQZSNXwTSHar5eVhgReVXmVrMCPkK1Oz5EyvJypwsPgg9eZWh23svbCJj8vzwyT0g9
7ME55AUjTLKYZuGvxX9sYFEUNzo9/rtl0gqy0i0TJRCgH2LgS7HXZ255Y2AJs9S0tPPV9Aj4Igbo
J9kg15Ocr2M9tedFooriXcO7vcKO3HKVmBfiFO9nKike3GBPHR317XNyPDLbc5HaEIGIjCIfuhid
EBT/xzTG9s20qZe+b+3Lk2wAeYpK31Wd8qvXqBcvwjN7hN67BC/0B+1jd6WCx09Wnm4DFzMrMvaZ
ZStmJloqVQIsesd2nEV5kde6++XOhOUE42me7HRinfzQUhdMfuT560UFA1+pFYxw7zqFoNL2+aVt
be9y486SFcgAIwRVkFfVeObfFFdyYGQuoxNKHeGISsOtmWQTjmCM7grdDQYv19r9MpGdTuCaDplk
OF3gDzHd2NYKX3j8B1kzrmdiSz9KRUN0u1IFhZtw7fbQW2mcqOq/VpdQfioItKM3eiS12H1X07wy
+cUBU196zFSOHvDx5nUIsQ2HvEB5EfAxh7jzVVT4phoUQhDTcAHVw/pVCqdRL0+SNdZOKHnNsjnq
yyHCKbkcYSG+DdSxqoh/f0jNYnyWJgHYuQ/fhuS15F9ycphcOf/VjZu/QuDJPWNsqNw6iNU9h/if
2JtFs5wPIUD8SNnFYp69hyL4Qhmn0eWW/U7ytws8Swwp5taCr9jqwEkLOigsUSH8wpaQeB5/JILv
K9ICZ7+Sknr9T8NMRgQ5ULjNpj2gI3B7yJ2CK7jMjbIEjQXA6DrgWYsrJ2PubYAtJqMf4OwCn9A5
wQnHPcHMWl5w4uww+Ei4Sa7DMKZiL8vcDuoevR2NRvA+aNh+kbHTEec4pvzIqrYJA1d2JsgHzsXZ
VjKmdbGgvN2NthPRZoCyap4TuWmuTh1IDjKVDOCxOR2I6wl8bwtY2BcAEhg4OQunZeCOc8k4/7sa
v7zhHq9jbpomY1qeXlVGWOF/1XjmsAY9NV+H4dDlbP2913V259Evefa1oT3+I+EfaMnV7jlWfVpC
Mefk+GknI1QT64WU75L6RPpRxGp8bQHbX8DKVhTOeVghVwwY75hHwMbjlmVt2lQUGRTDn1EWTzNN
UvD1rU2zHOD0OpddRm8nj2sgy2SltCQxR6hmN/JiSUX8tK91AiK9snX3+fv4uQfou8uzbLwPwjtB
K7zJ04GRGfp86Cn2yG9f+HQXCZPepchsPwuJvG2HRoDfS9Ac4aZ3QaXGFpMxyiTQMFpkNBK+9nLx
YjbH/z8PK8NWkAzewwRDqqfnmuMr8M8NqfztKx47WvHMwV7BAY8df0pfv7NCzFsbrYlpKVEN8UB/
ydQJs2a6ZFGSjwImA/U9b3lgci5UUw87DQUCUO1GS3ce3Aa5eLDdA1F/6fMJm9PsKGCB7ZCcQ+Kf
5LvJ5Uzey4wloFY4gc8o/Q5y/IP+IrPq9cZ2QPw+k3Wo+YV/N6ZnvoRVDwYjnc/gpRc0cBa4IJip
+qivfLcprDLaviWAcL9VTHFC9W2BbgReZwt+UGskLFcYkm34BgqgV/aqqmTA9n0vEKeMc6oy9qx/
Apbba/QzeuwKFsO0K0tNW4pB9zDc3EDFw6rjIiGnNFnR7At88sfQMyA7S5mwvbi71Fzp6FOjg51t
in2HiYRpl7EudURtjg8bQbQ5gcJaGk6HAEm85AuKFXwvzWNfyckT+EcU6ZJBvxyRSCb1wadL/VUi
wCkUuPsNduuWac2o4WAnsWppyKnDrYvZSwdpVoEjoaPgPwl+JzlaUVg/RUDNc/gWjjcLaBpFHyID
3Rpi0xC1m5rPA4sUv/a41NNxa9anIAbDIFrUdu/hYGHho3+/4YksYQ/DKcqlR419HOmxKnYjmvob
wEshSgdhSxLvf3XWOGrp6SuAISZeRoYKFzQJStzV+nZ/53PmOBZhzscTA3uRousiWIM8NcrEyl3w
Et/UfHcp/z6SHj2M2BFm2dFbHCKBBPy6LRdO5tn8iKjio8i64v6eDs7EW7dOjfR4x2Khg+SNFcLk
QQ++Mq3w17CD2M7cVwYGE+V7fjwExQ/UhI+JoJbHAPVdWZCaX36Y0S5y5BDbBHam9l3b4ilkttik
inc/Yuqe9gAMf4HU2gYr54yPpAtJtIFxMahD5/Ql88HCXlSC1eKYmK64kV/LpZlKhwt8XOkHA3at
aUmU+bOBVDXNdF4X63wunRNKquaZwIVq/d6aU++S8OBAwYe0iR+m6YRPN8Yy6PHiXi5bAJY064/6
qJyX89RoV4fcOCxWDhSSm750zR6sKlxe0ouHkmtLx8LrO3iuW/iQj49fJuJuS1DftHE3vlxLw8FT
/JRzmrbCn7BCYF2SS6GQUx2dsNt+RtRhTDwIJ2Zi4bKk/iOZFipK5bov5NSO6B2AXNvSeymruH8c
A54WqcD4ZAFaR3KEdmpHZD0JH9NXzBBQTNlr1qY+o90tANueJ1yk2w2f/f1inDdrrf0wyAxM+5fE
HLgfqtN4sUdpku958SIlODBsTMWSiRlFDK+WZ1a9TmV0qRRPm0b6ASOCS8EgFT7Mg0Ne0mnADGXD
KberOMlzRdYpJTXPDhr6xpAEaJhGieujN1zMrXw+C18FrvDzcH5K6H1SyRHmnQ5pnsQzLAG57MMO
VzJkUI1seGahytpm9IHBlrW1IvEjujaFlFlmHmiShlo/0awXYqt9G7WmPwQS5L2nXKW7446Cqes4
SHYi8bQt7dZVn6CdgBcc6CdAOa91wC4SxIIsC/KL9CZcFj5ZlWmPKGIRHnQ9OvUErNfC8wumH2pf
zlb6gUAUm3T1vo99u3g1Ubp0QEVqPaUo1tqlAU+5ZERaD1nM0LPr60Tk5tUXv9oHOUpKgZ6gfvb4
SDaFZ79Jwhow+JH60budLeNtgz10Kj8FpksWqioQebUoiq8Z8SBXhO1bbML7T9ekezG58S5gbK3m
C6MrQwT037GnYa6AtAJryDnXwA16hf1e/TG0n6Eo/v6aU6u+aob2s04U4rT6LKcoMFqJTmUE3gDq
96nWX4WwaV220Iq5VkIdy8vfqZuSxFXZuPM/XIG4Lawqa65Jds//kC7QYcRUNAc9y1/b8iS+Fn1f
RqH8RADcotqfBpllIDiX1vSeEmTZ6R3RwebUXShS3kbLThH69ojbhXsy2RYGuVJ0wk/kS6Q7yVex
1EogyQlzv+lvAzGrdaF3jzQaKBkJKjBk5KCyvl5MoYaAoag2Ryn7Ege+qtZWgs5ftivUxiACd6sN
Fa1rrY5kAFZWxS+ejCGj5csBq7mMm1KtNe/yA1XUSUaOStWAI8FnI+f/6tjqm2gRJ0lX/FrneVU8
c44mpkhy5/zHbQIKFpUk+7yPsyJXIxHsVAzFFVCvsuZoSPt7qcvWFF6VHCwjbh8hYKg+T1MW1NJA
QlTReoonEecyN7cwzpzb13pg1rPBa4XX9Z38WI0VilwyD5JHn5xoKaHsuvWPBGtdjNyRFWScuneg
oXvQ8XdMiNIl0Ci7ijSKJhqJjSV4qE1WVvc1BQtNO4+IXUsh4g/Ea00TKDhwkCJsutGwtezFIbFE
CAmpDdxhGuklNUm2wNEYyEPZdyf6iBXJRkAC4FgXuE4elOqvvjLGuYdqUjeuXZZ1m05ivmJ7nRDW
T5iq3892jT0y9kE1DrAp12BAhf2Mi0JNcgKLaz0WMcn32wTlqmRyQ7Mv7PQzPJ8P5ddPvcjD/D2L
WNviUL8UGP81vfyR5McMwvFun1X6Oi+/MneAWmq6vOiq5emZt6ddSaTLaqZ12hiqvWDHynA5Mn82
EOvshNlkMt9EfxEwlKrublNpX3th1sptr23JPgnQ5FKYlUEw7UhX+q5lLsgrNaHbIvVLrCVWJ2r3
Gr70h4AEyEGpUvO2HtJ+FCwSjuXSlFV6dEHudhXGo5HnRPJ/cKsiIzSps3Jp6q/MtJ3qhks4DCua
Xv3Xc2ul8cXrIHmvfrQn63rdHp8SMX8gob+zj5j1bCkJL7lD+ShBg238V5WeQdkgFw/mkQ2/3U8E
oKYmipx5z+E9isZET+4US6b4iFwe3UA3i+R6dlV89UYYY899zf8Qx7mbK5qHqhiLQteSQJmSdBlQ
/RZX0TYrYrVpIv/yUSWJCPETclF3bkswFH9ZbRd+5fdE4zwR7l25SV0fDg/ZDTFN0Gh4YcCcGis3
+dR0E9mIpDHqYSilogJb6WwfGm1wPZ05QUH5QKC10t35VKsTLFM31Zh017oYswdM9MBmEc6U3E3V
wTlHtx7uBznvqaAD/6BPajzplqiwXu97JBQHPZJcrCEMfq+FiWGqBgcisu1NmdW8EZ3LlGjAWBv7
40l0zIMtYRtm8iplVg7cIUBrpLEPF+OgqU1q2RAzJFRcyocmhI0gyekWHD5N1MuSNJQwKhEnS/a3
4cM+OzirJHhkuUf+6BCOwo1wr3D6sN9zXjYdw+a8bi1O5QgryMD3JNQt9MbYgT7Qp63G+qQWpjfV
78h0/xdVCuH2XBhYbQOa+3HoPLThSxQUCvw60fgDddg/JbhSk6jj7hmfZ4sWofn4LZzibrq/ifxx
GS1OZtRNuwWk1DBvVmc6/pWCRXsA6Y2tQix7Y4A28HEm03ZFCns6NwwrbV0Il4xFJZrK72CFKGcx
wHuiK4KHTnFhPDdojQEDc28NW1B6Z9YBxyuWB/076wTTDkXPFLoQ14jyuB9BJqKqx+7zt9+frd9S
2LTAlQjeYYd/iXVwsP8nRmL6xOPHdNY9xzoux2jEsINIFPkrBPvOOVR7JTETgyU6xvvvJFxDGB4N
Z4B5ruCHQAA7qT4wTKO/VezdiBY/IR7ODeQ9iTYWxfYMUATOmPjqtLgBKsQgvVxvAl6m3MnoMqF5
vvQpLPMyd2YaibELdiC4FRKugZnxLn6oz23WYl75cUdCYv1oc5JQj6cMwtd/ZC46MN8oobvT2cAF
kpVQtAE4/VWc0DYAcM/e4Bmo/QfVJJBtZTmFAkMyRhk4dJj+hzZr+gg69HjX6G7GRmz2zUrvDU2I
O/dqErSViyrXwMI1+0/8c6cDLA4fWV496CVnDu1+pAooNb1hMFBMQY9crVmTBwU2QDRtcswCU8Mn
+cXgEGT7KlUl3LwKK7nVS0RNgKZ3365G5h9qS0zO4eWonP0cydbVi6byXQ1dH9hn0HiInfwC+mWW
Z+rNQfoD/vSo8ZavQ7UMh5Lim0O5vkfDCHhMs7e0uubdUVy2rGodSYrjsmrGG8B9pqL3A9NWJYcx
7FW2rjjgUpjQY26xikf82DQZYGc9KnfmQO2j+EgrDc5/NXSSZNu+yzD7ILedJnscPfSsHgKGXEoB
ue0ifEJAs/Mek9839dtlevCDdYarSesapmKE+q39MFr4Za27+MXhzia7HgTp8OkFFW8MV+jNwvSh
miQ5R0wpARbkUd22CVEsQIyw2WyM4xUMYxvsheH7G/FhNzfDfnBKSFdzDF5EavL7kqZLC//2pJJw
jr14GIks6MoCqeRBLh4ylCq3V2mi+963D3R61BS38zfD5/SK1PydthiKaXd4XDvYyuxjKfmqixG0
Jd4Bh4qlRyDZnVRC/RwMwALdg6IxsmCV61EdbCQBkTFesoVCCbGLpyGWRwqsArw1n4ks/dlW+l7O
HjVwVtywXB1UMxxkdAinyHHLw3YK2CkUIcx0y7iBIQNxjxIJc2kHozTpclhTvTY7pDKdEfv/J4ER
TxZn/XfyCNrpthuXXYDK3mdJQhE9iJjvEZLGFp+9YmutE4jccs77zwL4NGpWC+904zACQJHPTtSx
CaSBLRQj54bHCJUxGhqAIAIFbPNmPaxSu9Ke9uh8kKQivtKV6LOW7taOgsSeQoxm6dADuqaBJr6k
0iGNFPH9b33zDDkfS3eTZHXD3dvYHb0rna/WB6sbqdfBXpdrpnROhj6hnWdqQDhWlvHA686HpYnI
WRFTZxHnvvVjBd0P+unPsG+m7rI8Zt8ejDf+grF0WPn84Rqr4JdeSEikNQ8YZ1V7gCrKJ9VoKO0Q
qKam9Ks5M//NNmwOhUu1XJtja1Mwd+0ToFpfFZuS/atkll2gEAvnjQd0bpaB0T54y5xbhxH8vsw2
v9qZblmmFxqi7N1BntTbw/ULbGsTT50mGKNsSTjAqm01M88FffQHOm1Yu2Yn4t5pq7+PTRJW08rf
dAAgevUrMW/dnzbLyZc52xYnRwDEHxKD4gierBf5YMMRlSGtU4Z0Cm3/wdgu+xIG7dPIYx57I6IR
nmmUYxetMHYn9ItAQUye2aBGghz4MpTKz07JpLtlVwixOxGdpTDkoWSj7vsBpAK0sn49MUusVtm1
3G5LhOfi5iqwZUNhiCBxYxwPJ8tuWLkygbcsdM8Zz46HplMwJEY1YHZmTJdnUvPj4K42ZnxLkxZZ
QTZ4WYdtPR/L2A8+aOhhHOSrDITzS9oKRPqfvSAAK/u6fts0OqWX96iTVcmQ/3I2NTwIK+SdOlEq
LpOCqQp2cFILv7G70+IvsW4eC5cCDXlogJpxbZ4E3z8rbW9DiwYWQV4nprb/45Ga+6R03obz/XFx
VF5xbnyV9wM/Pkgbkrqaf/4qzcY76ZAqD7l670d3+5yOUq/aMPTdmOMXBamLm4gy/pPTXQu5N8dX
mAPG7yEL9SIxzAM8YlT3BGm8fTk79cjzbVb7ohBMN03KM/aGKcWbfvGVxrJDhIB8uZYR4G0/K+N4
z8A8eoa8q6CZw6GMWJuw4l2CPkdNxyWr5BiHK6IC8Obxf+Iq+u53K921VfiEnaDh9Sg3QfmTshY5
KhCLpDCKvlcJuzDMCDwUBPz9stDMaZfNNakyfC9wC/i8rwWTOErwJbAuWXlVQyzVxWei9/vgolsi
erXvSg1rBg7wFgb7POz1zeCDvUH5Zm4g9k947j5H5l1528+Iwmw46dmoAj/vk3Mm0MUQkHoPZDZL
EiB/s97Xck/Wdn2LAIEN2monGBU4ctjOkAPJocS0+Xzk4jxkbLBDYGWd/2KJ59+IW3o4nYNDx1VE
ixmuI8NxhDRMZa1f7jYUGMEozGWgNRas1d3fkEK1KsCCvbQYoLGJRVM4+PK0sgrMRPVX9+Qo4LdL
z1L/jdVFL3MQlHdqlGPJNgf2r+oWTg2t0w+9F4NSph1i9+cdcqbMBcjiMrS1vsJnrGYtxple/PT8
KHJ7s8IrAKsXnYwxB++cRmmUi0RdYoKBu01pYeNKP8/OUAopxq7+mcjERG7rwAq1yHu2xHAy2pUu
h27nCzp6jxIuE1ECxRTchUztS/NweKGjcsmwlaU3FdY6jFeHce5BDXFtg8xEoklsIebHkjCHwnfk
jCGnS/6MGja9gXKoTBXLd8THIEVfbIrKgLXYR5t7UAbQQZ1CkKufFpqEud6KM3bW8h7gYZmZd2H2
Kq1mZ5J2hjyuXDVw/7TVY/+ZF8xELXzd5tpvEzXn1k9aocraISDYta7U5O6buDPmkYYGB3xksfLy
6f5hC2Ino/Zeh08dKnj1zVd9jz3SBNbB0yUJdVrX0GY5xNhmmYAVp8+dwfOl+v0Lx4JyyTvC00JS
1OoQPyhfJHakxYielLtUFR9/wlCfsxCsLBfez7qSAnGnyjoTo94fYaQStDKry9sysrY0+SOvKqbl
q7YwVnuolJc6gC0Zicbn46F0qR7g+9g/0FIRYcdAYNhwTeNrfYsPwvqVJu2SJZtc0MQont/seHXY
chALLl6hQNLetxcj7SYTedYYXoqVfI4o222NoEe8h54g3pyaMdVS1L+JI15bcfiLUnnBvkyzUf51
gcq9G9ir0spYtON1Jvcm2t5WgS8o0mdo+hvybPaDal+/y/TTSZJtkniRS66FTM1ElfIDzKjjch22
GBCa3LuY4lCNpNgRV1BpiZK+QRxS3SF6dRUEky7sFuRScFKLFpeSRWao3NRiLNA5XaPuHskWvysN
DUwxOnWE7qtHQ/GYrlTN41Jp2qPaZiWpdwQ1BKdfLJQPoh1Av0jlc+Yb/BFTY0pAg9nPhsi89C0W
HCC8yO2oPATthjR8oukaGC7IZ93bIsRjnZHejMwtTe6R474QnVvJFYYf8VkrhpYPEiomeGXA0VtH
3saErGYZp//uv8Zm6qzYrLoCB9aAHBwSCU/FRADLYIHl2kl0zrdwsdrgtJPyiuWdB4C3hsoJm6rl
DddFYrS5TgfB1YUd7DgkrcMtbDPf/BIDqsmaVjHLms8emMSIzYllnQDC5eSCdKZeNZLrYha70x3u
vnFG3pQNn8xRq6wV3KgVyYXWL7iW1KLdvxjUQrMDNxZ7NDYorijuSoNI++VDu/I4+9YwNSx5cYA0
Rq1Pr+S+f1OeuvlEfGHx5UTSqS4inF1B0R0KtRHZXGHuYoaOBtIpj92GzaazaYCqaT8Jyfs0Ke6m
nal9bgudQxGN8oD/JeZ28JGje7LP2AKjoKJomimgHvSkv/Grzw6gpx5nt3rQsFm1ctNW4z2QQbyz
ZBN3GdA59xnyd2y63o7nyFnc5rXp4DXQbVz9uxlUNIxO26KUmK3t4NW1/BGbHgltHwrf0+mNXWC8
q4eng2YOKSh9lpRFm/ZX+j3770UOGSLxxjn6O3sOwShbO65dyGktERmoHqM0sx+bBP3+gK1pMWhu
OcCmhKAnDQxU22v7clgiGMelj0oMCTIneC8PS0HJ3rKkzZ634lnE2jAtghKfVUidoA7539F7AEMB
gy5qNII3KK9aGsG1PUml5rPT2lzOTyApsi+GVMbn5u9SeYEhkUUwS1cmJsywirnpIK16IH1+uqHa
PGKDZchcoT3ZKhSjg8GdNWerfgia3cZqNaprk/uJo0UlEyffNk4+PPI3A1HNT1R8d+HRbYrEOoaW
rJOkCiVmKRp0Isc5Rzso+irmgqH6FoZBF2siWzLSed4/RZlqNPLpdA1d8Mesf4rW5zojux+rXwRv
VNlRK3GFt1Y9H6a7DX+TmioSDSiIaWN2RHk05MInjbXFfUcWZpLZjLsgNEDKoOq47bqgEu8yGftY
CACqEt9NVep2CPJSfTGtAGF/YY2ofTX2Ie4fXrp8zDQSDpsd/Mo2WleqinlXc8fDglZoYA3E76z1
hzcbu985lesCq3bAjs6gM5Y0YIrTj2ys5ne0hwZzQsZ9WygtZVTdu/HdRSoz9/iDUqCGFFcP4ZH5
ZNtMJ23ZKKNkX6KnQov4LnJvCreY1rqkUiWfhXMozaXodFOnvqIPV+M0evWAiDfGsRGyt0Lrrk3q
4ViXfl/lB9+BW2dNC+JMX2+UEwXz1QffEajxAgpAHG19PWHzjTYdRQEaRQ/UYxCHyfTN1nerVO8R
Y3nL8vbdaBFI0uZn/rl0j0BA6fhGcjodX//dClTS88CXnggmuXeqfgnbhHk08hpx2mGApx5AYYq6
JA7iPIKP/+OKuHtgB/DkddB1mDZvkEl7JPWkj/WG9bOJqc+4N3S9RTb0GG1rh4WJtbpeMy1vCeYS
glrPfg4QThCfcFDT9FuPkXsVUGdpmGfv78iiJ1S8w4S8yCt5bf4X5OzU3GJRTYtpU/GID4wn0H6O
60IvBJ0cDLd2md3k6sJfxgTq9BiS5vZ1zEj6n9moQHtLt99MzBWptU+QIGl8wDkDsRoyglKLTo3u
vUIm0KPAnvjvmF2w/+LALalW5xgHe6FAbm4ZLsy1wRE0OwUwJFUjo1wwwo/NDsEvR2FrkzqvJwCE
m9HJsNwfZpQXGpEixgHd50hV/dykoCAxz9ujbxTELwOM3nlfsibcU7/gW4AYkIY52eY1OmHuDN5y
PAdE+reJFnTIKQkP8DBqAcNJK62xqcc7GOPt9bLrAS9x5mrmiyj91gHP8eIicY56ntEFc68DACIj
wisjg+H3K41AvvLq/gt+ulnz//na7URUQ45OjPspBMnqRlenuq+I/yeXeVvmnbJDAF4YbKz9fgva
NL1aFnHEtxIzsFbJhwrVECyk1B4yb8bb8isIlHCuIIMrvVEkAK6F34Vo08OqiOgjxabEmnHI1oRp
krV9TMvtBruK/zELjceipQB2c4QL4bm3LJjAVkHhtVvbdZLMY4KPrRiqigWE88sbf50eZiVqTXVb
JBOROaG0UJV0qdv1RDLqoISo8P72vc0dhkg7jE7plBTBAxWmpRjRNKOQ4DF8rlm9jStOO4ljx1lx
M1Y2HkFnuD0NNY07kp71YvcS9nqfLTm6j4UHYNaNwouN1GqprVQypEs2VWEzCncXN/ahwmQzkf6N
60rI+1cMG7srJj5OxWJSpZT8t5HOVPu14XmDDNDfXCO5dS3FJTkr30uGOzMF+ou+Jq4jrwuLTFSW
XoEFA1HPkUAbhzZXcYxg1XM7w2RHt4qvb3T76b31mBPSTeH5OlFqS9tSRFS8SxLNgeF8egwE4/ZX
SMmVINWQzcvt3H7NQGHgQqLyvfQrEvmbZkwP09MPqLl5mXpA/CctI72CjgFvDlx6xl+g0gJS4PYD
eXCVboKtnNnNru9Iwg7ZrxJ3s8L2p7zvTlpcjQAkJqEn3bSiISuEBwl7m6Jgqw6hDvAa6KymGqp2
iW0Kou+fyu3pln+vBH6iXRitRGZ5M8kyIBpP+gBFdvG6ZJL0ImuprpPNRRIfbCCxxiWiA060FJ3u
7vjLZX866ec04EGDIhf80kRoMWMMoU76GHeBNNu/mUL1Xi0+atU2DjVYgOR53GH3pVrKDYsAyhA2
+FYZ1UOgbp/u23wxBfpaG+mq0014gLB1x3wVsfO/L5nbt9Rxp1iNZKl6N0ezOmzqpRlCL8T7b/+b
ySe6jQB035GFM5eoOX1pqkH1UvjLQ9q+459ug1LMtji1Byu3fvHZHaYmqMWHjOmrXBOe37jKRWVJ
HX8WE9xvzPx49UsPHGDt2fRzUTXnFumP/FBaJ0+KZkttCuWtBnRoZtmG6na3woLBqVS0zykAAydA
9h8HkAV4A5q/aKpS83ddyGyLx575p83Fm7IXn9pqwYgq1WUhy1FbDdZkpG/59Ty7u0q/7FQD8MBQ
GSQRpchP/GAJoeFDJidg7/sAIzPxlGfcAXbwzzD+Kb9Iu7A0liZ5hVt1RKHKqdrAh/cYGEjNEDxK
ZabXwr8/PnFrYdJdHo80fVa5Na/W0vtLtbPQDiGyHnwNFCAKwqf8QjNWIGCDh5PXNWMD90cAAAwG
7srh7NVH461kW8jC5eDoYW4tpddFWugwoMWoZyPf6GRIK6Rw/6SAbE3J44qMSiEFFVdlQWg/xZQo
tlLB4aIhOQ2xiOTGK3mhMqZGn1V8vKG1fvsukfmN3QhJtQlGCMr9Lqj0t87qNA4jUE4Vdz4m5+f+
LC2W+JruJEx+J00Q7Vett8PhEAuCo3TwTEYw5pmQZpdGvQMjCx75NCX0SKYWE/FbrUSVgWEegY1f
iCIwac3mR6LxTJySBaGwkrGAiEaeFJpyLP46GzBHzNd1O0ogHf0bDU3wXgn5IeiShFcrTdWascp7
rNxYjZ6zFD9J4xrTTs+sjQMUgnYjPs7CXVn+xEq9xJfvil8hsOrx866n46IiwOtsMQRl5PcAFFNM
Rl2WbnD0v7cyrEPKaHexQ+jd998VZEacqkmDbRU417d3rJrsFQufNjdi/AlcqNld+OCDm1Fq/t9e
xQWK2tN4k6IJS8qgJLvzVq9eAmQkmHZokwMk2LeRxX+hKhaPjiz9fl1yInbuYNRWUufGz1IjTk/y
Bccv7jwFkKnxoalSLkT2fB41SyJxfejx9hwbYd0eu4a+harbfduhbwZfaMu3SE7vkmFoD8qIOyKE
W1BY3goCq0pNWLLvAodxKUBFzrI4YfHPK7+ELOCC5SBC5Z+a7OBi7ba+2CqS/5bjEXxZL0Njrady
3NTkAYEUmKg1/DLDecy1Mjj+G9Ixi9+TdDW3cyWycGtgdRKw3nI4YaNseTiUC8USTqiDB7cAdGlX
MDqcsf14Tr5b1JcxTh20EYSfUd3UfyrtjVwIShFa9g5iOE7V/RkCy+MljeNRrU/9+LbU+7UoM8Q0
Lb7ee1ZSF7VmXsIPoEgptxA/bJyTl/KjX0VdG3aVkEY7nxx4ZSDgPIgfS9hWWmeNDJ5B5Wl0CaNP
SouSnQymT61b3EB8XqpNuDnqdZZo33NfU0xqkX9cFiS32Jc40HW6ij3U7IJSrHfznOhlUQe6Tg2S
1OalYkJQf+eAdA8NXJ1Ur3PsdDGyAviUYSPtG4YKLUFPpUZSiaZMqScLIgw4hECan7fgAmrMBWgd
/5yvcEklHnT3NRU78CI6TFGFKeBQ6FH5Eouz5/6VewJ04WaQpf7AeI9qIKt9LYn+HqrUX23YloZZ
sqMIAkYoEheLqgC4LcjK/MqdlWCKTBMxTo6hrXwOTEfyxbnE53u8V0Xdp+xafTjC1g35k3qjuRzq
67Dx4FOJlYW/nteZ4RPJtBg7d0TJk6QIniF6rYNx/YO8Ms5CZAhfd+aK0ur0Ng+yitVV8uck6B5a
t+ea2tvjXGcs8mVU8BRGMGAryB7ekfFS4f3YKkYEXicvv0XSMaityuAqqs9RmL10i0IpuA7XnqVc
YXlapPGYQNRx8Ik2B+Gl6oC63O4PRSmJ1vyjEurEIQSViPSY8jFXoCrwPq5IGR7AzlllPDL/GRWf
H8uSME8w7bG6Aphs6NYDjXFwr6UL7jsUz344xvHql6S8h7E3Kkehv4w798xQGteCmHLJpERw4PSM
nrxdFihoAuxqJMrflk6JSk53t/29t/47h3o4RY39iU2FVMwHryl7IPOtDiN40+54e/TYUDsLPRl1
S7wApL2RdS6fehvkuMwRZWzX5GioA/zoP6rpO9UuqbJOAyhjHkPEvE2qtQlMU4Q2FS31yXOG/n1J
AZg3cxpB3q3Rq7jOdhQOZjdpxticCekTvIGRPVWY3qei85bmyNu0JwDD16JDOjkCdoqsxUjsWELa
Ys1qQx2M3l4PC+Ts/PVH3vJ7T+XPjZvvmSekOsWA+VRBR4hb1JIvTQU3KgG2FFnMwN1dE3vlLN2Q
qUGUsayp2z3d50+GwvgDC3bzfzP4bXoZQsY2kCxlIv1IVqh1cCo1ZtjUrsgrOPol20Qa170vga4W
D+0U1t0nuyXW+osuywsy4ixMfmTcJyj/oG/Fp0ZVChuAoiQaglXE09pMr77bQ77vQM9wKfF9CHPF
1X/XT4PmtuiBC4bNiJm/PnOvmB/I3u2tvBf2py/5Rnu4HrCLNodUKlvgGUQmHVrKf30AP5iWH9kI
zvHMg1xb/UllnIa1gSYFVIbIfUpPAsrOFrX5xWk9ixXFvdXXPJ0PoyfVjkSeBaT3Zua3lizqZ1DT
hu2EsLL9Dxi4J5mEaznpYILIdId1FV2oHjupO/8hOx2Uy+6a1g9tAcUDI064EDoxR+JS/p9m5CLL
31JliWrs2VKmEHlW/jh72vKa/x//paTCBIKhOZy9QihaS3uaQMxCkSSRJivBTbOCksMuTmKKCIY4
4y4zXiQg4PVixem2UEVbhSeXveUgYiFyRzOOClG2TPn+oecs58occ03BTayZZ9XnnFGD3DqZ7NRL
HpziYhYsYPwH2LVHlJzHZifMQ833lnJlcv8h4tOcmWy+yTlQ9ELDB+AgFsHZa3ln0YPVi1w4Uy7U
OCXdH7gTzxqgqk1Si/JUQjmhfwAfpftbpFJefpZagbV5vFIYCj1CUgMksbC1AFdaJs4PEJR3sWnW
+54xI/4KmZpuoqyGVTltm4NYTDCkGiGd1VGmJjzqrNf1fWlWvtngE4WN4iTxlnQokr3vtd/JxTYU
0Li6gWJIj3tSxVC3055Fg8AsVAdIwhgOGakukfCkDcveEk0f9wWjhxLMwCQ3ZC6dpQ+RRvpSf6rv
0LtKDL71BRgYoBgow8y3rQZ8jZdZ+Q8CpQSCIGGWwmhF52FFnQfigWUMAO6ovDJbRGPUg2OvhOXF
HQnwqCNqrR/9U2e+JrPv5iXQL+TKtc2QDHOwzIUd+ApIRc6gWRvVhlmyZSxNNTgoveCgat5xHnKu
hHium8EHKpJEEh9s7+ndjeyuxFb/OQlbLHTmccBsZxDnR0KCXEVuUfH9avt3P+fFsdT4olhPIlew
hGFrWBPed1dnFw3RpSxMLPGMUsaHAGUfBscKAyHlB5tg80m/qKBiCbxCIXyGQZkICLADaZMCaQPJ
6dMOHXJeeF+HwAHOJ1NBeM+nQaNCfPwuM6qP08gcP9OW2KQ3xiWQmp0qH5pRuLyNnxuGGN9RaB92
CEvbofv77Yb0/pjFRMZz4mvPHUd5eDR9OLVlj1yDP2bYj9LbgjXe8zEiIjemm/1wobfsrWeSOYCn
o8LhBfPmoQxiP22ycYlbyuPTlE6FDxj1jlutuoCPtGyJDSDyW028oe5yCIXY1pKkigljbS767yib
tD/qjtgJ5kRHG9EbbE1rPaJ7oZZBnp8UfAlfZ+NGC7Y8gnXlhShiZ9PokhXs/DP3nWmWxK5kSTPy
xrism55n7LI8Zoj2OZ/A3DJDIcyWFDI/LYnweCxGycYhOF1wRDzZfYwhNnqxcDNZj/UlWGN2xAd/
oiECPJdOrEFd0iVd76B/1Z76EHwJBtXY8JcA99w+BbWvbAhNoUE2nD4B9znQWUdgTvdfyxfopx8H
QyASAmFoy5qmVbg3SwrD5m3bPk8GP2T72EAAyii/BudeUy2GNsJbxYFHNd/GIhjdlXn9x/g6gSOk
KkZzKW1aVp1E+wT2jS8L8J3tAlB0IYKOn29TYBvVO3HNP7QemlPH8Ta5Dr/opSUnW9hfPnJbjK0k
PUD0cpBKVN3Zd3SQ+rv5IquRfE8YwIj10hXtAVY1s6L/MANdVI5LdO717FLpzwtKfsMdAF7QpF6r
PwahCmESXNlo6SONzMBiIzVLYxGI/lvHtQx1je3xoTD74uDYtkWwLE+u3GS46uKegs9V7FTmTXaH
bZbYyhgjOJtr5fWhVPNvwr13yqlbDPXm4bNaegUcwm58+bmc6NDmHEQ9Y7FVjAYyUa7XpgENn4yG
U7HwnGZNXA3RJ/fZ7mGeA/b+/pBkdUPASKO5p4DTPRebDBjGea0x9FW1FyQ3jvubjR4uVn/RqUEH
KA8a0TEDTyMKBaVn8Ls8rRxVrj3SY2nUcRxfhloSzEE6U/oRlXp6Sg8DkshH63uR+AlbUuYynrrA
H+hb55G8YjXBcGSpYW2oc4vTVNswrW/aNQ07PmEjJnxW7/W8LqxdBB1T5MY8+KS59C+rRj86tJQn
dUL2n20SZ+jFTTw6MO9on+qdn/lpvSqyXjgvwrodcXfuC2+0Iw52GSxmhW2FZLi19EEx4LHiM+Tr
YNNZB0Sjmk6yi43aN36ISr8b9SpgV+OX2hjzdRqguZLcp8X88aZDDuVygQzqJ1eiuzlt3DNNQc6K
9wloVdbJxPrbEDnN0F/7yfS3fUJDdTUjIv756Kyq0mtqt2iQUC8z7w1re/rcOkBKHG9rP0LWawU0
yKdL512cgaj+uDM/W5K7/vWkusrOQhoZp6w3h4R90KYulIyy5qNfUNKQp5KpKgjTt+Y+pxfO1IzO
CQTTveH4w58vp4lbg/6Ktpw7Q8zqHUcJWuSJdfXswB6w+bhv60rTOk8ii6rqBeqwJSV+SEJhaZK9
ISrLUXdXJo3Z7xcSBjFH0O3Kwf8ZYnIsZA6nRoCinpLq3Ure+c+VnSGEAeTmvWn17z71kHIxYpWv
4LuvDWOcQE/bisFQYLIE3xXO/udPcOA6q5UdpPkD0mIU+rq8PsKpJL3sxxicl9lKuY557NH402eK
KV3gAQOzQ22H54cpllX8d6AXw0nloAXkm9rTIF64kO5encO7Xj7Xy+VXSDTe41JjOb8+5Vu9I+40
a7tCcFRBmRCVhPwjetohFnbe+tRLb0EyEKs6w2Vkmp6xYEMAX7i/ZJUFP7sBiwoa1eiyrSL44aF2
q+HIHIG+pWpQvUjCDNxjIfHuTG1Hqw4M5Z0rcJmuVetwEldJZUyoovKr/IxQrqgd2aS8+cIopcu6
2k+xuNpQgCwS02XzXngl9rDNfBaA9WhMDux4NQ0D307z2GszzeX0+9TLbwk00BjyOZ8hkYwMmfIL
ww9r3k+4TuvtFtWqv7DRiyUHIT/NSVMAcNE+n3GzqW2A0KkTLvWEyPD/HAQ51kG4rCC2m+YnNn30
eUkhcwY2O1xMc5d55cFDGHVaMJTiPdUYoHpw70E29zl6TCLo4nxiugvFao+XFOl7O4hxk4+f2aq/
aUJekVSvbWdJQ7GBLX77Zh076XkI4Jzn+hR41blyYOIObrePjRJq9TKYG15jEO5iARBSTcUD4TNh
4SQiSqmLbyxcriuGwWhf5vmjr/eC5oPhYlmb885x0kmbVxgNSzBHpPmrun8F1389YeCh2LA5MRkq
Turmpf8SMQuLKgTdUzCkT3C7SSghO/27vj8Zqrs4NUalM778OxBTqUPcupjuMgqwxhKSUtxIPxzF
5YXjtI5Zd8kHAtdvVDJFHOPxSR5RWbQS/nz7eRqjMvlLIV9eloJ7ByiZdVXzmZ7DOe78eN/KESPu
zpHbYLDdhG0OH9ypC6wT5kRsZBTIoOeZXN2WhsLIVol/acjST7mp3UkpArYk7FOkzMNLsXxvXVvw
A73ppyT31DrZ/A1QQ+7eYq5MROPJSMSwvQwRskmLeUk9c0l7NwodNryHQE4QhHH7HWtQHcHsdjgF
6ldxy/DhGXCMs5TLT/6Znt8RMt6VXaBcu6ggWupZP4tyfePaiXeyDidWJhwIssRNSBRWc5WF48yb
qv/u9DggGTOz0YidKK7d/BzLUIDGjIypTICgcykAcJCTtCJRi406Jy9XzSrCZHuABs4CAB+P+IOg
NfZI1FxJT/MaRbLtE9R1klKzhQu9KHGzEBhtfuWOJYxC6GstvshAs9BmLYrDYn7/orwbXuFvlMBn
cORNK+X+RrxzmwQgTwEJT/M8FEG1/sReL33UWjF50Gyx6IlAOQTZ8PbrCFsAMidngv6p8Rr3/VIJ
tTs8HbJ3SuRM4yashoSOoRHIm4+kdqpKAHKwRQHvBGvidpc0HCXKFPieiKrtlYyi3rSNvErsh6uk
NmaG9CZ260vO6/6dZ4Oeqe1FjM7G/C5vhDEqAbvAu9mYxfJ9cIZOk1gcaTZdTVSers2R2lJWVUmh
QrK8ToI1IvWiaQN/tWGuwZJYA4k/beWniqR9V2TEou3tc2TusvISGnwu4HOuNTyGfbnp5pvQIs2q
tKbTsNvVbd2/P1shd6MqyEeKsSOfFDgZhST5cuCilJmB5nAVDknuC1UOdPCtdegS6KfjvikJ+FDG
R4Sp8fdwCYKmZd9GmpXtV7xhcBv0CHnKjJcmJQBWpM1OxIOKy7De6SBJKH7iAm555vTY+l2pADWl
dJQ7CI5r13XTMm4zOVk0AC+8jxmItJkQJJl0LUuUXSwoFm8lKK0VS2qxndriIszNSLF1LWdj9KnH
6XEd+A0W+yGdlsVXghg2H5G6/RAaNa9QusjzJTVmFLYUhut+0hWjZXABPAdfmKLdAPTUJSiU6+8o
R1b+qDlvUiFV12nnuPVdf8zOOfORl87f8KNLmYTsdCWCtgiZv5yJZhKYzy4LbZOaFKzPZng1P/Jk
nWCbm8aOLkQwNBFw9G3s0/FzT880imBimJstJirYO0tyOdqCceEj/CV5o4xxc4dK+ubilAClM7Cg
KS9N0+cnNjz+p1N9DsmSugUbjmgpNLmOdaX0pY/mlq4rU8r5DoCoXCd7I7j4rQo2lFnaK9wiA2Bh
sjdxqUy6rp3PBWne+KU5l2aAfEos0tI8gDWAAYOXvuov+9nuag5BjYT4TAXBWGSDIJTRMtkY9gnW
aXDPZALbvRpswEgMqNPpmgDRMM4TU2+9XLo+N1WBNogmUBBCR5KNoyuT82xgf19qR4QxwkvAdrV9
uUzuDgM/tcyV5zZenzj7nMDLNKjX8r1E9ijRl7HAfRtWY1qMMyi9LfHXnew54v+XgLqEOxtItmtO
9GVRt9AReDpr4rgYY2XBdHQE5fR8G6awIcer+GbOe11nSsJQz97CW2g5kcRfhHjjALdb4a62Aha0
bhtBVOl6RBc6IzrQsJiJ5ew/TNGU4s75vknmC7pHzfx1TwYAS2GgwwFWlDVJyrqvjd8GlfjLb9Li
rqGA99LPqM7JvEjWNcfMxkRXlUAj6fgir2EIDOUX/QbUXk+HtMgAxh07gMxwPZrzvUX8KhbW8Kmh
plp5yP9w/SF6Q5pgmlNYDmEqpPSL/XDV+lWPm3a6hFGBh4EwDSZeppMu43P3cvUqzxIV67S266RO
ssvoJ3A+hg4RaGRdqxZYT12+v/2uinS9LvVNzVwos51vSvbhe3sgBonIinAeFNq3c/EQjbygQQmm
3JMA4TtTTRL2cxP+0Im0Ts38IUQy4MqOR3+J2V4R1Q/+PeORO0uW1S+PkL+4MM+v7I1ZHAeS6Hi+
OJLNXBlioLlGXwv6F1iH+CrKseLbLMUD7hbVT2fD4SqaUMeav+WwrnrZdS/OUMlvTaYlNoIxkVrD
MAcroooejn/C0lL8Dwuwz0kxz21G6mGRbNwSZMWGrKcSbCM/enWG9uYLCvcWTbxt5mv3UT3WGvFJ
MOsRE4/YnB4bJfzB+q9DYfsTHlCmObSNXUW05hv/6c+L9uipSeLAB4/wJKaevlc7v7ctmC0WJfoj
DLDx9kvMCybFYd4/nW1C9Ku7BK3weZWXqeU62Ag2jG13kPG4Vfd/ZweF7/Twi+wKbDWSXnL3eExD
hwXMWGvNxUssVh3sBV8uN2MVqIaMqFaS4RG55wS8oDa0HxbJfdV7cDoBRI/rv6NnXx15Fo98eFtX
Y4MHtR8WL32pdowJgQsawJrBdQAHLy5qpGHEqqlOsNW3krNw889oI3E9zK3V0b1xdLDH2FFCVXEs
ujwHVwcblVaBWgbn2lyu0n2A0T/me7AdnTCQG2kwKUrMjEcqV9Ob0a3HAKQVspES8eifaXsgpDjP
9Rsex2qpUWTFN89I171K4XC5yROVTPloBfNA2tb7f4EYOC5sEuAcXDZsjOaa3uRKMQPFsDGh6JeY
ZG3xDoVpXk7Em9bGLUhIsIG284vc9fMGHCKqdCbCsNQZgHm/hGgn1LhpFyjlRg5h8/6LAz3wp4+Q
V8jALI4VLkhMM54tpn0ooACLr/8dJhFbAKxu1fEQdX9M6o++Uu5XG4uJSnswlG3Uqqo9Y/0BCrYv
Tey4zmu/dJGzyKyheX+H0VvLbCjUocMXAzJxnw6tjJiPT8pMNGhaff+n3TN86Fo3SAFSXprOYCWD
9lTQ3UC+1gj7aaYRxqTL+rBgGjFr2vbr33o+5qvII8BFhlTobV2lwFO7qlDHvQ+secAPCcIF7nXT
1xQEEca6C3mw5GZDA0Yj7iZoWSfNZXS9O8mhZDTu9F5MKGmUHKG4LG4xhSB4RQ1zbVY7kbCbfslq
9+LxurM8+SxwQTPcxJ6Ei7fE3EBtgD01avf5CoLhuyKTzlEA2zSyJeaVTKPLi/kLV6c4IkSSQW6Y
RpbAnzqSuO6/sDbU48XBBcufRS0yU0avEDI7BIjPi0pvOCxT6yD7jA+7gA4deX0k+g1Bs0dZQrLZ
nBnm4bIxRY7GDlGCgc1w+Vz52Eas3OMeUb92bkGgej2sQQoMWeVNvR85LEDL/F4H9OPgQsyAehg9
sVmxmcqT9M8Xlr2v6IBFDouXD+rF3oo2+IGnR4tNN279eSCRRLyF7ZnWDAISsS7VuYEnZUi3Y+ji
IamZD8C+gQGbU3HP5qdfcGKql7NsTdLAuU879N+WltQ7Mb+yt2oETI1eIcluml09MEUz4PuEG637
3qFKR1GTV/fpq/L9Vb1jvzDLmr/4OIHe66Yvc7+XivLES2Vai9Qr4vBRwGkRZCDzjCR1yfLqKS2n
bbwlBuYRn1v1lTDl6dshTeOtPVpRGY1HEXUcOi39uZgMKo0RcpuYNreQh2EDyMQpnV6B/1W7Dlx+
k80LM843OGLvtw2xaW4h+fDjX+bku6Iz4jYoZI8LQlfH7fj06btPpDsWWq9InpSoqM2tRKQ4Zhh3
/rpBj5h5eVTsYEkDVye6rfjFrUXnkjp0Q0I9zU/xBz03WHVFiIEmL5tF6AeCO8qbnDUSwc3Bs5lH
VnM5vpvcmpMda8udG7YvhqMKJciQFcTgPgoCgYSvOTBsrx24xffVP92Zjt9Y/pdq1Zt3YTSr6NQq
u/wS4XDB95GM06UYe/v8DqXCGzrtO6EZYknu4We+ux9gUrbcbUM7kYQpF/XUonkQc4by1H/GQXHv
6MEEKkwQf13YenVckRmncVqQjIMZhX4wwN8wsKAsye5Zw6ydX2mfHkQSOmXyyUP0NCmvP0UUUvHu
xHuHanjjLIj7bFF8WTi8WJ0NzuVnO9WwszN24ONyiqm1bfnn2UzV41gkLTvwAVWUgbBg/Ltwgthj
KB07oyCPH6kH4N8kZC6klIdLHIpmwcCB+wA+kZICwKxD7LEdvHpCqlOon9w1kXG3T7EuyrwViUJ7
qH77PhJS5vfqQmOQKBwYib+M49hXgzZoacgh+AQGxeYiJXt6m4hqSqs4BNmIqJgzfprHk+M6oGo2
Lm7pqORUgAPE4wtZd91GVDX+vPqaAJ/B8MMPWwHS9P0G/C79psYdsqOwsuEZoCz+sFYeYICJcHnq
LgVq5EMNakvfW7hdjrHGULmJFemjmh8p6m6LcUEEqvb8+mJbFugc0C82E3NnDDN/NY0vaTkr/uVv
JaS8JLLh9qvJ+fI6R3P5OkFXMQdTHVITo1TsFJA8/WIEnCnjRTeYwy5FKfwGUgygAS/YZxnfyuPG
iQkt1hGS4rLxqzRbEGD4JwxXark8lOAera+ExFMCcsspa4ps2/0Op1LE+iAvgoIlhoiDSn0KFFM3
xuzYGsl8bNeUSlhJSyPZSOmzscdEsXp5kTtHNmNLhhCEtJE/j/zmUr7YLvnseaYaiQwXSDZBUwQV
15UA6q38jQdxQd/KB69RdqCNL8wrJIKbeX2+TrwbsZcCV9iZaBUl4qqryxNSVcMNAr1APoyf199E
KYUeInHvYdcKRWG52uvK3g7Y4FFgvmI9p7IGXKrKh/mo36f6evn64mRkWxelxIAZLWDYyCG+5ckv
qUixSH8cx6ehz/OS6Zj6nN7gx/hpKXRrquyraI1oE1duZm2gjUjBG0QKbp/cduD999MyNuQ36wX7
1CDsVNfjy8hayJn/K9HIzPx/RZheVbrWJssMYblXZ0PMqf8jqUi7NxAhGzaJ3K+NnwUkrfFH64FO
Axpppc/D4/MNLJAqCFcZqeJr0DsYe21gN/QynBBEI2/ZHDbR1eHxVdMttH1NIbkJI4DjEQ/GWMed
LaomjmWwvFWbetFpdj6hG8jNp4Zq6+FL5sQ7PIhdQhOz3l1/kqv8/E4m6DnYQ/o3iDdSAhPgcDfz
uwL0BknACB021yQD3LH7J8Ok5F6b62OvN+yl/tGMKMtLNThjg/awf6Tkqo6DNfW4QGxUPg06PLr5
rFxXKFuV637BRakXk22kzYK1e4JjlTsv8/3KQnAckPsc7cFTzxCxjQtoNKVajA2mgNpcjkL6VhdW
c0M/VKtZSbvRrlBv7HEnjHoyVT3kfpdliqaMZ9blh/iVWHREvgCSGuQERK+HHxWKs4hjAUVxGLTQ
dSp7Fyyuy5uc/MN3ROxh00/94mBL7Re34AjKRN/GPE6BXVOrtjshXSnHx4xbEWKlx5BGLtgTakoo
zRsSNSXdLRbs4PR8aLbWDkruFtFjpfRWpoakZGmEB4JYS2OiY/pYOrT6S+ZhXTD3OvIWax24h2do
pWgHedyM0B/RMHSDZOTR0SvHKVsZ4VwFIARl2cw+9SmF7ZO1dD2xLIvUMpd+5Q3uFK35ORqBozC7
Kn5r5en4TSv+gk/ikute7cxoB4tr2+ta9j3BD/SCSZMU1zeyvEUt7fpFAPsm/qd3Zb00w6YDAdGo
JJcwW2QC7fumPzSP335Tbvt2bFvDqUMXfHgfIXnwcGKbVoL1UQaSzuH/6Ug/TKymWTvxod29Og8C
/Y/KRVA0WJ75Oj5Uw1b799x57pLaYy6iDoTapf7qxN3XEZetJG5KQrGBTPxtV4OEkWTcAIplqX9D
01DyxetKhhd5HysR7aDSkHf3VCLYEPuJVmmacyO73cgDAkniCgIv+QYC82bW8ZJPW7fM4LAst8eJ
x/rDPww06RpRz3waTeQgrPFPtTBV1ZIZ8dl2l9ErmTv5sOxg9qZOa4WDGD5DhuhpJAsJtugYA+EH
UKffMWEhINI0dB99459lr6ceLdYH+zzH6yzYhzca74uvUCfBMU0usCQpWuPVUQbLLQUewwzqTjkH
BUGfU0zcadBJ3Yj5AWAsoaSeNMO5yOH0apMTRwwJ6cyAzK/lPS4lP5mfrNuncgMQbSzH7gz9CPAC
WuqJuNmHWt3Pkl9ed+lPzEFhoDRT0sOG1hAnKk8Y5P1JjpMaWCHMbmW83t4Zyl9Wkti0NPKDEZbe
XBUK4H6U6SuPWg7nxZvMKxN6KCJbSNuS0hQbylMiABqJ7aAro/TfjBQCXNDQhAf1W8vyVmT6PMP3
jT0aCLwjbCXoiGKXhSqTUPem31KrwVWS/PCnj2cp+mLDmbYcFzzr8pgRxV/8mJlA9ZmuqtwAwhGe
47PE7Ro005HEAZ8e3xvNAryKy8uJzRbHNJBwnTCuvm5LrZtoS3a4rtlL59d9lw84vp5BghrdA2Ph
zp/wJmzJstOKa+s5Bhf+KOfuaSoP2PZjnqc+IG1RVRENvYS5PqwQCUQd5I/kHruGtcgeh8vcKRHE
VgUstFA8wVEOdzOju0IryUZZCJ5ZozY0+5ET/Q6mwDgbyugkmtcCU9xutIWs/Hh23u81TnITpTG/
pS0MosFUK45snlM9HsD6H3a2d16bdUtJ8jkIgW3XdNh+YvRFthY+qFb83F9w8oviTc0XTi14aFwf
2WwTu590JNiuoyTJEBoeY2674AnErHVjzhF8Tf9rgPGV9uXgLAtVYSwZp63CcgvV+usrxY6w4Tcs
s3iWvglDAClua+awYLWbak0EGQ7aL1B1mKqIAPEjDSAP/giT8XDX92LhxhjpFzazRG+uRKJsjdWW
eEXgAWPtfVkQdHxphgDt9Njz9h0fcvDhVJdD6/vbQhjgXBPexNh6EBh4SrrcsIWq/OCngK28tfOP
x5B6JkhRnSdBsOn/xNJmdgfAQZJyx2rKRERgaaxYdWPhXErF6kscNj3qvklL/Pwq59ZFalVQJFKw
VniMR45DhR1FaLNB3MUu+AcFuodoCa5qj/SKi+oFofaytCsQFdLL1hmXJpeHGKPYVp6oSLzGM+BB
79KYJjjCkOyxI30+3swjAXGfea7pOLgduUsqjdOJty6nXU6FeQJyiybFPOiXHLmYR3eG/n56W6g1
DSpQnX3mXv2s+qHUDxBnZFGjs1AlO3qaNZr7KpSBjb0jQAtN79F78wiyuLletTVMAhz++NDUqfq+
+cY/emb46ZzARhqEOwoyvefYD4FvUXeKttaDaimUN0umenQfIq2MVy/WXP1O+pV4VGBFE+rCX2aG
D8fpHKsb7LTy7JQ5WQh4OXWQ5r/dxhXbNX4+FP0fjlFeB1nmVpFKE5pXBUctNqKqEhHBzjq6yfQs
yWqtiM8xO1NEH/xRNl4wTmActtQGGbOm+jYKH2MKQ1s9lUYoTFuk5D9mkcf1WQrjIPbmBmG0fmsV
p2wYQ/IhSXF9pJnl9ztXQttaB5Ih28nzTlVVhgkg0vGCx4MPzEdIoOplt0vvpIgwa6ZN5x7CC6Ss
OSRbf03q5U5TCGp2ZeFqpu6Ii7qLjGs1OGNTCRadWRuEIDhjB0jEizFvfuH+SR/Y4LEn4pHiWi++
x1xnzuI7hdbIO5wKpx5tVa6FERG4uuu+dfjEUPu3CmkJWdQEfdgb3DafCQ4+9ALSYUl9prtdf7yh
2kAJCcM9gCRLVKvDhnjqSQN6xxeu7BHE4kOrUJHVsgdGZGE77T7nWAqbA0WXTwMOP0UALCftR6g3
45t3TJHyS6D3RQNn9g4lDyJbFxwdHSY2QAMl3kiZHzpI1hbjiVf2nv4yWypwlwFoqdZEqiENe2jL
R7hhbD2eDD/r4CpsK9gFZqpGf7rJXnAd9Tp1x6RaUGN7xGW+VcAM8SRt7IJkmnELiICPgBi86WYR
BCSvlmk4HIn+horr9EIZ6p8O0aqsecku0jfrEawxNvdMIJvzIFfNkfi6lBrPTL0XqKahNhU+B5hT
Q0Bptp15LL5qEfPeasAOdm5a4VdVWzXMaHcO+2JkBeuNFoFRtY/hQBkLhu51/z6XCcxrfp1ZpUOb
M0Te4/bMBJ35X/RlnGw3xvlo3iDkXGorBG9kuED1Ssb8zqiK1OsUwpi4K6hKfpxcCNeMTyMcbqhZ
cg70fY+yq6+hKNBgMaKcJkv/75nrcfuqn2U2tp3hXgMzQ0BpGW2Ge9q1LhH/Uym1eCBoNvagusqT
u/5n+HuuMV5DberGH/NebkF7QCqaeH0ohK7gqXFdOVG2v6JSqPx65Z7PiNMABpIcDpYBMKb/MwTi
XQMEzvqXpxmZ15bIVfvAKI2Xk7KgGH67nnJ7iM0OTrfBUERrQGaodNNpBFHvdbieQRc/BO4xGaTA
Jo0DnIGMNbXk3Hd3EMObTf2g6cYIn5+xzvfDFO2x33DY6Vs65TpWrU9k3vc7GXSFbOuAOnZjz6k3
xmHr63YbzGDLO+ZQ/+MjqqEIqliLS/OxFMJ4FYaFPZe5DEV6tH7emzXisw5DwjjNZs78k8/bRWOJ
zKdifPuNcrbKpNmzE1tBGBhCNrkcwCp3v3vBEK3dIteho5PPLWGsr1X1w9/NCeEeFjaQHenDtAai
WYqSihwiJE5n0Z/UHA8Adx7GK1wKn515yDF7lE8V6+7V16ricCBW+x5/IURP1YG2E0vEruJAbIGX
3LJe+znpH6K4lm/rVFaRPq3VYgQqjS6OgXh08HglsNHpoal0M+yJTQqxARSzzfjwHfK6OSxcyzWK
8myKcX8dCOCB2EAwLuWiBoP5EES1w26YdCTfPVwPnEZ9VstLW8xZCvyFhuGgNvhePilLuoKZlBrw
joPI6+fHELjXDSbVOJeoWWHsSdZO4iLSr7DLi4V09z63qb6AGzcl/pyOUDCL0HHJqQUQS3B1uuL6
kGoO2Er4qqbPFEs4xu93roEFP7MG194yd/TytAPZh4BwlIMlxKtppds6Dp5r31QQ0tEn/qV7p2G0
TH5bWtW1/yFK0iqKM1lekqTxh3yzzlXgA/jE194azPn7AGLC6Uxm8StBE/cQxbh/DmAnpDDEhTq+
6LaZJGgBQQVZUqLB/L0v6/gr3VKivW1oxkA0NGugMKI5Kue6rSCgnguFTW4g6skv7ST9VExgNgvF
3Ko2WcrUaSNtj1mF9TKMOj/hqWoaz9lJb29XR008g0zFC+tL3qzVdHyJTVAQGsdvbuXJWm+7yLpj
JkEBu8Go3lPhtUijBILrq+kh8Vqflm6nO2mp+9EQDvERIJZro6M0O3fpnoJ8UdW+cpRZOVtzz+7n
AO2AKL3iDgqHjjNmzubDlpWWJ7uACVWXjaSH3PwrxBCbN7s3mNlfJy6ZGcQmD5mxLpA4IRmJkhNM
ToWfbbDnUHCbKwAjkm53PP0DAyHizVwaj0Nmb6zipNSXhjF8ofXxUnkPktSd2w01EmwQec7Zo2cb
/Owz81gb2DLe8yz93HCc/B8YyntUbJ7A1EQxHjkrTgkMCwG+R2TKqq8Fd1IFkuPdLuD9M4YQ1iOU
evOGgddoQODYlUHmG8APINe3IUxAldmZN2fbWttekky/SmjEg7xdnwZyA6HWgBl/AnIydckTUOYJ
WIRlBznTicJTfEsA40l34BuANzYq8DMSotrOc1JMSWgqe0sdetpJnbXSq/8MgnxwQyEOlLhT3/lt
QETLrOe6gsCXJsORyYG8KgNdZQhlazubRl1lJ+XP4PnNpvb6dC40DJCKEADssujfq0Ol5lXvTH6x
W4uAkiPSyQJAcip0Ql5QJACxPnb5esncAE9eDrXhRgywIB1P7p+NcKv86eJNjr6WOZh6eEG5Qx/B
voYA9HEfJOtHwHwMOdQqk256z/+9Yo6x52NDTgPE5dEZyQ2FcB26SKGR5ZdhYjvSfaKM5UTdvQ1w
R0cLN417hBONT4mYf94HVSgtpeuWbA1iG/zDjrzyPFtzGhDzPEeU4gvrYteOsKgKEiBOMR4i2d0D
MXoKMi+SvWm7AMWDL7sPUSQ+hgnsDxmyivpm7EZAD5OcmOpQkG9uoa8rl6GXhpBRX2GXE/tMb3PX
+phVq75Eqb+trZhybjr9baC2qTxr6MKV/aQw6RqzPIuRxu7UKw6ehySfQjoSDQj0ohTb9c75ai9/
3ivFtXQssDOuJ0f/1EdWNnowa5qk5u0ItEsfOP/bwji1ZVQMsammKOjuHL1JHMNY/Mf/oYs6DF7n
sTCJYiGpWpn98cZCDwEc+zZWYqce+UZN8/ozrc3KsmRlD+CBtOQqqIlBJtWxtMWOhvG7Qk/eLFNZ
iKG3EjTaU/txPwzZf025MRipNn8wIyVWIHq6UA0+uC+/vbNAeet0PDS3gHQFHCm1W9XT4i5FHCW1
R6ygGl0ZodQ3YKVHZDjw79kSesV888mVPp6F/sNRULespfSakcKAWKrNlMV03UZ1POKfqlJMFB4Q
qPBwc68RnOpKu4lcgLbvtZgQTk/mt4PJJRwYzBxY/ewTctL2x7clHAWSHJ7mfpHF5eujU5uNYg6G
OYE17upSwtn8gNPsA6c3e17o0Nrm7csQu57eVwrTYSgTbrq5ySdLdE8MeHzbsvbDzr5l+uQqu5ma
U5XJblpVTKrBMnyJZM1qbMx2vbGTDY3i+5SUxTEl3tX4jZb6AEXicXH8wEBEbS53x0tSrakCtU2d
OCfHseL2+19GNs+/cCNQ3Fjf5vOevYrQCzf9QlBZ4kziYAeecDIB3MTAQDhfGUekr0SqS6vqgG8k
VEIl0sECqPsoecg4XfExdptdTbbNzmePyod0o7tnut8mrr08h77hC28Z3q5T1zJMdXVn3XlziCZg
BVkZrQ1HfqLDL+lbYuY61ctKLc7G135t5wIp3j1LntCm/jPSvK7TM6pj3X0KWD1hXG15g93HvHF0
F+6I4PnGTEjst0o8kQVwu9tXM6uEuN0T6/GxLtXbCgoJlUhBlkpYsjkU1/GH0n2RLYIVuFhbF8UD
cLiEpotagZKcd4d45zYgTM9pLz5JvTqJ5l26Mf70UyUmbL0+KM6XFOZthCtD8DonhtdQt7ZA9AhY
E6SSvWIHHCECHeU/aWp3A/iZ9XxvSbd2DSpfptugIaTAqb5fR8d81PcKCdLOy7afp7ouXlb/bzYT
kyjI5ehA78qiRtzY/WfP82pfgAcfzWgS5jKJaQhsyyGdik5TFZVf/furJPkB/hHnFqmhBdnR347H
advgcwq2Ury1Hu/JY4ryHKSNrBm5XIo3Ftj2eiF2Nv/1NkFUj18JQxw6JZJDCNcjpt4lFNuwB7LS
RwKE+uVl5l54fKEZKy5BnsuED+jblKmbJc1cwnLvdZ0MaUA+N2sZuOTFlX0aWK9Z/avAJGCljAEV
HxvfX5Ar3b+IAm/IkheKCJu2LKpvmT7/KJ3bwcDv3hwTXevseEBmU74sBjfH0yTn7jilLfML3XhA
ZKZp0+BeHBAJo8Da8A/UH+0GZ/B2XNCZTYbbbIjppp2V+7C9F2hL0Y9sVxwfhqNgEq5Vf4d4V5j4
BkhADNh0eoVRh94Z5F6BtohgcfMMy7ar8/dkJY5UJCmil+vaEz3WAtXLizr4Byn/WIbD5MQJX+L6
oxCECMd5waN8OpsaTP9pIW6PjiN5bpt2J0OlqZ9cuVYRbW2sh0iIVx0Q3zfRQQ/fNhj2yC1zhEsZ
627K22c4Xyf4cgRmLZwOTcfV5MaNct7xJZ/hfS39MS0LqzSjlKzx+uBtfAUsfDIb/rDYI7eqNZU1
ZswhsmU5xaZ4IUnZzJ9A7Ld5me0hV4Blha60MPeQXsDNzxQJdDEw0yVW666aJ9UeQ/6gtO681KKB
s8C8EY4H6RQhUY2cod37QUV7gjOPJEt+EaYziaNC03sCS9GtoqTMp6HJgJUob0VlrnyaGAmD68DP
TLsQikUzraoyUlElicl0DYwamSNOcT1f5JqP0tlpHD2F3mYUXOCXlDpu6SoXcRil05Hd2E3bkbXr
PbLERKFI04qA6YVLqG0oj4Zb3Q4r2IV64iY6ZhlD7YQ/jkDwyGoJSXPfLbpc9gvkPlloayEDZBGH
JILxjRsGkomeKBX47mDTtq3hNaQrv3Z0y3Jz9Vkyx44KJgQzfMx3BGhdIzYe+38sF0dLsegBszcX
ImIkXHqDf9UknJVLYGV9wdVNKE6Y/pIrSZuQCjThk9gU1HUYfjJYBPx1Z1BhZThP4gkbEowdYu4c
VFVHtrdXAM7xZ6YUi2Z5DuN3YCFiRmDOFQvLKJ6/X9Az5G/iQ+p7Kn+OiQgfcPjac+YLiXvGL5Fu
FjXCDneBL9KGPR3SvUgUj6pw+oliVo3mcqYn+h8tyGob7vBDIHJHNzJgSp84Ibin8nkrWltOqzdh
q2pIou0mMTykwEKd/LSDRzxjJgNrKzaEGwRBqp92Wo+Qse5nHeykx+invvFUigzpAWE88wgzkm+F
n/0UMXcHU+8TIsA/2m1GI95ntz+94OkVvgxBu+qZL6FL/B86rj1vZeQ3D47stTdccCKRdXq2243X
P92nueVZx4vIQHz7nB26UDwtafUD3FFirgPjVGlpIIzmhKW4WKkzjn72DzABcq66praKhArQSC6B
orDsgdyMlgO5BBfVsI7FQiptK6NGuD55YGsWZmxYd7dslOHUInUb1u1aie/9XJoOU7Pd0ZhsoJwv
GQB5JeQ+kCq7I9O5ByKVVyiLC9G2I6WlWx0OcAO3jpP0k9liCE6/Qjniw5xtnqjHiS9iWXhQyvNT
AlYb/u37z0yh1DNLuiqeaMy4CjAK1RyX37k1apwXcV3+jVhc7UY4bd7P+KlGL+6QHp0kEYBQm5/g
sXzND2VJApz0Bld1GQygStgfy2FanwQa3f3Ff/kbD6Tc2brsNTJ7nulWD44pARyvUReCzJJzMBGr
3ZD0gte1RAns9o1TYJ+sILQxeuTZt9FcMXc5gHlbL8a/KdtxiRV7e1LRLAOjqvFEe0CKhpCxD3q+
2/hjEnw3kwEmDykARlinZ1qMWwAJxeYSc+szaOcfC/KUL3nawhpHzLZbndIQioLj+N+96PAnISjN
iLAehBJ/a2Tx243QyDo0X+ywv2w8FgHz5VCSeqwyTnbG1J9fO5DuYxFj0ZQ5NANULgCKKayN4NAL
LKETjUmHEo9tclx39H0YJbv0qtR3205l1ifynPXzz5GB31y62JdiCCPPbsmYnVJN0WuCu/U0X/tk
8yMbrucEpg4L3rCXefbi05/pH20eiwrTRevTERUsEpd3Sizu4YCaPY9MttLMXdHAar8WBukgDjYy
YFOQXk1mjGEy/Fl/3tv3HncOJFDz1uKWdTD9sBp4kubAr90E3znkgdNTwvYaMLJ8XOWKme14WbDw
yK1/gPPURGBFi8irEazELxEBhHrxcIF1kRx2bwVKGaJujYOh05FDD8pWeaazsEF7/qyr7ClJWCsW
1cJVwHiWNtZPI8uYfIdHq7XieGix+es4Ja2we8JlnHcu20P9MH4j791QeTYFNjsfj3xE2jn9GI30
wnqbGUBboeguTHKddk/ErlF+CrKR3wVykCuyzP8oMNylWHImqjcxQXDqLamZrQMDDIasbtkDPp05
l7jtwc7xI+nOX2P8rLt52d0+LfSZjfEJhShAqZ0chFEyov7r5QddOBO+o1Ppy1l+na5fWsptYapJ
R9WYtRPoriP+v7NphbHJQGyegekV8jy8UGFYD5sWUlrCCu8ybogVtLwK8A6W0MFYe7MTSY+qtX4S
a2ypsd5Jm3gH3ltqjA8i+R1cM1JLEdAEbFPj3cwMZnJwUCy19P4Kgmljb139WaKsjM3VM9pkqRr3
f4m5s4W+3idtJWw6KGB/YsnqCnIm7mjWtbDOpZECvS91opMMs3oW9IlGW8RMf+FiWRpf3rqDwX/W
obeVQ5Uh9FyvsnXzElazV3LlfjlAjIDfFC7L1SfA/ufNmwYg6ZhIBklaNvF5mQxO9cJ7zN6LsI92
PIrpk2Yt9pwcbtOxwjy4lquqyuuKXy8qDCpL1II6P5vwKxcLt2gZvjs88K+xmGwHOVJv1w4WW7aO
1DFL3IvSHo+WW0TfRmMlU/JehpZBOF+KciZ/kTa7ZFYHVZuP+Cghk1/XvemHOtyAyxVWb+DUQDqe
IWztpUteUL2eIFP2ltZxXPYDO7gIlnIRrSLkLl636NfhcVQP49U2L//zmljC+MvlrZRID+ygbJaB
k2HN54LNnBMwmxaE0Sk9rWj7mNlSqHJ63+n0ptexjz2vGVpVv47G8TzSM4insKJxVHj4HKVAs+Qx
3KQcKFxImmr4/lptS3ZsL0yXmegrBLMK8RZMGnS4yyAZCXmmtaWzk/cFuBiA2TutQn3ARE3PkEJr
dcFf+/e78p3yY1IPK0oH06GTkOP86FrFkts6J+M9cZjg+ouQ1fPBqnKUnIEtecT9XFliHkEF0iTz
+NLXoLbpxfHiDCgpUL2M5lCEdcosLRWxHpRJcvzX1WSPnz9ECsG58wA24HurAtXM+Ari8phKx0E1
R0Mc3DwS4JkuIAfPtEF0uJxoCFYliYoQAufTaCQWJRa4UIDvf7zf9xmjLSoABZEBjUoCOkAdlGng
KarrGb8o0RZiNPYCljPyFbDMK0IyUf7sR/EdY0kKLIyq1pDk6FbrKazfQJvuZGJKt1VE2DHR0No8
vVzB01c+cugWI94RRdVChMSef6mWkDat0YKqap5DN2eMppvjOzTfmHq+iXwMj1pWKHkiuIGMg8Mo
ZnzXGHAgiQe4f1k7CD9zrBk21pC6OuGwHiB/lXKGjsIZ4evLFyy3Jope0zShxTRUVvcdYnegkYjj
h5gGETT/Wczo/2OLupydNZe7EMEB0s1zvX6F/ZJTNwQD05bRMDBUnBDSDB1Y/tSYsp5TV4/fS2ig
FEZNTVCJkiht0+Yn7i0QVY5Jg6Y+AEgWn7qKYwBkPIX+pdQmTTqaEW1dloO7pNwGm61QWR+BIxgF
fmjjg2+NlbAo1EFQ9Zbv3AaEaW9VT3OX0IlfpYiEzTrnMEA8lCGXJGovSFU1hIFd9z4NcHulD+0D
XEwfLcY4UeDCd1P7/7nax951FRXLoSsS91J8l1KivBGOV0p5kEpocJW0+NcXIhNY5i1rF9lm49TB
dOxTMFLMLvB75W1eS2KlSUzf/85iqckHzAAb/y1x77k0rIk8rUydJPD+wCyolVc8RF1+xLtsC6f6
pwJtqUq6w/4S5zuVfd0ev2WdBh7/HZ8DjUGcXLkMCJIMnsvE8UUQeXox1sxU3PFyoMps0Y0A243P
VtHD4KTMbYmhdmfSe9CWmNwHMw3uwkdcDSIjTor6shA5cAmRauBLhtFfZo01Kh2wHmiYcsMNzheo
HSlz2A+OId60HMYkIYLA4sOimOVa8QZ3s9/6Y9RFjKl3MSYLuFmnNVoqTYa+W0FGqgum4BX6OfzR
77Y2bW2qQ//qVuhtR46TUEU//SWHROn074G5bgTGdHtq441eRubA5WY38yvUIQYyHzEHt1qfhm+H
BXGJT+GWv20qW71l/OJlzstVoZ1yNJlZMxdfULT/E/fQbBNBl91BrJ2fnLl4UxOlD1rWKYJrQ/uh
6a2hNQ2FOKMCogVX0a4Ktm+5UEQXRxTQyo5OoSc08IHeq9TImikNsmt1DIU18elXGqMg4DcBx9Yb
TScToaq/1v8tFDQD7HxvLskZ+ksrW7T9XMnNTSW4DaYurBeepivsaijL+okB6r21X5/8MuSRtVNd
/vd5tvOoSvSmPt+6xpsYZtEonmCNYBn68geQ0KVIpAvbQKUtcRaQDNRqDTbzlLLku9KhXd5kguVO
kxxYZDHhKM2+7QYJawsTBf5ufJVbyVFPdLsoMD+Qq2oyLVNRALuKZ5iYJ3eL0n64yFY20KiyfERP
RYO16jOpUjxYsc5hzv/dxBB93JriuTiwMOWWiQOu9jF1CwpDGhWXXyRJrnnOJbWe5e8AP4kdt/bw
z969soAYUDImv3JmTCycYdUo+6tKnMsWq/zDlxmHwuomuZ1OC7/RDnA2zuWqB4lPK4k5RzBjZNsd
krYaJlIWDPiPgJA8ZZYmhKWs5SDKgo91AEelcUA0pxa50q+cDWnw+rWvmL9zyWNE+/wfA1swkNTK
Pv+y5rbUWJfBR6zzWtGXva+RQyu4x6N91kKkYOOloHTBb34cxgZK3g078imQ/PRDhMAMSzHGN077
bEavT8rygIh30zb8XtJevDUrN63oxwXr5/rh1a+aopXi68U4JzTsHPYiAqHqGoGELSYieyBUE2s+
dOHje2Inxyrd3waXHBFrHThGoo/5rpez5XPatk6y/m7/ligEBgaJ5bIKQHZFL3g7XwGJ9x1OwkJt
amZW+uDHW41gcVGs1UZBcFox3Rf3Kwq4BU0W1p6f2cXJ9SRS/7ydVkkq1Rzz7sBiXVas+bitOOY9
7GSlmlTgT2H8aJ8o3sabBykxVwp5h4V9QazNhbSIt7LN/LroxL2g8wIyHE54BtMu8XNAxSbD6CJw
e/d6TLAz1/si5SpupyzH6ky7B1xD7bf7yNW8V8X2wjntoa0JJ7Qjgu/VNiw9AUfPJj6pwHkHAhpX
SZAmmnP/4Tcwvvwwm6OZH7SX6FoHm/HBq0O4HmACidLQV6TihzrE61wEAqfexilTs1tkJ+AKqq7Z
bIX8HtZdsFS0Yv/EX6As4l+9sqUvHWYY+cYPB7OpZMIOqaMwA+fiTzYMa6Mxn3PDL0Bno5uLMIhs
/D0irjaa29z9oNZsi9cwwsNfoXijZyUPglUq8qum/2MC0g5Pp1WJ/nNenoehWcTtHhz2ohfbfzUG
siCHzj+DNtcWhMv6bB3+l6a8UNbvKxjuLPmZyTJ2V7yxDBiSsxIVgbUIdKqo5oe+frQgDzvXL/Jn
Qi5rYfoAhAJJQfVoLoCEEjjVn2yherAP6OtFsyjk9KAN0pnVGNoWFEYx0H4uURYZPXnfOjUSR80C
679JzeY27C9aHl8WkN1fbyAhJHPyTF4XjpUSuhYpRoZo6dxv9FdN/fGp+QPSYPdyDNslkk/RNO4g
PEiFqkctt5YSdQ2LYkw9oyzzCaw2QVfw5Kkv77cBQKwo0Ya7YcliQsTRWwzZm29xzJYzEjdjAVKr
P1PlOs8Fkv30cib/QHvPnv0eyQp0L2nY6LTTR55YNXLLjoyIGX2eqogJnXKWjnlCal2sLwz1GKX+
sNYIOZySe9VB9GvmtToLlhyxOFzrH78IPpTAUschSD2d//+uO0TfWyiEhCB/SlUYSQwXVbTspZaA
qIsIRH7xyA8jrwGF0UcsEdj1YptZ5kc+vNemsq12pknmtnwefI26n3YuP/sfXNAbedNGMiH2Agf3
Jea6uMR4rg1hlvnjP5geEJao5F94I+G9O6q0ADnEy03blvZoQ1NZ9Bh72Cc1NzNbV/eNZRBFL8KJ
+alQDyerxjKwgq/EMl5u9Q2bxT7Y/4Wj+FRosIUNy3o8nHCO0NvPvosXYpvfqfO0PE8MW4cvTh+1
ZtWPc5FAVtlOYBNaUJ5s5e28V35dorPaWmRoHyRsbZj1wH4nKWecTo3ePy6hKw5xU85DY30z632x
b7AtU5tMgwCax12eQoMmIfx5L8fBL05XoWtyu9LToBkwq8CRwZhruQ02ngfYn46YmbjrWp1ZsSUk
piy2CsoCAv6gn+GvWtrAw4St8Aept0m75IdGLwUZztruUC2IP/s4lswzDvqsaz1Ub0aM5kMhi+pQ
nss8ClAbw/cHG/2IOV+UwsNn5wrJP2+VbJP5mk6Ez6KyFAUtDvvzq4WvX+0faf8lxVbhaLG6/Tjs
wGi64xuagVHc6g9+xJqVmeylmto1b4s00dlJx8FQztUqkNMvFoZClm0Mzdl/FeHabLwznFobY0y4
xC4d8Ab7GNzMSsOgitw/c1TKzSwqrINk2yx0sYrSmBfBM3RzdQl2udrJSNPgxEfxMqZldNnr6t/s
3WGmC/528FVUwp4E+yNmEXtM+nzGMx74pCz3gcGqWnndcDJYditlvTYsQX8Cqfq4zYXMx3VUO0z6
/c0Nok4FKPqVHSF1YAdeeUTLIgG7IQitR3o7YJEVqSgok9k4sia6IM4QM2rv7Tq+F//x/YEWHXsL
i/+JMJkPpRZ/C3isdCGSjDWEhcbnZ3BjHVlaeJTRDZ1tWV2K7DDGO4l7eMUkSsf8XAzId3unChDa
B5rcdfP/Cpyj81jpJ1YEKLZcaOdfce/AdjsrwaU3RnvfdQRL23ZBWR8kDRphxUAj9e4/bn8gClji
7OYrl/uLhJ9i7/lcsDYzVicc2rTFny/9ZufWHXTSa7EC3wrQwkYRXPbUHr3KIQsxEVbNUIUqU4O1
bSpheFBa/GyOh3hQayAyNt5GUlyx7X5liD7k1YQLOFQ43czcrz+Jw+mMa4BVqQQcgxDvbd+XzkeL
mWAh/+nNXms1wBL2gGO3UB4Z75EA2aJhcftLKHTaVVTiOqO8hwjEKwGOU/Q1DPMrJXzryQ1qdeib
IrOteqKblXhiuXTdJG2L+JiSLvZfBnNJTxyE+3wVWVHPKa7q+1GaIvnrXSbERzXEFQ/1H9jNj6k0
zNZhYz5uv0AxtrLEa2GB0ZHu26zqsIeAXVLeqLpsFQgbC1Tg/I4Py5EsG/60b8s8zPcBskfjKzhS
ELxhD7j+ODHibYRWCBICz7eLkP4vuWaV7+tmIMuZIksapAbj3Zi6ucncTBzsN16ulnlUVInvx3ke
bhUlD4rZP6d4bo+kREvBxnWCJ26f9zkWmrX7BPeOhXsCF5TNyiC61nk2YwFiNew4UEWTc/QEp6oq
vvDbqCYvI/FVmBgEMJRxoUGrR54v3m5UbM5GwdPAOMyFUg9rOhNqykTuDSVxVLyzwbII11bdC2vy
MJM8V5mV5i0fg7xhQ2H3+NwevezrzjXbzqgPAK1guKfAjgzWXuiDOy9TzexpzXsYt19NkD2hHMbb
kxeJKB2fVJiILoDavmBRZavZUmZvFTOQ76tMJShJWglUjDrrYjQfdUJZWgMCRxa1HDgINOFKsFTi
s43HDmopvrWLtxtasrGUYS5STi/mpw71ODyylM/YpL6mfDdYrBcHi7RYTkfH8w6SEn+OldpmOvxy
L3EK4MRW+QqeNE+2iucAUtjnHxj+8I2YaUz+HKRFxZsfBlEZb0uCJB4cxDPcrylIidNM3I2BScvN
9QjvkpX07xuDKH8Bp99OcyHKo7Myls5dsAs4gBIXtPKCf9XBCUqbNKS9QL09Cwhr79ufDaRlzsne
oSWD9FiKwH6qCHKtpEXHbL3k8b4OP8eenNCZe6Pj38jB6jE+KDDg+bg5K4O5/7C9tMBqx0iKw8qy
CAd/6IWws5yFzbB/uFGrRdNdC4EmR0QnoFzDZ/+xIQXKUWwpzIKlGbtjvhCC2Is3Q+ZCin9BbP1i
pDfsepB2Ml8JcjVIlvFqIhiqT2Ww78oN++SEgbuwrKCJ2EWGztlwZa4slmqasvTgtbI7j47OLvO3
Vzo4AwID/XQxTEAyH612Maz/Ve3ebxKcsnhr9JEQXTNLFwc+fVuFj1rVCIrLVJYhRpFfR4Eo1a78
P/aYCJNSa4IRpwS/TWOu6JisihB+JTgjwqr1E2KlBQgNsveAnznUfZ/1MrkVbq7P93IG/BzJiBwj
jH7bCoKhZ0mXVt3/E1tuA1xlvoAspS7NHDnv7qAWhICwIoYQtfgUtwiwlmXbz6qLXsZYDg2T/I6X
aSHh7UlQMVnNmxHe2VCe+QaeejmPECZXzpOZi27mTm5XuMAgtU/gpViwKempQEqwy8bMAnyqmT91
1mBvoCBkDhuQTRBnbrTkKXDlyaZyjeHyb2zBhaklLGy48p/uCIN0AmhILglL/e9RmmFYiyNTU9uz
EZH0CUOAS5KN2Au5e95QDI9ANx3tAdMtNPoquEyePjuSk0Ivc3DQSG7dyAqXEeWTpaIssjcbPSj7
nbNaN8OSt+1SJQU2PIpOnLQv5bk4bZ+iFHAi5MZPnHgk2YszUEGw1oeMU20CPjLrRPEW7ntyh9fJ
RgkcM2mjnwD6yenAWYZvBXh3U1QgwvRp/Zy3xkUPrgmuSwgz+cStyiczU2sxFb0q6tJKagaNnZtm
PzkN6/mGVNvTucQ9Z0GS1NXBAUw7U614q3GYWzDVnZfkTPkIVQajJKXlnGRjrln6H1+xiq2YHgf0
h8LEhGtRnuwkBUpI8Fr7nf5G5ewdHGAEDLZOEfloDdAglHQ8xvlv+8zFB+RW9dP9gMFlUYnAe0+a
6D0Yp/nl/JDWcUJlOyctV4MfyQ3oGtNyDDxh7gbx2GiPwYnofAHk9voUGgFzNVX5RH8EQ46uz6xz
1EVMS4dPvnVztzy3X8ZLOY7oXbgmltnTFpTyC/MEz9E5G8byEM79kdxQV4Ez7zfEIpXfS6OS6H27
gBdH7TtwlPVfkWBtLTK12ikt4/Mx+dqaO4UU5mWJT2vCMlD2EC6w0vS8haP6gplvar23cECMnuUo
mD+4jyxrZSGjAfcCRP22EYLbANvr+3vwVe5cvjS65g+vymGymWAEBUWr/y0Oerxt63RLMaSE1/Io
1oLgK2eet3UW6WQAOv3moBV8n5Mf0YtNOpD02DX06xmE3jDgSuwvwYsUqa9Jk/VzLANjXdyHmvOX
zhPDsxexm8cwFWgqn/5rE8qPofpnlM69Qq/dtgCp5C5MXqRN3PelwwsciQD6Xc2sHfoUYHT+SYNS
fc8akd4r1pKSKe6La7EyNceiN5VwyX6lZewTob19kZwvW+4870ljfj0oo+Sup9ZpaaM4WmBPJaKc
ssdkhlYL73vAgXvoE6FTi0LPU9DkGvHHLQqpAQR+CAS2aexyf/A9Icikh9LvsEuZR/BNPsWsHiRF
lxj+hA/SdbzJ37S/Z2RuN1zl34EtCu2gHpovHokIkwvvbeaxMq9T8hO4ZBUsV6qIo2DvDW0zqkrv
TrRJnk3AN7Bonafqn2mQoWdqRUVzKxdcynazjRnbXStNPlk+bSSGcq3/OHMp0+gV8a89TS+lt7jU
glObbckyxSNYuDelBdgcJX7nscNF0QCwM6aj22ogTjY+wkEZpZ68a1ny87LYCwnlK2DSej4kZ0fj
WghgxsNr9oXMlCaXhsv0y/sbPnvaZ591xyOWGGO+hKJ03+FIhuPoKdnB1ohE9lt+z+CChEXHjr6i
bsd6CnUkGNJTK9tW+lL+lxkb0WxJYfNxjHu9QgleLgwHZZxNi6p3t4v7wf98mov8qDUkGQx6lN3N
VEqKXvQafipnxm40tBEmmxoMTtqPovs0XslKOcqZWFviOIHwIzFA/IkzAlNJ+vMq0pWGrZu7cVIK
smKhpnOxZocoGAgMg4pwo9GOsgAab2EZjt0pRz0XNrzCEO+KzpKNRjgnUuZE+2L+qkPDAIikTpUk
DcDVy9AdlZCOQhxOXVsloUzxPUC4gVJwQj6Ev3CFg6xyC4rWrLvdSoahfMkfS89HJirgR39Kkiso
hV+DHIhXkGY1Z9N4qbfSenwvVpSq6QGvo7huNRABbTYYILMXawS7t1pnlMSKSoIpWe9vR6xBod4D
Q6yEGbUHXhoOTIv4TvkSq0tAoyzIz1iPb+ZGNRx9Jkf62w6GCUi1mtjknuF1R75Xbm7CAkhQS+8E
5xPEVWAQJzW4LiFEjump6/YhhxgTCKHu1qBM25qOl7BvhtaQnv3inNgly2duSQ5CR+ICieBwVO/0
PXGccreB7VLwHKPEckhupg1mGlXjtbz+LBqFwf6DfZ4aXdTxjo22tkCoSvc1GB8h1trXjprGwzX0
4/FVmdsGBIVvBKuR/Gwe/vWa/ngUiQkFsfrOJx+GU/rpOzrWnVD4bI8UsiNMvgGo4vdyAzcyIAJZ
Cf7c0VAWy5FSUwhC2YWtIi6zVIOZiEbe+r5fisEIaRI6BgbjW5fPfDs30iHB84F7DNxEMML7P6kx
xrAp36BcTCVz2XtcMjjZboWlDeZy1BHv622n5V6sZJIPvltb+Pb9KuS3X2PVXKTAILByfNyaaGTB
r1r0zZyeQ+2nFop1J+l5d8xrZGRWFNiLJQRwB4fOWWPdnhgksm+JJFcfsdH/3cfYq6MklEWzjBou
VI0LIIGje0L68f1wKxkq8cGMaYOTBQYZtyP21UpT8Q0zODiUDAL4V32PToKVS585hOFVTAg2naqT
SDB6jliJ9bbWv8JI6CxC8soujImYL1QRQwbPvDDlMu6mk1500weRF/bmlMjOdRlT/naWLi0d77FM
YNLk7myumUSUicu8zpmbcND3hcJ2JSb5ma5aVTjMKshZxFgaayplRP9Kewlh/IDBPFkzRSHRgfeA
CWnrp+wBUcdNU2nDQULzeWsfqpadVQNjOPnPRErdDCJ1JIM9RrF2jXhZ6OLQq9/pvU1/4+WFL8Hl
4fngLsE/u3nrIWD5dtNEaFz7TBG2ZokfO1Sd/aRlJcWGf+N5KDJQiEUyJlcSkduQzB88FwWI9AFl
sOYWB1tvof8y91AIuBoEj4FWSEQsKW+sVEDiN5bUXExHNfgDB3A/4k7gsR+EA5LY+AakyXb1vYrD
ORHgx2qG7ffBZHv1G0kTpPXlSRQpkWEc3iYcnqQ8TH0A321Wz/RN7XyoP32eDySr8NVVQxJusBDv
mRxFvg1OLP6qINxnG7OThavAvsabhy4K9BKNuhRC2dik3pxQegtdLBsQy58Qj6UAkQyCzud8V7p6
O7btRDzQRxGYRaQOgLoWWyFU/87rEfZ4loh9Yl0iAeBfPLkt/Pjc88e8zlrCF8buN5S+HlEQoTSc
XfOj11n1IMH6trikE4jDZn3HYoAKWE0Z5+xwOuF4GVpjd9jzBzd82KOb96D1U3x/v68ExUtsci9s
BfTZQbGpBVG6ezCazyJJOMH1W05I9RIKVT+0Ls7ggQhg+NCCU+fugvyM+ZtB3Cx2v/46uyYv7n1z
4g4xoYwYySTgzHB48F6C9vqUYjhvO/7M1mFAm3YVHyqIM7glByaIXOMMmdgPD85xKxQ/F892MP9T
9sUYYBYNCRN4nqS2xN+9ZRWTswjsUWHn61JTV2vpU52ZeeAols5mDLNOvl/0w3a0XwQh8hSIgdqr
QEICu38S6f05S8FmnigoEP+BZsS/l6jeDJpqpGJ0YnvByVGRdj20cEVFE6sS4+DAERrGOw99kRBH
v3hfjpbzQkt6TM8khlAhyGHOQC1/Epa8eJNiCdCSSVK9UjL8nKnN+oUp53jF5og+54w1bqv0ObyU
/8S3mxs12whPnZ+0wQ9W3vWVQUXQxicuV1eA7+xxjXln2I9RpFFbqDJJ3ZxxbfuC5zju0GPd+/pO
+DPg1ESYS7sjcehHhE1BqfncbB51RueFzHwRPR+9iIP7BVjLQR05utEL0iJGEqTTQhV/WNVB/c4q
eAPoFKPib5c3lPNIKahe27rToeACIPAfPvmKxLrjj0BlVNKlB4lbbb3tJs4QJoDIwazsgYjU6hnP
iPrHlbIV6CQc8cCKaRkxLKDXXGpslR0k+BInAeOOJUSo81oGb6fEV2OJtRNqFYE+NkwqskqUHlvV
c22utYoQNCfPsB8/O2f37LDjxXB3YCN4bu5bdRARGEadCzJvlb6FeAls35yEG3hWiN+T4t2zO9bM
fV76JT74eKdglbbWLbqkfJ/WbDHi4QuiBjAxaMpDmI29m/Q6VFAd6ymsKuwWfEdMegBLqtb8ctqx
zv9I4ksiR8FXE6vewgob5x1ctl2c6dxpQqP1iKxKQauVr3ZcZV3QF9xR36ubeOfo4fw1GYNWxeB/
EgfJ/bsXTe8HPVvsPDwMvrrFyIsmwB6G6/LcXNrVT6TatZNbZ0TS3/TgPIFYG5su/nsAVDnzgYok
1gCVdvTfwqrxmrofhpFtp/C6mp37bY6nCOcFlIclWy93eN0Lli46Yye0UdzEUQyvYO1wT0yVf9l6
Ij/t1oHYTM61GckEPHbz08CVw9Aky8tU494wrEQEevQ/8Prjpoq7UZB3X3Qo4IHWqPkUjXrkWQKp
C3auZZC8F2GGpQsAiG5+KFtmA8TN3Hg4IP1GVAD8L+RgAxVT+TClOBLYdEgbr8Zn37Q56jbg6zvI
i/y/dKDjTsKmP8vQiVWuu8BitSXsGM7i07uxTmA5nZdl7+trtL0p0mb85aZZ7XzRge/XiXkiJmr6
wPDdWZuV4f7oUTWWy/B5TSKxp/s81As19K78HiWdO6IADj0BkpsSSM3azzyX6z7kcB54IB0VgVCB
To0YuIN7Dc84xjQ20wdSzmRhY4PVDh0lMzjajXXZ1F0mQ1RledvyGSNv+5pPvKICxaePu5SJUV4V
8mqcMwUYvuPUJ5lY/CWwZyIXwE0kGY95IRurNLi591D6ko0VtxYPC7KJqnOV50KZIUewNLsHiiIi
9EE5Kf9n8MfeTV787GMjB7H7HSzr7BFOcKg4hJHKtbkd9QPseOQhuTq643D+pQM6s0fcgSuGj1qq
qM11nbm/FAL85P1bpNRZU5donNi/ZbBNMpKGUImgMZG5T4O27nX4MXCAcewp0mwNU0bQNq/GZVKZ
TlSDctC1Zc5aY7wqrvRsCQKgUe+hhzOQ8RopeVO7OAIChATuBC2OzPb/Ml4HfEfMwhqWo529CaBw
FvQzihERkT6aagUg/qFae7DL7GV1+OC7n8YHmv10FAbcyiqHjLrwgDfu6Uy+RabBvy+HJXeXdPjj
FUtkXy8ncK00sFeZn37bcoJexqhnN8hW80IFZyqiNzf1UfvGCZBxdxUwpsc8ZckvFDHsjum3bmPV
I7pw8awYIkyU+cnVSs3EnfZ3buXYHIeDy/KXWQcLtE8BaZNc/BFam70ZG5hNvAnEqaFqBHkVSpWR
pQZFK/Vo4BfAGi/H6FFZlKVCO05e75seHfyxwJMzUCcsWoPFwRKDKmXbdajXewF0g+nypcpFlqF+
NRLDNFVfPczlPi9UHo35Z4PMSI57A76xdvPDY+NN28atUbmRlb0YUK/zcHuh1qu3drMaujLAKrkg
1H1/gJmQgGAfEn/5dIV2lkzu2btX6VktGZKZl9fbdd90C7PsyfYzbv5hfhjNBQICaYwFT0npAkBS
6qwQzNeEMlM7WZplnXSTnsGpOMfKwvX2B9mCQv6P33fM3Pcc+IM/VaWkxlRVcdlf1UgHmwIpOzLW
Dhzq54ayjgPfVFTKIXKRN4G4shumG+1xZUXDShwsC2LFaJ6avwsYA590muqjfO5j9vjc7EKeVll8
pnGgE8TyXslKtTicEROHwVuGDVkfmzsGXt2OCoHPRw+a9C78iuGpf+PkHdhmfX5c6SUhhPgRdP7W
FwV/Txa2ZJRQLL0f7bVljxwfpShMhKqoAOev5VFB/XIuwqpWkpyWMPhY0MHSfkwLoRIyQ1gqenDy
LYcjKZRm5TugKJP5A1DFcpykA6dyBzN00yYphyyCqz3+yi10o+b61Jy43uvEUFV3PkUlo+In3GCy
gJacqPpa7Y/pNLY7l3iQUeo9LpqcooRMIvTjtbeu5XuEQbm+zuNGR/lrXBRCI9HYMJBQE5ZP0dKm
Eb4fEGUDjergeLt2evCAnFuOH+/eJRfhfX/cL22218MFAZPj9FcdJMCc09uq2jcLHwyFPtgpWiMr
cAYnE/CmykR2OwEiwQGG7nBcIx37pEP18mK5njBLdHqkDlhvTkHUhonPbHj9S7q4yxEFIIDtnzSd
QOtLioQ1FIff9hUz/diCBwKrqQYvI4KBT8CTnl07n3BCYIW0LiTIcqNTy5D2ZxPCv5NvI14xFcNf
5Kn/85dqeUufvSnesGOi8Hv4GbWWG/XFZsE+AI8zpW8l5tDzvy5DxLdQOrrsI0ozEIZRP46EMykr
ZMvFQvR5XZm8oqgo51a0EkZFl9ZDHXW7bzFwwcLZyiVhBMk9c5ET+E0Vv2GCubFB2kKjSwsMk9Gs
j/AifHq+i8KsWLDcebTyz5E+1u40Tc9akvEJMvN0nfr0kzpAl9HVw/4j8YXrwuzIVGWs6+vcLs2+
7HAof8yf3PT9Zwx/vThoYzKXhFRKCUfWlbFLgKa27Med7mNEZ+2JeYzAUaggJIsHvqyY4lrstFFk
SeZT4TmZdkL34qv4wA7ft5BUsFj74hSE23Rm0jBNM1ZG+uWkl9z7U6FCEOwuNl/oxiW1m+Luyb0h
rAct4OZM1g4Zxndyx2pIpX+lj2muiEuZZxXonbp5eOhUnONq2H7f9dcptAWrEeGpOaGVWQ4YnhY9
vdG7KcwFRFTKCPO/54Opo6WX3oTZkR8H8nr28Pa6ZAUgXER7O1ATVB8F9ABLMOLR5UtEdlHqeD9o
C1xG6RLz8Qiff5geVadtswmj9+hsb2FmBm9J2YGtSo15NDw7RbrHJo1n7Si2CGXYMGan4ox6Dc4E
72KueqtvqB9zAnzlcTtQ8Pbxz9BorHrP/lew8lpzgSLDWtR/P5Q5JxK0pHS2HHVv9KdpiwhpZCTQ
Mb11rOBc7tbOkL9VE2DF+yBN3s4FVvxhWBH4D1pxWc97lrW2Rt/DIWwtWeHfKnhZK/jvvRqhtVLR
7KCahu9PQfQ69aTOjN2B8uqibHHxkyic7X+mjZEpDGFBbd/p78SLlJZUBKsNzpos5lMW/moFVr0e
A/T/9XO+4/i/xNtZ67mF6LbBV0hJ87u2RuWZbxVeiLRTbg7rJQc8nYDiCs8RHWQGOIvLirNf5FyX
1AIwrpf3mxGCQ+HEIlPQJK1EjlI5aO4vv6QC6XDkoUlcbK0MYRgH9biUKWw57Omb+Xef2ZA8Mdkf
OaD8QsFspy5+maRV8bLrViTsREuuLXlWSZLuDwrsZHOBGaoZ9iCdfloAy5UFLBYZYeSYFxmwTHIR
5HAwelWGuaGXWQKKUwTjRmGUGJDMhLVxauulPaAD/0PIZCeEvLifez4/iOSGjnYsDrKggSlv8IgJ
BJljJg08CrBmIWjoDQARo8LVfh11Mqmny2O8lKh0RlvQYLcnGdMUvXoos2HMWI4+ujgfPuqlROtj
eAf/koMPs30LHRnkYBBtA/35E0mV/e5F964xNWWmFfBfGgkqH7jkmJl4fo3NEV/u9r7q9e/MG6+q
KNw6Zd2YXck/0uiZ9j/oN39fWT2v3tBjy31pk/eIFvxbcVQ9IzlhFYWSXWKgy8zo/SxexTBGA2CX
3+x55tGfyB7HLRg4MJZMUQI3oVt6IdvT55VaFF7KSJ8o1rWWIJ95Tv0Jqv9bjC+LQXKplLjrleB3
rlf9AvUos490jnz5XmUfhpLMi1DFsjPPZ8dBLKkBP6HSrlD+TT1DmjVDI0pPYzRSilSbeOh3UAAo
5LruGVuJB96SILw+ZUs8GmXKkA68DCd4DQu0CDrzBF+8AEuZ15ySCTKn854Ep4YJ2tXYb4dCwv1c
BQDIjtftaxUwT4BKF/NONUTtPOeE9/oLJ5kc0vWLDd7nWZfhUYhCMBbuIH1aZV7OTmCI0dk5zjag
eMTpHmmmX4pWAb20GGU4+0Vz2PCgxW3jmngj0qkJ+hT7aWslRTURLf2L3cXLT7hVTi6QicmEz6hT
IcZH2q88Oj76tSp0eG+whQPuU3FXTDZfpVMrfewjsKQgZJS3MTDEH2sfOnlLZLLFfD1N4/p3Jski
9UonxvGO0KLlF6tq7JatFzizJfAluFGkz0dyiD8E8DieJIBSFxJ/gV3N3UA6SDSLZ9R/5KIkP7fM
+Nf6744Ksgxzf8TqlJOetMtDAmOuPIKRHdFzj1GIxAxnHJ57Xl0bV5EBSq5/ARp6rWuWMCPTjoYa
A7vLcWPf3vI0MLn1mtfR6jLyEO+4/ujWqcj7SJ3v5fuvckgqBCrqtE79/+GkXTLLYf2vZ83Jddr/
NFC/EPLsgl9aAYGp6bifkPKWXTHf5NHlZBHt3d9gJgS6ANi9DutTQttzEjWtZphUrKJg1O/mSShh
xnsQ/d7CFFoq5tmtYR11PMqZG3iUnX/qMBQhmZMRfvY6GlriAMzF2mGlTeqWLaz4Gp7dNwmii698
63PQ8sVv9RcyIdlhawZEY9fxIr4zXp+RTb7LQRDDu5dEyNQMeLs34dqtyKz6mTYpLBTjp0WQ7gjj
MgtgDIInmrEhxw0GY8DYOBBjBCvZQO/OrPU06uNcKq7ddsg5g2NkR6/szTBzCC2eHS9KGoXzui63
W4dnucYOeWPJMOthL+5QLVAgDF1WPK6JtNY//mQfT0XBfELGeh4GvP9ek9qsT9B0UQD782D2H6mp
3ADjkMmdqP2PDKk1DfFTl4cGsTTqDFYxtZWlsTvlHhYh3iondFe5J13itjUbBRqiNLTtDuyMXgO3
pGqNrQJuEAuIeRxPe37aPy5P5gSjxRCvjyEc8QxGjIVcr/lE9R/p2NvYKeF2kUP6hlmw2SgJXrbq
vIhucc7svaCrCbegO48rTNPYgyrhBLC1HSRfyVwMjVtfRAahOaMPvVTVIEUh7PZMkgVxqnYANuAx
0hq2PYwpdZB46ROsigcus4oZe8vjn1/8v0M7Ha+TddVGCHonTZdGFPStcRb6ntCVHVsrJFcmbKpL
cirCkZ7Xq2sqVC3ctkALZsflA9HZjfgY6rFIjEgK9ISign71Q4+AVz/1+IUqE2ks2PRN362/Napq
Ic1axdZZ8eeX+DGkq2uuFkf0yx/FktrSdaTcke7irJE3vQUa9MYdOHTnOp3xgyw3yeq8/oKtlHZx
HkEgKnwhiz5Y7YoThzOFWF7s8ae3RGznxxQm94/zhQvOx9/F3MXFaqNwE/f3xZ5HYY8KiUsX9nbs
EdsYIBqCW1U6Ej6PBL7nij3oQPCSEluTapN1ATv7TROdFRDaqzOdqJQzrLPcSOtdfuFHBo2lCgXc
rjEbvvSdOYc3q5NLmHr/N80bWfiE2De4Y1aBVa/FwZupE8jRdM7wbpTBWVMur2sCtekFLqVYJdiB
2euEh+sPslFBmf0oL51S2BxFBtAF+B6LSKPLmMFUuYeP9c/0xGg7v0Aei8XZSKHO12cQlC9u5jQN
Ex2LLBfLY+pLGA0h+L6ZHfSm502Su4O41gWqnV2FH9J7IqNVj2U/R8iBJrzhAuK9Kb5sfAr/YVmF
QjWDMAw7PbIYWWG2OQQgDEfIpOZ3YE3GypiZZ8GDkgbIGNTM8ClK2mdwba1Ej9hquvgXJpEpwrCP
RwaDvcvLQZUcw3rmyGGwdI7qICbFQHoRsHKOcW92nbPpKd/Tx6U4pj+nqJ19LmYLJyY88cQKhrIC
Xh7viLFSVyYsbQAqPAZu2wRVK7O/X/sHhTV1EZYgTqOWNZx5prrNxXieO60fM0ris5C0cpDRq5cv
WgXX2uFOuhpVofVKCR08j/GuuZ5hNWcugHNbXN8V5QIok3KdoMZGhaOJMf+WyCr4eFCP6gXrGyGe
s8heqO9S41T+Zm2zq/mvu9qhCLxaYC7NOmiQfaVgEGlpXlksLKeWA77cXlo/qvftVdyzdp5yczbe
qjesmUNzJyiV8jVq6TeM/j9U4uurE9KVQf9+RBZDAEtMBiq3zO7q6445Jx0PvzzcIJl72g5myZLC
oPLIEcCpERT72LOthjYfPSDhhHENTZKVH0p1PiCUWPmKeayobKWHkCnv+XibT1cFeablpSjwxdRY
2rvV1YbstcuoF6cvK41mOQ4bcZk21jBU0XXbJFQoVvd52drc8qBFawsN8DKlp5E+p+uiCULPM0u3
GWojZKCuqSlkU61luerv6sKjGVRjYtfTWCbTy4SSpMVk7c6oU97vbp41BI3oZ+p3qeWgQr5kuXl8
D9SQHDtPtRr8gcBZ5qmIxnL93qasHz6AItt3GQxW3q66RLgl7yRGxFLWZZKgH2pzABjYoAMIz3im
dnuN2Rb6x7sP722x4TbZNws+NOpyQqaskP8XP7x1Z/qcjCfznxgo+yp00y+oXGAS89th8n2OFgos
fgf1+a4E369Fr0JNXW1PMbh47QvHDpK3FQFcAqDRT3tB5AceM1FiNZvpg4ltuacjqLArBuxF0w8J
owyA5pKBBX/6w8jTEABIfmAPRjfcgyyphldqTM5HMinAXTs8HNBS6xHpHjnKWhpdvhW8WyAzy8Ld
LQ+XyAGPSv/9wFzAHmnGulrwkuQFZ397NQEMqeMH3ipnNgn8PEpj0IRRdlOmtfa5s7QMkt6c+7Px
kkuwzvqaSarIBKrsD1k3kdz2SHr1UqMWjy899bfhaTMsaUcPIBxFv/kaKiLHt6kDnHL5XEwVAzWc
iuuldALdKx3UPb1aZAsN86naNQC4uCTkeo0szLQRjWlqJD6IuefEOHvX5OKaPU7ZLam+6hbJzflO
QJFfb62odSGBKp2QAU2OHh8/hhJxFrSaXjbhFzrPSkWDw+MVzftsWFxraMG+9ZRtWHh37k07mAQ8
BO00fnlDUwYaRCQfzgu+CFwQZaNbNwRlro0q/ZMlqMjEnL5imAj9Dz9+6wgeTP7XHfBs42IRypdB
dN0I2T/iMHji1al0qhmKtRUuzt8iI34QJ6z2A2nxu9gIqF9eydEQ8nRCuTMD7JL+lY0Pmz7vKru5
Sv85ZuF46W+y4Vql6ZAsgRj21i3Hf2w3AHlyAqUKCBQ2an61G71Qk8RPsNWMNDeZDJOSTBfZ4PzP
N2dpsTlcZHT2bnNW+RIa6736rrtgLEJBlcsjYjZVoRFN/e10DEItbHx4DfPmbqPDgsOyQ/nVer7C
SI4Rf8eNgGKxMN5zSOu81jeybqN8+0cJ4c5RGgKaUz36rxxU8FCJfYYN7nJnjT0epYzR+E/sgtoe
kHVgx07rFgIL943Pnxzgkji7MFlSPOGrjLTLAgT2IN+QXSBxcMDhCLB2B2znjeI+fFupS1YKkW1k
hgpPgXOTKtdkYq+eyuN03RtBDGxNdcdmwnNuL0FO7N5yt9CsbUizJ+5HjPGL9JCfEoDmU5DGOFhq
pTCR7MEG4X6r/13CvqBDg8EK8vlvLITi6eZQL+tSYNK0TkREXatqRKDfhUxU0VAlByjCaUQ2HVGi
GbZJ3ls3GIJdRNdCqYxAWOs+lfl1+JvGAKlWWlUB88fIoBz85YX1/hEA9k1asNBMuLWncGiqH4el
cAaLTfHCT5vO6U9JY+tU83YnJCIckL6mUyzjyRaRV/XqkbP0IoDVNAiEaWjMocBvALlxoIm2j00X
cBiG6Q21VjzIizl64z39juTJ0SvkKCT+JHjcFjKduv5zYEHOW+xOMnBKHbXrNF8Dfpqjzi53+PPL
Q0zKHVMZO2tu7Lr8huAAqQKYOjWsCImLAdH5T3GyPON/8fwkzEiaJMKNkDDj/NlBjTQZ+THZ0k3Z
4GXaFCASDbqkRzYbPS/2VauXVdgBSCX7QdjDQp5mA89q0c4NtoRyfc6WqcQd77iMxZzNzK+3l0lj
5HWicqZotg6tbfPdIRUah0dGPnUWBHihJO+q075OwXMQpg83bD4eG//9mbcMbuzrkrLOnohGXxd5
O+9f0KJg7UC1h20skm1aFVRstoENhmS69MpCxjxy915f0kXHfovONaqcsmk9g2oZGXwPw04dg+zk
s4/+fId7k0RDq9WqkCaXdJpGGiTwX7X4zo5ADuZ/ouABTwBDhSMPojRQYYVYHhtYGL3y7je0xJF0
Rlm9g4JC4xZTi9ZYFNvmo26aWmn56Np4Q/mfFZGttnJFQCXjrUuz1PN4V5X4jF2SoagjF3ZDzvgR
J9kslBMxkU15sp87gVlgEkgbuoOgJwgJT5qUYqrvhzhrc/jAkyOqOdAxuQUtxbe5vpRZFHw0dzPC
PG+kB8FBB/SdKYaZu6YrbPf6StORSKGQB9l3ZAT8OkyMpT8091RiT/rWjc7SmwPH777HzEgYvYJO
kBUJuzqdHzbBp6XpY+VWf+bsIFkzUKeEwecOPKWfIuIEwtXg8w4KnsH01OZtb1PjV6oS2NKoBbhQ
/K3jojUWuZfctLRvHL99exV0JkNdJOHmM3AiyNsUmB7wZEoHJAUPmjEYhr4PqxxzLKA9iDpeZ6n3
rxSzqM7bCqJ5Sd53hPyrk3kyW9Nh4G4ONlXJbHbIoOUnJjPrBEJVu9VOHSwv1pULzqMn8V/TTCCl
w1oDJ6Soh1GAV0gyIqxkGElZrxLTvlVTPuDOp7gP/CthJOraCJo9L2Sl/uRsb9ZgE1MGWqH/eY5O
Czu4kAM60FWN1b9NtQqP1UfgSub8bFQgSxX9zSFYGWTvjwHGzjGeLPH6CpI0JnmIY9FHkI/0JOhM
4mp7e4/6rDdZUTtqGcOHjbP0ubDp24l9ZYJaBNUDHFCLXocUaBsPUOB9RLhbCL3+hUF+dWu2Q4hc
HlcGfkSLMWtW0eOy6r4wa9Yrq1VSVW+NMWqaj7zYyiVXRbigkn8H1D+eNKFoxCNQhu9aAvfotrhm
V4YmBcdLlFuHJ9yH7kksX3LMl7SHY4WR2Ee5LvT4loOzQFEgTynLB9UZR+qJJh76yfuEqHWcEnvc
bOTvG8YOZn6waIeJEACLKq2BFopCqHrnWikPzgIJK0uW3B3pXkiObndoGd+wO8wEXHX+IMtz4jO6
JPIml6qfSampLlTKU514bewSZgYy2lD04UKThBl89vG0Llb2l19Ogwi6nJucK7nddOQs3vVDJb+c
HxZUWCIYOTmB3lnJ8WhxzneU3StepgXnZsPcRDTRdtm8xUj2gppNfexfWbSUGDRv49QyKDQlQKKP
2oUYFJXFKxv/y1TgB31tqR8f7PWSyVlv74OuEcUop78ZMK7rRn1S9hbwQSm6xlCYskgksza6Dk5Q
dSw3TMebHPtIipx4wYGRC0ojaKMtvGP6P8B9xGnjF4IyInsO8aVVKXFSQe0+OzP/Rl9PZhtKS5XK
6GdT721K7pI8TH39JzRaIqisYTHdBB02/rkZxULSID+Ylf7WaTAEccLBNzX5W4jnH7JY0KA/0Flm
OY/MpzWt8x6sWEMpDJJRxzLKjkJLwXTFW3I8dcwpwsz0FluPa6xWJUF2ybUqeuMMoPi8KeGEdbvB
acsYDFms238SPtXCbgV7BokawPsaVNR4W/O6TjfhXdqc3xQDsLwKbSz1UyNK/DiFMiNr/njyMR7B
TFQv5Bkrc7qYGgE20LoGe1iWmDff6U+aRmIdS4iJNE0ftVnZ62Vo63YNorrb0FudcS6uxEZQi700
10ddGhjp4Jr4vOwLNJyT0gLc9jEof7JBPEFcYQfiZyYLZrMXtSbGcE/Ck1g9H0/hjUGjrPekwkZH
2WlwAtBjnMUwOJIGKf1JqkEoCuYntqLd/yfP9gF5mptjEoulSshS4j6jTkN7U5rwqfpbftOWywJb
MTZPkaJT3NVW8VOok3ilcuO3xktCWRAvp2p35Fd+hmBQJC2y8h0jEPUj0PfVYcj4gL4EO3OVM6pw
ygPuwseU8DsM+EQhQ8gP/8KiZ+0iuQIjR/2xRd0p8rl3U+vV7GegY12KsKBooI20EsZaEQih4rQT
GgYr/ETXZbj+ffahVpoJZaysCQh5uTvsrOe+yNKmgGAvqq8sJ0MpNQKpge+jV3ylOmqryq0TTjgx
mT1xsg60dk0mUdVIpqbAY0Z/ZYFCCUpA8sf9xYRXMrXX5q7DlTSofdvw+q8/scjTLHWFk5vPBRo/
5zkUdAObt1QCHeXSXuVhnmDXMv0X5q/OkQkD7WiVm1I9kdyJrG7JNt+5+tM0RK1NWkTCsS/C6quX
3Ls2z5lFuDH5GhJCvxvLekGDHv3S6bV92SzRYZwiDdGbTzdecdqKzi9SdQ45OqJlD6ES/bOf/GUB
hrFIpPXBAjHOm45tDK/2jqsy4ojDqZ36QgBS91IcWkQDUTLTggGnkeX6owTQPuK6QgJvdvC2WLPn
oE78iiKY9lfEYd3QHfqLFjKguqmaf7KrpKT1p9uyZOiYv/BgIMZ8F5oCBdpzvRgTVKgqg0JmTMgr
zgL1T/WRAzLr04o5k4TNWTzupr1eFN1TBCinJA3hVm13mjaA7QnztmdwT37MgRHjFaukdELsyeUn
CLxR4xG1bJoDM0ZUxRu9UJ5fThauGvVUofnnkRC/9K8BA/QZjuPsdPl9f4/7KE0r+31AnHWdoz5M
Bf8whBWKJiDy0m703HJLX5OK9fUl3vL2diFkMnXnD84eq5TKp4XHyTbtslW/09ktnDSOJ/rT0voJ
VbWof2WrDUWJ6eRznqbP0iOXfQoDFhPQPiMDyNA6K3TjR29UDlw4YVc3gBo3TqX0rOazu4rInfot
/3GHtVP0NDJKEhMtjsKP+Rf3o712mZezRAasoHWZKMRPag6HgvIrOg3/5FSdPoL7NiZlhT7URHVu
JfV1BLyLTBT1e799pMCR/PIYJsW7FPtqJ6vR0ibaOIhVca2p7GNyRqehJK/jxpVCk1jwnxKC70dG
W4DzrUi0VvcoWw5pQ1T/g4ZPA2Lb1G6POF330NztRUp/ZkBYLMyhfPxzftb1ZTfsnDc8DnQjy96m
OXHgEicf2dtR3yyW1xnAOzcIC+JPy+8EOT0AuKZsPaXTpIqMyoGrnTl7b6YpKmyE3g3/w74rOjZq
S84znTVYFPD2W8/Rly6UsUJsvQnLeFYUJ026TerBKuU3zjkeYbUNyni47Cpez8kW/6q+sGDU/64q
JDfSHhw9l557dKyrzh5UxhR+6QgI01SzerD0nh/qB/ssbY5Z9FlIAHvfAYpY2tSWNfxBZ/j20q7i
trkHYWPJy0Yk9pVAjyTZEZ+xIr4T0am8BNigZvuurG30tELcaHsIiTr21xcW4Jkn9ZoqTJsdkcIK
ab9eDJmG/EnUZuDV5P4DLqaHslcNbiACZE5k9tHXj6CcT2y//vL278VmkZ3NSt2aSQPX47ud3LmV
tLjk85c3IDJbEB3VBuPbg46KZ/vF914jZCHZbI1/VQgwn38lTVei4IHTFg4BNoj3yjEqOLR14ifp
vQB++bzJgXUVo4poPAkDW2XBCPGmmteZnq3EokiUWCVZybGwTYcAO2//6ZxXZeRIeMeetKFO2XYa
XoWyIcK6F8qX3CZxUAUF7xEGjolMz/ilDhRFvwrkYl7ZVpZma7zN2ohRJPxa+eNVeTc0NYmYIlnA
mOTe6GlsM5LpMS1kiO8zjis1AFHlMYA2ucObouwnM1Pxn5Ce2mzZJZJxbHj26KvBrFpUgrKEpqXH
4ucilgdoAjOy2M/naIiOyLXQ7t7Lqv/nkI9hQztBeVCvq071pHWffk64u7z79uDlbH3JBdNaUNO7
WVJATzysVtwfnXJZkUJhNzZimBER4jhIeSq9xZ3iA2Em2v3Py94tFnA5LiDDNCx0z7SyZW54ACJz
oMJPMjkURbypODpAd4sBVXJOjM78Kd17e0fTHQwy+blM//43q4Z3XhGMxQ452Yo7Z+BAyvOL9GX6
tNplAjyVVctIkAHawljIV1LKpUkjloBTIQ4/tbvtuCAWiaozcclKChYtuALfkEF2mRviqyA/ivdy
3S+fTeVwmbwYEu9SiT25+dNQmknrEzp5rc8LzomEY5xhfRqKr3xHp3RabFRAFnO4tUC8RwuykZsg
R2Vgz16Qo24gdZDd2Y2t/HlC8sYhiGrXgGUCVkkgeKIOfGm2MJKZuclX90w3v0oYRooVZcrJ8UoJ
3T3SLlM+WzjIG2/aXaRJ4pHZ9VHJmbZYxEvxGK1CCCP6rcGu1RvQMQz6p6TNKQRIDXBhAZZYWp9f
Lth3IPMpFkBAwyxHRG3TLB/MoaergMt80DxyDviMX7kW6ZXcrxUH96J+4AncUu3WD5GAo5H66faU
KhnVcZdqkHigXRkr5itcTVE0LyY6OVuKCkaeqAqgTAAucMG5J0RJKxBVS5Xz2OVZBcXQe7RSOEeX
7D7ar7xM6mrtKB4AN/N0vWyYIrN8611Qo0C7gsnWY7cn6VE79oQwu7gQFcB9bUtaFx6lQJ2kapGP
8osxj3uh90XbeIFKEdLMupVMOdL39vrhyr4aZ22S3z5NCZR1paOdqRaxsSECOzkAKlfk/efM5YWN
ok0zFy6EQWnyFcUFFkqBag8FDTzoeB/XRuVt8t/W4VMJKRt49w6MpGo/4t2QcUaWSbuu2eI7TQnY
/Ns8kH35dm9qKWAzlj5CdHvF1ZAcjLiuKSaUpuRPPoG+gxmzfm6NLfnjTACW88BB5NT16nlyWOuD
QYFg4+kAt8ji73tVdGaqgb0sarHKoJhan7w8GRaOA92xrKlk1X5vOx9Xk9naQNUT8CQsol4S3Dl2
YUNtIxdKRr6GQozkQbbiLWlonHkGmsTbOSKGCNkLt81A9iGWC8xpOepA6Fd3vDhl2S7WqbksXEb0
6+8NDfnq/VtwIknfBfGPjYLYqFLTLo/EEHE7MHkZvh/d9xZiNXGVWr00D0ZVu93ya/lD8GZF0p2d
c0v5NRlFBIXL32rMIXxVMxp8MZye6JXYm5WJy45HoCWG6qC8cIt7NPgJ5oVjCqvz/NzDLGrcYISe
diygz9Fc6T2LH+yJRQcZM7LriHF1D9faZoqLIJhuCirbdUU1822FJEancIi2n/fGjhRyOlP5Ld93
nSHBeey/+MwLMF5fVC5uFSTc/US5lR41vuBpwvqMFsQ+UV23/CD13d8wVWRMChCwria9qbDQIPgZ
qAlDppICeYhfRE4+RCKW64bwML6NZyAz/r/3kM9V1ABsddAutkru2TI23EDBrc3RQ1ENOR7j+/3c
EwCnk9BP8AfrPaMQ60c9NmWZQM8Idc441QuyhJhV96/zcW0Ftt6/83U0GVzunNtFaFv5PM/f8aTx
NBpPw6g4/ajgF+YPBFVIWyhMMnvNfosGhcLdd0tU0sN519/vBkcWE0fKFJ95EGBqWsNiR563L/Yb
0ostHeTC/Bma0G+fJDmwUgH/T4SzAmd+zgG7srybkDjhOMRBL4VUncN2YSFUnLal4pDWttxckhPf
sM6jM22LH1JSW+UnipawJyv/ty22wDh/aOL4W/SXPVfteTqO7E4igkwblKEZufSkC4fidvr17jAd
whmK5if3jW3WXr8+bgF5r8MGNHVUbM6uwBuprnp4gQdubyfbvSp1E033A82QZRxE+sooL2DfSroy
PICEpXAPLF3mDXY7RBFnMGWD9I8YbBuaXPeyVG/nN66LyzsysvZOGoI8RX6MCbOcVr34C2QxBW4C
tkJTInXK6hygrOn4jsVoDkh4g5f8dhkkyDnRu4lHTUjc7Qbvlo7rd8T3MhHid9F22z8bv+VWds/Y
R10Ao6fueZ8TFIC/AJBgq2AhFzsyfUzi9FgVqAYNTKXMyR/3Yt0nIHwpZ1tmU/mzKYOgWCme9aSY
if2HLFhU+bB4S0EjNjD9UFLXVS1gnw1UGt9refSwW5fWwuL2wt2edWmtW0kTNZocvKFF2mf/MTfl
boTfHQHDbtE8bfPTMYA2V5BOQmvt0dLcvZVwjM7Fwq3/GGh6YhCkN8eyTjHhZV7Ex5gwYz1uIWxM
fkx7OljTw7s4OHKIKKZqI47ykhisU1Y8/SYPw/9SVaqTLBFOkqR0QHEXm9iMI7U/hgte8m8GiVq/
X3vK73sU2dz3iPLS98ZdmzgdP/7kpKmrJrJ0x7RCQ+yg0cF4sOgSEmlWw80RMnj5vYldx2jc65La
kYJ/Ql94+T7ZO6WLqnP2PqpObfhTWKdDgQXNPpOmFoRdo6xPh3yokQc7cfaPPaRIEEyz5khAH5Bz
unUJYEVarVktv8TFQWL38VgaxAYJGBi+8Htg2epi5AGji7L9AbgDqGsgdtLCnwW6JI/StO3xz/UH
bZPnD/YHLY6uttlh7t99EufidaFPx14LUO7HObaKoViRAxva239pOelFq0OY2Uwnlez4P+G8D5MC
g1Q31hgO7ajD1oUUaKRKyXNINYXsGVXCnz36+1DBpZNrHaQnRWkewxaVYICBRRfosuBUh3wPsaXo
uL9epK10d7Cso0OLpjGZEyLA0fou6RTJu7/r3dR12L5HALR0CfxQuVrO/os0APW64UtbhMarj5KT
aoRe1NftBFWiBBHSJTJN1sb7E4f0ohmDFbFeJ/XAQL+BTWm2LeDlir0PpgDnR/KAFOBx28lZdxbd
1cOJ8KgPMfaeeLnNAqNEhnH2o2WeNNO+PO+Lk0fcutk123DmKuNdkU8AQGIpTctt3OiW6oRA4QOo
0NYzl81oDbJCDwBoomtu4mMlGx0PbqI6hiMkNDgi1jH+H7afSNlW92WOnHVeJILyydd7tle7KcOp
JF7PHMpHLbWYWcJcY0MJql3Wjc74famSswlTFhHru9ltnW1IF/GCVHz7Cszjdgo1z4YQl3aWapcH
qfxRxTBVRWvjq1vpiXG471V8WL7ZaZx2IMpKGnTTBjgknfm/T6KuemYiWsB4BBG+NBcYibhy9W2O
hkC7fBPM4HkaVXd92mZ4xFZrar8WPGm/0yMRKbKzHNUiqo7dmIJ1C/myMNmNSqvJB+ySkVKQlWB9
tSl7RqJwSg2tZlUhcjX7sbgZgDIoWgJp1encmipGXLBhc3U+QeXWiT8Qq0KH+qcioy5sVdEO7i9K
8zrd4PqyQuI4L//G6vLYKiKlsyQpd0a+bCfu9gEG+F7rsMRMpeA4Dx3Ig3tD+0I+5PYIyCmUjrwV
+Zumc9WN05hTm9GT/7TEQALjjIYUqltI36TAaZEQ1ZabcaytOxfyjSfW3i+EHzJh7qvA3+yUSNNe
Ain+SkYCEsJXzHQQNQSh/gi67qJqytfv7DOnN5AW7HOoRJ1zeOeBOtornSPh/fgKd/eAkzeJBxvz
4z8B3l3nPCQeCRTnkZFumfoHCQQyEb+Hk0vjjbf2dhNHmHGYXtO4PiDf/BK+RCxq43GSs6e1iMpb
8pBLr5XxzBZataqOI4Md9kCSn+wHmfqTQMb7CU7JWgAyPAUw126TvvYEQtV36tBJfLlR1zGgx3Mh
Cnjl72AhINWkVG4fUnZSw4Ly0ZhFBbF08/HFSwEU9qq7X7NLzdz0axV04EUj3vcWDYncMHdrTk1h
nBj+mj+Nqk86fRAoO9X1cRmCAidrVr0MMaL6UMiiO//yexEfKn+IzmkHcGo36mwUl14TnVL9G5jf
d0grglXHLZlxvxTLEvS79zRaHOMPDehknKSD/fH2kxuR3jGpYb6iH0oFxXeQ9pY2kkF+ufeKDCOO
BBBWSrRkruoFn6dHGYMGsxupJAKKt71J/78c01fiLQ/GP+3OpbU873/q5eXAVBYtVly4h+XaU/z5
rEf5ZoNPm8PwlJzn8E6i7xl5bDBND6h7i320N+wDGXJeIEbai4toCtf6sWbAKYrGL4v+gNs9ksq5
ZjYlQMC7g0EVa7aS3Bqhbmg1j8WtKjDOFKQKbtBmdA54NZBFRqn+htcrpYehoCTJy1hmwQofU5oc
Efu5e7cQgkCfY0p6ERUlLgEK1NkXEMdoJIzTWHEaiqvJhbIBTm1w/Dd01qwOPuSdy1u8hhNfGwzA
DkDjzvQSuui4XEEYxWD21nVVQCr/KdAJCkfnJu2HlSzcL3YkHSZ5KTq8qH+eeQP+dokDEqENWO2/
Y/VYqKdZOUX0/lbXNZDetMLzCJTnJBg3Z9ka9+xcPyCvXstwvbKG1Nccl6x9BARjL0/lIH/5SP0X
ffxhEIHa3jJHMQUBoYoVhXZWEKu6KMh5DJYZx7LsR7N/0VWKH83AXrh5Z9ohGIbSCqaId+9WeFfX
HoQbFM0qc1kXelU6gJrFIvT/cDTIzr+t68xDHeiCx088TKL9emFpgN1w7cnmcX1MYXShVl+ryv68
OxXGjBbFdQDDZKvY5AJJY7YVG4BFmJshoS/O3trvoYNlHpEqs8qLp4khPv4U/kSv+Kl9q/JEKtO9
pphlSelrNyKCWXlTrHm9q/msadF/+bZ+8n2TS5LkROTWj71aIsV/VjKcuFP/eHXYMuCCQmzVsV0U
zseriBGkivuxQ7XcYWNFAaf5xES38188BI5cNHuItrMLwErKlQ4JaPRUBSdhJTbiLcAXnGXKjZD7
JgbJqAMBAwWOMcGvNgieT6EuT+a4eLOavIISnTPpAiDkNZrSn7OW42l3EmmBBeGSEHh8R3xaxlZz
hH9dhdlzK1lEQQJtZ2kvv2FWJ9XZAgTz0/zICp+F9rgNX3Pk3ftHwPlvhp2VEj0MqhskRpBvHNnr
UxPvWQz9POfrbabn3sHJT+XZagwpPc1j2OWHrl6x82RixuSZLhtLI6ZqaKxoDG1MFZ9uOFSN7BIo
VbLHDKnXoxB/YgY2bUrX+m18o5k+J4owzNC0kusfyivVy/Wc/VsR2L8ot7W4Whz2jqeL+A6r0+Z8
BGjemfsVOKoUyiHSv9124g9SGCdxK/0wWXyFLdAqZgWZPk3KPGSVfRZ9OdRCCqZslY0i6C6MJPCB
XKdH0a8ZYvPY8XzojWr0xFfhdoXlMpLHiEVRoqDc0s/hgP7nMDneEJC8Mhk8MdvCDqlA+SaKPF7y
Rowj0H7q4oh2TRCB9KAerXJH1YAeXz/B0+sjqZCTJLUrgzxB7AKUVRQt29Hz3zuD+DFnPTIkaHnk
1MbpFHsGVDjf8YgeTHg95RdrydPtomdSDJ5+jVluu28jB2qNcSBYKokPQ9wlPaSMXklpgMqr8K+X
M4877t20Y1SLdWPZ2K70gynJBDcv03FQvm8Y/JzhoJfxNsdtEzSP7BOjhhwqMA6xDyBJrQVG8pGH
5zx5I4SqgsaqSP7HplpPUjz/HPqQCMRQXGn6ItPL48OP6fTg0ETy846I91vl7oOg20le57aWkVwr
wx2Viw9JfEBW9EhTgTMTR17Jgd6evlmxe5Svfzm0z3v8oOJUptvRhyRsAG4Qk7aiUOPU9FsiM6MW
0RAms5ZdaCua/clQGVT2nC3za4lQUpOawrVmrOtYDp/Z2k1vUWvs9JzQuVfGzahK32QO7tW5yzmb
7aCu4K0Qumyo2kiykgpuFrrqI8wisKhvAR+5utof8A4dQFVandfFoIrmWGvubvPChlOE21IFrwfq
5BY5xS/+6ZSmogzVrEy/H+bxgbCf95WZJG6vSf5ZwAG35+2ZLUa1v0Qi8H6fJpThH+daoiDex/T4
DCHS49t+9RII5Or2xAdJvHEjMAH4TEeyv9U/2Oai7iyzwgHBwnAUrWtnOCRk4bARDjLqHJY/vFaS
5gKnS0LADq1ywaA7Kxe3D82XO4MvxICGJ+w+3t3Ttjmc3kmexP9Exo1SFtzZ70jMLUS/35aBso0g
Fvaw/klPBTYUjskFQgpZpEyfGPFLcqTrD+ENc6rvh8AThHrCSkRPEFr8KUdM2zg62K4pQbGNBM+T
7WYHfGOwoIjVGiLvcoknloZnZRHSql21o3h8M2gAsLGF/NAS9kH7qgxynpHFbGvcNZV24bhB4Y16
ug1i+TnVH8hIOM81ADgIOjd04/tzOrk5N5uCgVykzwkSrMd2JFk8qgAruZXjVwLUd8HrwcVo9Vwt
cdkkTiTHJebaBXwJrr9gELPiXu17UEfde68LytPn6GjpydQlJzZmRGb+GNFqt6kFsy+15MChlYZv
oAq+akJheWVyEr2Ishbzchk1v/O3wGI5KjP9AcV2w3TVFnsoe4kF5FP2DcnAjBkIEqOUDERBgbiK
SXUzQFwmXdLCG95bQH5WEhKg+ifkx+lvUMd3B5dzAEJ1Cn7WC/ZTFsOclsR99839OwyaAGSj/Uij
8gjjc4gHV7X0HKG6I/tw3dbHj2Orz1d8YOoEeXjXI4fu3bShtzJppy5IUNeFfI/QA+yic3b5EijE
+qFRZatzmDV35TA+MMif+NW8ybhIe3Hkethb7ayH9heJATGnAL8HKTuMy1M50srQlmyKKzfhevpD
89eaq2yaPNEBy0HM6F9sCeJPG2aq2/AryAbW/LTBxrnQjnJXq2zQqxYVLXvyF8LbplEcyewmE8la
J6MblwOe7/1MApIdHLCdQx0bC/9ERPeyHaCWvsc0DDTfFeYABQRD3yYgJ1T6ifAMXu22kfe62Rbl
X32tj1UI9zWdInvP44C9tcVVxakUIuTc+mwQ+YAwnAdGJe7bWClTYkEbrPHz3wuJG4+40U6vZKPW
AKmwWsrrtIyMUO0mXnF6c6v4XdYy9GgUmSdDowO+HoidsvKMsyoGcIP3Hw5d4DPBn8oafi6Hohzn
nZL4CzXo4FObmUYOUomg/TR5K6G3yqHkRlbjSUokbVlct4/J5ewQb7zewiVTAd4wJ1+cWF/lHcEl
3rDRSF8bFaQoM7vJtwXSsR1a8SjlwPibUlNBdzibJPWFoAyhCQk03mEsK2//fyvxwUuZdKFc7ZlC
2m1CL/t8HVBe9buUBNFudqlW9LeeOUwiKnEX9cJM+6YWU8M63Pukot+ONQo3DHdP6PX7KwL50R22
S2pskr8lFGv4l3sK4mxhzajI6UGJksSPziiHULWzDeaH7ioiXgu7YJu9RbbVJtElxB27BOJNJoal
ZaaDaGGL/FCRHRkG8qHxRDCxbm4OnLSQBtBU497RJ09XMDlkzn94GPR/zAL0KezUxi1KifrOPRtm
bbiaYz0yrx/eng66Zdq87igSXtzWMn62PjKQpoEN+Yg11BGzYjOEx7envhDBW7yOhTLu3DglCt0Z
fb5AkeLZp3daj+5hwq6VZrL9qrm57ty1Ok1nl1vf56SRo1y24aw6uB44mY5GjGA023k23zQgl+/B
O/N+FdmkGd+g7EEVt2v5mE7Pr2vTE9hy1/bKakxmk198/hfLJJ9avnP2dJL3WjEYq8B6m4idkgXO
Hm5ji93EZl4FL8cfjEhqHhAB/mqAuAqEZv33X6aGj4eXzAgxfjdT/Dpr1MDuJq0k+lW9RJrgW63g
DtLC4QunhW/W7Tx/RZesbjMfINtTGLvglomGDF2bcVJ+Lf2VR4WU3rTf1nr+kLfFDcd4quOzl53T
pOYiSA4RVibJ0iuslHOUpFyZGYk1h/WcF/xqmLW0MrxUGC0QlFtsnAJM+tHDuEvN9twFbdjG53Nv
qabTOGJkEsEMvStyawQ2Y5H7ya+uc0WU5ye1uko2PtWXu+OVmk9Z+0bSbeRQSNvDGM5GtcVuon7R
ShmramR4Ych3uAn6+z373YgUND37jt7CnmdOwVDOIdGopu4JzjhMJpJxILf5+wNrjMN788jZEACX
Qc/bzkuFAAWSCLYJbqbtJSn0tDIA+6OWhFRZ0K3y8ST4DiPhjthxnDzX+/5Fw1bsbg72PlnThBtT
Qo6nzJsAhjhq0E9S5dsx0ewKyXOWffLU/Vje4xDrmg6H9b2rw/pOELbnzKhsGqmDbBcCD8iqKBY8
8CrCLcIpTiDUledLAuo5VOOxRgrLqqzAANA+otXjW6Tm4NPvPuIEYrcEpl0H9scN5YfZ1xRAlr67
D+Qt2ecl++OxVL93zhrm4b9RI6HO9iHE6MoTF8o4wCf/LVpnll0wdtPTNQeE9pxKG6WNV24oy31d
pCPWJNo9dsl/03GiGs+13dfzp5VWK1quv9hZQ18xi0bw23PTbqFi9ebivQrg3KP1c3fHvz4wxxSo
1YvxhzzYDKiR9RZg0Y6MDTDUaLs8OK4Ys0OOZbzB7HGtMkoj1/GHiH5qDS5LAyX5VlvxtjpMVaeV
qonX89QYuOYj0H0FlU6sgq1mdRUdE1gPPnFZsLGRIY2daDrxeXQWfNVst1TUFFYACGp4YDvmyGAm
T+DmAaU+DxatLnF+aEXNXXx1zEZ7CxI+TPQnMWcR/18K3aHiYWzIbMn2qNlsVkqesxUGz6oMd9zh
PnCBSKs1buO6HlzwNbOloPHK0lqkXs32JQS+xMxaOoFkBmXtb5QJaoHcmePMxvhj+niXSQertron
DvinCms3Je71QZiMmjrpoqdMVH3kCOUvtmVhIfP1WkdUV2PEFReBz8+FwFPopVNAet4gWby1NvO1
LnJPct5iK2FrPXV0Ymhc2JQyhpJn9HDd5GmtPANgD+fBNL8yoLKWLqLVWJ9UKMINAR7QB3DaZqv0
TTDvLFDUrZ1xjVvHSx/0LgSzHcoBlmT5jL73dfkXwXjYyIhDVdLbSGwzoq1JV7EFdGTgUHW1qXWL
pdR5ciW0czbnJrIlL2gRihUG9fFgmQnjg3nIl9gQmsw6n2UjYaffsyw29e1exQlVzLQS9gTOcT5Q
KLkwGBmohlB6oWGBbUUtsEpwTt30KHyF1KIFlEOfmFdc7ODN4qL6S0iLsMvi5lglNaXr6qpOCaFq
WPxyyQCGgH/i0yCzPJ6r3896drc8qsyy3wJwv9zS783uTqDlX184Cira/jT0pb+Axao9rTAb5ZtT
UCWcUv8GJed2pIb0OTPdhvFnw3dNdj+7DuvyhHNrV7q2+us4a2E0TmkeBe8vVjfOU0iwvdvX0LqU
CgIc0WFV1woHywG78aebyojkX8Xjg7HRqKLoAzZBv+WgLEd6wOMiQ+48ZpBs4u/+xq5/K3ruPCXv
aTspfqqlxaDUKsLTDUPUSA0aS+KWaRobbrKdi2Mw8QJYxgt7x+JbbvSxKUmJnxxUUecTpfOq0sAP
8b5lKelEvPN8xqMxwIGT1IWUQN/qmMgx2zlAVc7kjcJA07dwrGc/pHqNixOb/wUlkDjWTuX7K9YF
9hHX/xt91vxFoZ2bt8RpeoH6YoTrVSQU+8QbwpEr48of6pYk/gui8aLrOImn7a5SBgN5gat2hVoW
N4Attn/NPD7Dd1G5+Xo1s7/86qAv1V1kWJdKtcDNYWpIHXGj2+CX6ChMJympAFZiZa4pyhcRiZhP
NioRjbv973jfwg0/AZGVJo2uUjMoeF+K0BsIC0XhaB00MQO8TfXbY+NQlhfgPtmsZFZit+pXT+7T
DEYJ63nPG3w8NyYfvj7DXkLrTA+632yB6mOgO9KpU7r+pSawVXpYF3eBscqIXCJB4NBy0IAnyqHv
5Wh0rSYEVNztRSn7E/bLGhDxk/+pQWvt6fWBF8/Bj2lXaSNPbEVyWghmmcMDULnXLkHkZltmr3fB
NF0zri/0UYT8CgLKFF/gS+R4tJRsV9KbLQkIAfE6c+ilQL+KaHkEuFNRMqIURWgdpw2TAwjEIAH1
n+GDSsD/S3Vnzi6zRCaFJvM00eNNwafTJQDiwYiBcxo58W9ENFMHUHuZkVZ8pg4D0F0UpL0I7tdj
Q0lsPO/3NjTU+d5IdhjcYDFUSApsIJap0vIaXsiv9Glg07mgG9vxfIzfU9oos4f7pdg0dUajsteF
jmmNi41pzI7Dkdzw+hWeAMWqxCaFBfNKK9LaitgsMPBCLb4QbJ3MzAhny1YyrbN+LF4mKLxUeiZI
t0C2fbfgKtTR1I1OpcWvbYqhKNV5KoZjPH/8/dGfZJWdPEBJQQdMMpk2GbEIbjzcT5eJGbMXd1Ay
iSbtld0BtehT2sY14/9fvji1hpIs9wqTUPh2rdjIcA6jzdD8J1j7hE2nmpT7Ujik+aUblCAfXpDz
MScUSpl1lNmyFxwwD2jHkc45hd0VwH+ILk0d0CKFg8gBPFC3i/lVqdRvi2w2fLb+QkP+1rLvHiU7
1rKQmIz9UaMa3d70x4uVAKr+ofVsmhVwGLmiia1MKAj86a0yPIzm79w0W5Qgcl6q2VVVhotmBJ3v
fgCyle7lg8foNqoyvDZkokkcFJjAoMMRz8geBRtm89NPlimNW4sAsnH3zFwVXqoPSA+1LVjpd66F
XtrVH+kKd61VClJzbifRRO2chE9nz9y7dVQo2XTjKHXDWdWYDBnqS+RAf2pzflQs0qAB1gNl0ArY
ePUonpEXO6PI7zvU6iBgGa5c7v7p2X45mE9z6w04+nrW5huuOYs8GDkSGVRRTkRIrbRfzL97rLGx
HNl1i9tM+rmpuBaYSGWBkEcWYjsXoXBni84pkZkrID+2eLK8H1+E8qh8yuxzuAWTPDYTkcRL2wpK
Au5lWpntQ08JljkOTC5NkfiLThiGAGCkkl7ZxGY4QesWI9LWxWK2HC8AYx9L8McS2N6awFh6agFv
DNjptQhD8n5saVKb9qjfg31wryi6IlK+X8ouyLxzxkQtgO+2hko8HAIjHlJZ4/I30g7EJHAuEpbk
zSTGlmf0wEJRRQGl6kILhiEXmVfCjsTgEO+EU+jSbnyG48bMZJKw2QKU0TsTCEG7mQFWAaJlI9fs
9u5Xca4732phOpDSOq846JFHpMk5e+C+RHdWY4ltj10Iig0eQnnHdBxbQeNeaVwP/SRUV3w5MUNa
v6lt9NhDdKSMUFYvq+Nat+XIXTHuZqLIIijBRi5Jd4LJqgBC0Rrjbuob60tJEhFjhy+AZ1XRC2AQ
dxp3IoLBQed6PeGwLxTwiyISavZLUUJ0FKYcTOujOZNomGdYipvwnh62bF8fPiteQ665hSxnlTxg
50t92+XhQ6sC5ofm3afMo5Df3mNhrpdXH9XJUJkHIjoPJC9rZGmd4xgcZSyRRbb4Bk2Z7gueJ/gB
AvruPpCF+UZxNmZprCpRTZQtRoxXZxqHCZi8JJhoDKMytQp0FX4oBNFk9f5LvGuMhvf4xxI2Dfzp
/HcvkQfzNY5B2Mtx0t3uBECw8w2vZFt0lVyDfwIHdI9xTWkeViGgj8uBuv0xW+zorN4ZhlxGxLNh
oQNeNwflX2inUEVT0FhR61VJs5fRF0tK6sbLI9w0UYRYKRc9cb/PZfqzN/UO4YLxkD/KnAvS3tWx
hkVDB46SIVWC6ByAuGH1wqBF2sqEtl162sF3phyo6wq5+6RIgCOVCNOTcIC0ruC/S7sdJzFmk6qp
ke8gjvH2NHqeTvb+vS+ndwDl56fg5yFOPiVB9tbJ6X7o0O7TFE1vfQ48sDH4/Ac+reW56SYGPVb6
knFIOKsBiiOX+WXeoYByEC0uIN0RCQ3zp1g60BS7WOJvZDj2BZv4XJKBmiErH5tlwkQqteHsi8dp
7zVjlxJBs9DdjOS+y2SvddENeggeE5WijP+gH0FUtIYHxpQ/R6Zw5JJqgAUYVbqaB+likqBwU3PE
rX7jCQ9CtG+wx2A3Sf4qI2qIALjvZc4Wxu+XJsEDlOB5r+J/AB8/iElMH5Bnh4b3UqpBYyr0aFG/
dizQDewhfPTlWf2UsPFE/KoGdhmQ9AdTb41vTzgLtZm8/YKssy1EW1b/I/GCyzVEdFhTGsBBtSkg
gG2H7o6QzQRLbbAW1tL0E8nHFP0VZwb10hBZ0lMnRT85S2VIoeGjkYQCGwJE5p3wLm7qYFypxqLy
h5/Qd7ktqZRxVvOoy0zUf/PWIdxzk4elaEgChcmRmJh/BPvl+0B5mkZazPkMmhms0plQaOz6FCy7
3thRGwpQpsKFP5zHx9DUbGn3XqCBiu7odZWIbf03w1ngt7zYYsKp5eM6/s78mmTlAU8aGPeoYPR4
LaNvpzTYGM8vSKkGxlT/lPZaebCPmqr8TkFazo6PEM6salrg7Ku7hsqiFPlCc/n8T7jVYW5HUOSV
z9IAgGkYmKf7P5GWJ8FWcCSCYdqsvZ3RkjrZaXp6dRdyrjbwidF2B3+wPeNFlXi20124xcDlssAp
55l0rYKAZtq7816DW7ltB09/b4wOvHgR0kOBpzKP/N7OiHLjJ705GMRPUaHgIh+SojHor6tv70Ee
S2vggyuo/fXbwBMhL/Le5EVRm7kaRAu9kh65c7BJb5R3vhZIAg01aBPYjlWOA9EEk9MLAHdsYxnT
EyXUpyBTDYmNIZEfCcPdW3oWhst0BGMVdVwqG0qBCBiEhuE4mux0bjKgyL8KfGF0DCWwJoFUybiU
JMgzG4kHtakl736cWNF4cxvZkf3yQQfOWJsIijue8df0V08NiTgAjZUHqpvk99pbLG/oIBenLhR9
oPt8VA5KOaZmxSVHrx0IOXOdswkPNSi+fHIYOJRZzPdn4v3JgdSpFEk+b1tmxUhjOpmdcS+3YX9M
r3IHX6SPCyMFNPOnFr9n2RYFL/US/lwxpJfYt6Ek9oscFHOr1YBkN0/FaUovJv6uVVnkB/jKyS+E
D4pZUMq2BiILr8l70t75397M9bic6hURzDaxRfgaDREgWtp4lTIKPvKU4/yRF9DJHQPycu5BaJYC
79FD2z7zW1ndULAtusB9A8wgr2wMUgc9pu+hhap45qjN+dRWAd8nlCkeZmFWNuGB/qa8c39xLmFN
esO2xRbpbG2qP074Egq88FQKc4fsn+wowt3lgu5tMX596LC9AQoU8Vz5veYVYMMJdO/CVQHF2vmE
whh8WngI1AE+8TfTTmVAdoPRspmbhSQLxR+ndrZNI+v3T2eFm2S0FgTcm5hRU3IioCB/jDcNwiOZ
tYARroYiTn89Fn1vFQUoUqZ8eC8xNKyukpSD1u6CgVkPs9peN67+Ry7hEeb7/7P/PBpYEC3d+jBS
vRi0YQ+EmzvY9yHY+HfzfOgFoD/ydLhvn7vrfvKHpVU0Lf/lCRswMPrkSMkiUB/3B5iDAkcWBFKT
rQASwSJqto8CAnqljugstyMbWIlRMAuQlQROvTzS//3ZiH1Gp62gVzFPRXmJK9Gq0w7LsK0Cc7Hw
YJwaA0xXt3lm5w2ARdXfsvHnZ6pyr33jUuOSc/WEfi1NlNYxGAAy1y7T2DCX6ksTL5+btr+ZfGD2
ar2JBRfaJDTDYOiT/8USQDt3maWIGE8mLNR9fZs+Av7Joht5SsSxfW/3AEcTkqTQtCycjZgBC05K
hY3zCBApd6Zfi9Y950OYkz+n3QV5Gd/Hsayvdt8HrMk0XFRPLWJ3mkru6timFGHlHJr8KyHFeohx
0lP7xQzCv8Io39sh39E/tOFPW88fihTBDBT/RZMW6MreVT3pV9wlbNJFMgMAaE0qZAyoYRqz9M9B
o6U1wcFUw/u8zx1AGxAJ2KVRYc3D1Qm7AmTEVxfWAD34gXry4gOglBARrtQBjfTMg9+eiJF4Rk3v
ogX5EmxBqy/0+DAgynkb5EvdN2QOz5S4R680d3niaA+ArMfHz/C1eSSwM9KpYn+sbaxgkWAvJYja
tjhxf4xFGtWQvhWM2pZkn0ejhWMKx+nX+ASAv9UlHmAT4jxTo5XJAgTHuD1am890nKQFSPBu7Hcz
uNdHXjC4U8Q7TI7PfvjCuyJZT0ot+9aAdiOq5jjj1AHJve3X9Utn11C2Lq4IwP/cviThRSRtf1HB
pModr/VYbA2Qj5K0cCcq1AiuEqMHREAjml80svhQZaWcznM3cU6HfK0ohuMUodrJJZcdRdCgnKvZ
rAsWL/1KbUBPxqKk7eIjMJT5qe9yQPXLTdtKWQh9COOTr4y4/E2cwp0kilIde3o+b3GJPddSj27p
nDskqL8qsI85XziQ4uTAc6Yd33AATKtaLFTP3IA0rbxf3wtd8xRJN/zxyhfGYp5O2JEyLKpilN3q
YUw0IlMaMRoihkq9U6weKKxP+6UZbZFkudG9zOMUYpkfpxXwihlJdfV4VJa+H9Z7DZta/oerDYKs
vV7m888EE5WeEjRuW0a+MSLSoDQXtfwddbFxoHwXMgfoRfdAIoc0oSg605vaBd/Fp0ueZyyZDhKG
TOIypw+PirF2GaG6xyAvY5RPxEA0BM5MXDmC7F9A3vEBSFiofi6M0N1uOiwXTer0AhDhmKWEE+vE
26YY89TwGbBokC9La5tKFoBPuZ9iG3iVREWubkAC6/qZ0xqngUUaTc5kBPmDznKKA3GQD9qoIii5
Qn+yofV8CjsoxV0n31hoZBN5WTLcyo7g9t/o/14e5WOL4Nc011NHvTR6yu4L+8YS28vRoSEMhXmP
gB8OFQbY+JBdJ+mSLBRzzmNQexY9QeFqmhwKFhX/tZm95occQ65Tdu0mPUrZMMUfXFuHJoM4VFok
n69oW661js+ZhJvtzSV4mNFqRon1gp9IjYEBMaljxZR1zIl4hWUO6HczAVKmbEO+OWc8ASWVmhZ3
w2ZFPFXANdnYjhdwjWFbRLhppDcmZvLsu4dCFRWxZBnyGvQcZxxY4KuwObnKPi8/oXnQXa8tAS4b
f04XNm7zWbn+iCS2f7FCH6XXAQCj2rWKPXTPFEuKMRDKzTlSQ91jrEZxrgcxKInlqIypfcC85X0x
mo5EOqRtlxYfE3KjPnj01h5TV+Cjfb3lMTrwm8/MBzlvZppK3qhoG6Mo/GZLncNcaX6QkKDa/k52
3czk/pfbtKMhAW3CY+LV6rDh9U7rzjnDWV9k+QhXHKfKCH6ql+wuQWi9hn4oZ39eh/1mVwHz3g9L
bnDdwQ6XJ49XPbq8fjpYQsFSjzG2ee4TO4Cg1c+dBKypiCzrAHYaIVApSb+Anm+/SCHs0JG2qxBz
3uzsR/h3uKCFFcCM650ygNMPQ+8oGyEPGqzvXR9gyMX7Fq4yV9T9G2m4K/GopOFGyCO4Qa8C6G67
YrvzfjkXvtun2wFiHu1yeX7mI+Ju1MfFso28S9mkeqbPsH9ttwsizHzOJT5pQp+yekE9MV13OCv8
FCfi3X880zBonx/V9kOHOn5Dt59/2ewBxgIz3z5cxV09F4l5ltki6lmUxAn0o5vpP17C5+RrCSuh
hpRUyYLi244KKeOR/yJllvwUfeTDYHihzf54wRfeW5qkarnb6Xm04wL2oPKUXlqbuV1VQa82AlNZ
pxRE9Z2dEFSKHEHHZQUnqiVJHErrtXmrEx1b5zAUfpI3xMl2gxxKyrpWrwp8Pet3L4Dox8k80QnH
DXQWjGtEfcXnH9BSMp0m6z/l2R5JQQ1PPnWv96s/qVYkiBgdoVMhMflRHOS1ZFguyH1Z+1XSco6q
QPikgNyuSvF7wkxE1s9VX9IUvaLNsbC5xjBdoEYjQuseE07aSlggKJPN0+KkO90CyQnaUpVIV08r
btlVIL1r2dvm1xfYCZc8qRAefqPJx4HyM0qy+i+s9iSjRF7ucQRwIxGsf5oUyMX3TLupEZ3XePK/
QoF2rkSAYuGdr5KP/ETcWznDfxZnOeDEyPLW4G34TciOd13KAGEM1reQHgK+AzvTSZHg7VBFpZDD
LellMm/hfalZOqkkIGHnl8aS0UOruDApkfuvCug6ghoLhkRgJNxQMpFs0+/Iwb7zW2c8DAKeZygJ
RjPu6zPDK+yI82GcMYh2EHo6etLDnYYwC2J5hIXpPVFuwWlh6qEpSkPTR0AbrBu5O+xf6bJ4cq4m
zszaelaxJE9iAHEWDG0i+FVUO4/ysMYgmpko/cvOKcx1H9VD1b6Z5IVzgDUvMivgNsGkbXPGIAHW
qjV4u4UwcChR3woe+NP8QW6oOs2mp+gA+2aITMxX5vvZwA/oCuVOMs/YB+8LTHW/IEF1dL5E3P9S
biE5PqjZOFNMjF5luLXUNQTJSgMd1x3V+36Gjtvz+ONsJan+adp5zilAoyQof8C6ckGwc4bk7c+c
hX260YDjLV4nXRiJX1nLa7Qr+BHL0ihfuCgv2soTAD4jKrmMop9lda3baFK7yfzr+jkuY/8HY0vo
/RsyDhzrHMfTZ7jWKeO10lkHg8mqCBouaEYTEgBCEj/I0J1LS63gtC5tQkN/Cl4aSNS8H26zDIOg
wD1U8EVurSTodXj4OZg3r1r73qJ7t21K3dx+Zd1jTQfHnzR6WCM0227VYGJ5tGMu+DCsf6Ta3Dkf
K8R6vEc/rgcVc/jcXJgKZMCW0TNoQHXJNyxidifWEnBSnoozPbRojkVkPYlh31rMEnWoSsqT1VqO
LWzF1B7ljc0p4Wv+8c9v0NALGYIWkEIzY2KXkXIh1M67SLKWf41OL6biAerain2IVrQxeOAVmUe/
joOIo8oT3KvTHeGNFauO5U80K5mpm5odrnI4keRm8/GUpnZNEGeU3ETqPYN+l+vvElBqb+21WQmk
84zHrfvSQEG0AxXGYXICb+dMO/Y0Rq7ACtsm1V3hDC0gfOrbi14yh7za2LpM+1tLJYb8eVTcjpa8
1VctPPSo/+fA9eNmzmzP6vxFt6oY+UWmeA3nkcRsW39oIl5Z/TYFzIXKmP/+CN43VQWh44tLt6z6
7+RNubwG1Y0f1yoYy7GNTHFS66SAmwWZ5IBkvs0wrKJp7Fww14yIHyVhc8mglERtC/bQv3fg81vR
BMs1Rr6BCX1Ec9NSyZnnNVQbtnSZ+OZvnTNqWpfGkTQjgS1lm4fGIJ1SnPcmWNzaEd7RWoolqdYW
Qca0gmvopeYDyCRplYUJ/1X01J8z9E0tEy4nnhMaxjH45FX0YNxy3W6qDv/OCIH0MPNDaBbTboJ8
OBRvFtAnO4MhRQ8hb1Tvc+EXtq2LOlz0cexAe9+BiZeknImwyvXqZGcpQyywZCAXm19hGlRSONw5
iROTp9Pwa9egUT25BVSn+cb5S9PLua48PqDFW6jrzHZnjutke1pA3RQ3Voh8gj2wtMNS6mcjdb/k
J7zVUtZq18f6HlzYcinFzmvhRr1212IZ/qrcVTtZXrnTEZtQPh+ymyT409i2XfUCS6duY7659tzb
uMiFiRkoIv+qqH2u5FAXRhN7Fpy7uRUrePZLyRbDuAKp+UbE5qtfBEYQ7nd7cxe1HV2S8KmOWOOm
CaMjuZOOyS2dLMxjXPji9UNXFU6qW3RFKahBq4zwI6kcxGRMOQtEzqTOxWsa3yUWl75JKMNPIaWR
npr4BMnGa6E91xQLOmPnA/BYx//YN5yuxRxKuk//3UVWAI1WLLeOUF+fPNeAaA8GZybFB9bWXgXN
37xUKWGHqhlK57lRp4wsbc2Max92SVxKUOy7yMOCxhJAeXJXb407ArDYeTFdbtQ4cbry9ntgJrY/
0zAnr0QqE9B74U4QlcDLGBUAtpbxjfbk4zN9he3dKUwqDqkh9WJAA+Y0fUGJwMpWIRL/ugNXlSu2
5+L9gikYw9cVGwoAIPVrwadpYw3Nl4XVuEkpnaLMb55MvM5jB8blwwiX3IBTJBUbEm/RDMKrB5qq
NE0mmP21NuZfhsx0J1bgbQ0x7kf/TymfLnw+Oye2k/Se/jd33MfJ1sv9Fkn3GNrIhqtqxa/l1Tqh
Ei+BBrYiur7X5SfnbdazgvVqP5wcAJ99h73Uz+OhNi5DpKNUtIfFw5fLuK67BYv5tUvaOytGNOCK
Xjy38Z7lNHnR6QrU3iKxwyBcVQTkHAkFthX/OcnOPBTu5jCdWcTjxSvlWejFWGr72U1yWSQeynuu
frPQLAW6knTRDFRr/U8SFN0tNvHu50/7u4b76i9WDSO2RN/1jPqoFyWVGD3fWF22SCCyw5IhEVul
h7+70TKWmTg8G6Z/yqqnP2sClNeoLByI52U3jQPk2DNFOVJnD05zYTaimBeAcONgXMFikD95tcn4
+N3JJ8q+1+UlQlhdZQD3ljHLfEj+PHS1lm3ybjqjbK7nC4cqWh4d06zPtaoP9w0u9MA54i1I8RDZ
X8k7+uRnf61QKny1CGR27BysDomfXSkTF7UNg5GISoB12lEXj6whGi9XR4uZpJCBflav2bFAnPeH
Q8AtRAGiZsPsBsUs5515Dnty35GcBTaL6VHBfZqdPq4H9UCmZtlJ0bdEuUJkK026WRWhMQqucpBE
u5WyjkNTeomQgwcnwgAJ3u8PD/htVLN5wFCD5ezYSYVVeQp4YKzA34SMOSnaIh5UsFu8DmKS4ZET
gxOjB9QXGi9baVcGmTrw70qZHf4A6UdRCBsxMnDF4SQKgm54CCauUvTzNjlOjRB4EKlixlHkopdJ
iTuDLOag6W783pvePLzrSwxJfPvGjRaaPiDxFxR51vb0tzFVSAn1shX6ikWhWkjEFPQ4SFUMSdcQ
EUktUBMdlX2qTTqBb95Jg95GbLTjgcx59/fJfnt+TDV64Mi09Zd521k4c9g0IxDO/oHjbL4K01Ft
CywYI7YfXWPOgC1kudAMeuO0LNbRugv0yldlSIkiz1gy9H5Z2MZx5C+JFNvYwINUmKck/6M1QhG6
fBTcfcpdQRac999WJxJHxcQgFY5Jtz4rZJnzSGb5mxVn8bXHpu5ikBTILyErLGdZFiQ3z0usY9uP
rk9u+0CGRnX3Cuww0Z3cCNhcoZfHhuFp/k561UYBSqT1aG/WzSeT5bCg9gnIr5T2pfvEEXahFi8C
TU1BV0nqXX7eENrnwn547gQ4JUrFbdpNbI3yP0qPr/St1A5yT0Uwpwgo+uU2C8ViISpCe+Bao11a
ax6q2imay46+xl/OzesSghTdgbKb4k1Um6aqKUjPB4GAJwnAM6nOzwBsmDKATGMqH9Lx3fJgHgd3
mkKYThbVOjMokV1vjvtkhk2Q1tETMCIyH5SRMrnYhXK55fhZ8zTxmuBHPueKIxOgnQFMFsnWEW1t
RZmApoRFGJzKFd4nfMe4Z5TGERljpkzf5xa8Xa1Rg1oY34ENOK5hPgIiwrrrrzewd9mYqjMsnrPD
RSGw+3Ykvju5ObIwqePcZ/fgLQJK7/uBxEsar+Dcw7fW3pDa2ArgnBnS8fGwJQZJ7mkQDPxW7vKq
dN0ZZQ92KNtqfoXaZ7bb0A7ETZIQBYbj1/PX+85yOnaZfAgRHdiAHu7bOe2aNIdl3meCjGTD9xZM
fJVhEZsBOipWgUbZXPeUIqgTMYSWHqKE9BCnngqvhWk8QozkPljYPiYCMxG8j1a4Jy3XVuPsBMBW
EcL1Pwa9qN5Pc5/pAoPwDOHZ5qeCQdTUuYe6H3uRd025YfW1Wt404gharlEPVNmqikz8bfb42dmS
MOhbGlGq+qeACMtU/OCGV3rOnkSL5soU9O02tKZiwd8xQFtcq/+CjJ9ftK8JhxKcB9566yN2xDvC
tOogs4mzhzxpOTyOAt2UdkkDEKbXrFzZU7u+bA1uTSF1jAokhWk8yjumer9iP1OBNwbObnn9oa3S
f3A1y1CUr5E6WICT+IKA81oBivFBq2iYrAPjY9PJdFfCoa7B0BVkcCNBgrD9mzScBFFJqRe607Eu
N3K+3jQoSPWPi9R2f7YowSxA37YY2YRpobyOGeC+D4vKBHgLXH/3AdjEXqGbEyhYWXgaDZhh+Gid
e+27og47iJ/qrYUUnGbFvnOMRSFyQZbsijluZbRGBUMN3B8pD+z9M4vwUylVG5NhM1ECojxPEDjT
IfbUWP6TJ1OX584+8irbyyXmHFShxT6jZD7+6RF1X2zxMvjm3s5D7An0LATuRFHRM0c0AK0cfuJM
/H7StlTHLjuliT/6so3ujAhbfvcKMbnqE6zMCCbOHGIS8FOJ1pZIgcWf1sQ/pV8XEzbuY1eG8roU
TKFIi0Al3Jey4pJM3zbyAPgLe7Z4DCSVWgq6D2GpsH7ktqL2byEBhi2J360uN5Z3rMBWi2l4sAFx
tL/jz4dfHZjTqCK/5XSvvQLljrx1WJQl8sLuLGkHMkpNnlc5jNBERONf5vLl2gfkssS5G23nnT5z
q1HA2PBK1vbqwHGVqzwKsW2QnB5Oac5Ky8xkEpapxuujFVfoQeWYKquAcOeOe3rfHiICdv18xt3h
PHRZLltl0UNk4/HZNIUmWWMemWH1m3SPlnwHsSbrs98dMdmG1AioYu0vqdX45Hp2qMh/LFAg2wC1
z7QWN/lER76tJZSD4XFfS8mjqWdPzuwb2gGhWYcILKgSzBkL8Caq379nFEDilAxDVp/sHiGNVj5i
Rpwj6HqqnCwS5HnqVYv1YBwqyiGCXx1VAFMB7uKQu2x/YRADnEyOpKCLAmTLdPd/GQaSa3fGCAR8
r0rGE23V9A4oLYRXa9U2iMf50G25Bw8SrNKq7rtKcodOehvttMth3InR3T+mqjykkhcWsKpfyjkP
FywgLSZwX0nLn1PyNEQFVK98Fm6BgNRylQBk6TkULFlejcYTrAnWTomJ8nKjyvY0zLYw3TtXH9XV
0Rk8ltfAxiDYbME3qY57Y64xXc+dnUOZZoEx67ZWBoNqF2P9gjXapEg/UJRFoOdUm9TzAC08H933
N3mdG6ITrH3jmNVCF1+Tsza1YhRgfNE1GnktjgOvD/YQl7dONw1SqEM/mLKrzV04XgbwictW9Wlg
tm2ieDBirWjwe5oqy5LO9dz5/OaS6jXXxo7ZlNmoj9VId/NKbDYcDBWlMiICJW8GmAsYNmyijjb3
YkpRz4by+fkWbTKFNdbQJRKeDoyXSkohQr1RwCeSar64S3QuYNTK+6oR30NwYzrfZ52InTqMYadg
6lF3wd5fOJJwi3Wfk/XD2UamwM3DmMdYIPCFjs2c9mNiE/5ZR0yBir8jbiKyzkXeaTgvcZSnsXbh
CkTL9ezojeg/PgL3uCWkQLgJgRq3EJHfc00KhOoMRHKjHkI/x54XRfXMHPMI4bSRdgMxw7/WiaGt
iK90OP/+rhV9z4EQGFu2cZIkcij56b6geQQRGWu7dfPXtSfC6nf+POgX2s0GogJVhgZurOqPKhze
uEYzpdK5dhaCj1zK1D/2vqCad8BZjsEminNf+VkbLiZZxZ1Y1QorSYFXSwJvt/jd/39HeDmkkpGt
JbT49nCCH172ioTYn9nSO+Htf+rkGVTYgu+5thXk/9pGhPg+4BsE4tN24MMj4aoSGFhjtSfVQpoI
bUzKRv6/F0/PrYT6f/7TAJRkz3uvgzMJlGcrx69Pj1KDCBpVyfa4ZehzLndLTowQDum9zbPbU819
jhMLZu7NOIKs0Gvcs34Yrj1p7EicdSRp2L1G0jlDWZbNebcnXIiIs05uyVdsxiUuu9MZjdx74jLb
S8GR9eooZd9PrPCJXs1h8dz39Vm9qAhgpI05a7JAlpYDEzGJM5WdoYTdS/xrfsnplN9iZu83pePb
yQm6x6TBmdsuJN+mlqTt8VKknTJWgiIOfb1M4LEdDgx0rAFRanK1B2i3mJ1axGSepusSgRlGAldd
meU7WSsXUCLoSoPtiyNhsi0wlhhMBE/5DKRXBVRQ8AQ3iluWQUn3Jvo5MhmT5Jf4kEjX+NVqYJiN
N1e5AOiTx66xzK1sA42jN0g4K1qlQ1pBYbpxRLXh4XixPC51KESzBf8glSSCXG1wcnbTOfUhP5K/
wXwyohb3mo9McjOjF/q6BE1/PpOAc40ex+VPOzXrhkSMYtUHgTcxEpmZ+uCsss0yN6Jdu4yOPTT2
jQ0NMwoF4PFOQnpGuj/LPFY58OIn0oc7gPgarP7bINg0hWC+ggpdYcnDOA2WfPl0oZDtrvh1a+46
9cVKNUUV39nKlQyiHUN3Em+wGzj3QR/TORxKu5NOsh0bzU5OQ3qZ0LZaEpzXn3nH7N6ImIAq0y/f
pyCSjbcWGb+PIV0CYCZASnuLmTrXiHP9oR1qNtdv1h7gyT/fynu7IDL0mcOQVsbsEVrNkObnD0Yh
qhfsozbP99usXPSzEs1GKt6diPzSqcVqvD32n9EkBEhYqH378gFO/7rlOrKOePopiGdEDjtQSYhI
nZ/FlZ5Coaa6UdQWKxl8qHpFeUgtuNZWqTC/sWNgx6OXXeGxU1NTvikAM31Ip8aDfEvHYFL0gQge
Ekp6YnQHZv+JnJ23ktrhr7ryyZKYQzWK/dykqBQaO5Y5jkTMRJunvr/iMrxqGBIoAIr1J8xFaZVT
sWavuwdUxXz3T3aZbIKqtOII50GIaO+ct7fmgofT5Q/uj6t8AfPbTtabP8O3CNcHgUgCy1QUC3Jg
ONenTOgs5NfMoSTVCgNeKLDUMVoicx1VJA6rzwcukLoKXXVur1WOFYLSO7s1ab38WRlnSj1Pxtvx
4pYi14JEvzaJ4GR01pjlQUqD8JviXg/SVYWyFQ/nlmzoe+uNofz7tRbXVFnt4tLJAmIhkWsUkGWs
ZBxntlLMLzQtHX5ep2I089o6mAAZHKsuNf8z9cjjCh1r9Rq/GpOmP1SYnX969JyOkiYh0sJTy52W
xak+hnke3yPFN8qRACKS8cDcZ8mFrsYOrzjOSVlmqqEDPZTY2J83AARSCD8mYr5VRedgup/mThMT
VzSRTA0x/FJff3a2svVGWuPXtaNtUcZ/kh/V6zg6YNJH9H8rA3vYKfLA2ItfSYb+hIsgdlGj53eq
YjPxk6TXwv9LaCM6xQH/8FLJIfs1/FGqIwYhQVRh+DMEE7u6CloMwWyvZsVuIthMT6NSCZGFKAZu
84nZpuUG/z7t6ihODxV+dGz1T13mVTK3IWa8SPE1Qt+z6nXXSxSEso0S8/pPYx3ww47lG5SXLhfo
vFjDtUmcu7PUBWLay/5DR9XK09+3N+Nif7jJUP9YchFDCpdciGvBoXTmoNmUGvmtP4F4KtHngWzo
nlPMEvundj7HDUwxASebh4rjWhYZP6/u7j1np+ZN3AW1E5AC7OKATc9FM6+ldgISNfKXjmAgCTEg
ogABVQpxv4u2Tj/4cfX6c9KHNuI4gHl0c6weZQLVtK9iEh2Nw9EdGBxW9YwRZ3cMCDIVObnRjfaJ
rqTESx2XKXuGWfJfBG867lwtF9i9x6ECl5XrfLnTtHuWuHWL+WQcL9QhVJpCUVHdI3icx60fIGP1
47ZhhwCigeMI1KVysXx9sEg11ePd0jVcmeHZjk2a6XrjcvJPDOtbkTH+hHNjO90Q9bSu9kuWmzwj
wZ+EvqirIWsS1Oo1jQvOGmgnnP8fn+Q1IIGdIjw/CjYuEMdLtk4+pAGpYSDrn4TaoPBpZmfbcIS+
J9OGZTo4QvxxGvwU1QhDVFChZBxqkbejTrVn6it25CZWcFBwD6VGYvmVMS4KnX9DE/Akm552u0jW
60/wsILhm4hGiEbCsY9AYbmH1RdpXHFXaoUNhTFBFe+vxoXSPYizu7t42InWJrpbmFYybR6yndqL
zJ1LdVkt6LaaHmgZebMuMmMZf0DCIOSvMd6GerYX2axK+Hsm57cTfjQWXuSQZWKjKaCpwcR2hDIH
jfH4GuI8i9rLD9CcCNf3e4gHMNPJWcMO5CcNcdxJNlASUC/m/BRuS0qADaZJ5iZhJCIgnuJqzyAP
Gbq9Lnl32k8HYHA9XmsC5Grybj4BnDOwUK0ynbdjmABJ0ZxXr0IMUEo6sgfbQyPTxjaK+Tf4GZP3
lbeYod2mP4ogfNKPw3vL63Y7GkgQGEbHLpdfF9zj9+rxqZh6AopGeBaF99yhb3lPiFmOgI+dpNT5
8UYhuqMznjv11877Wta2Ix0BfzeQyqZAEQb/9l8jzUJN+xx9pR5o2vu+LSDvgGfYOrjIUhobVCJZ
zqUE7e3y0va4+a7nSJle0YtBJXqfkC/BnR/LzY8I8unYY228lvEFnQIe+1IzqmCatu6BqtZf8UXm
eX4rgS4mdS6xycctKB6PeLlpoYd4doWpEyDE7MAL+KAQH/0eVybiuMdP2+9wBg82s01WmrDOLK6A
onUEpF0xPBPIOAb1H/KQqRXXlgv+mC5GEDm440/Oekj8cO7pkVSqjSGjsxcJ84WJL33Y5A7LJaZh
gAaEtFqy3i0JfofZKovImnSP6QUQsuv6IvOkeW+TR892bkPDxb62vlZvevOTPVnFup+qj40MvLxj
l7cf9m7JIp98B24f76g2Vj1AkbJ8mO/WClRxEzd+lHZ0tdiVobewtexxCAv/or2w8urRUEkonOtB
Rs+jpZmvmzxCZMoG2Z0r5nRCJcB1pUVyz5JL8a15VXBYx6+Y6mObljVqL1vT9xgzAfJEJ8LwT5vS
zA7/JW7wDLc6FF3TrFafPEp05lkEzkWXis5bVZ/FdwAZemJNN07BREIvpzJb1pdYrwvxWBkaLGvL
3C/qbcNt2gMw/jk1VPaBULMprHQT2F/Is2VUOQTaaGyPi7wYvD5S0HbyFLPGThoXuW+oJnMwJbjv
YtpKvMCOiq2A4UzsshMt9nEus7tTzjMRW3rUEwomCNPZ7Nmz6pToRuzFrQK+0Ap6Hbth4XnnFddf
Cd8Kxd9e1JJ+3mKhvr9i82PEzc/OvcJfflS0cYKlKVZsECugPyPvAlJST/oPhTr/x6/gM4aDsNeT
M8hC5N76gxcz+lRwiUGMzq3qVbBrrHcFQ29uJTCgfP01y49L6CU3HowHfDP6yuFFsxKr2rRhq/ku
Od/UCUT+HoGI9XfuOlUuzEK2C9jN2KDHegUq8d+KaAaU+57S9Dz0rHHXCaK8hTf9kdYhLBG98xDq
isb9z3p+wFXMPl9g1HQiqRcOfNlDYF0o81cPHS9tRG7CfQAWk2QZD89rFrzf/hNDRVq4bYAgTS+6
e1nlmbpBTDS9INzyt2U218wXbl155BUX3ATEiKESNwDueTb93df4NF7PDttIqpyTCdOe5vvMdvac
ng/QqeVZrV4idQkWSaEkk8sANXV34AR/xPajY5OyifE0oNr1JUUAvVjC4Hf+3wcAuzcT/1gehgCC
ueqfiPA5HVphsZt75O+zQcEpb6ohv8/tA8yxNjJVplYuY4w8qaB0v1KAQM8H9EHo3lnUoGyfn16I
6a5RBLetmoOGe99GX2P8K7ViVgsqnK3nQ4fzJme/EIqGRwdvi/fkCHzoa/Mi2xflBlpD1Z5TdKb5
Lu2p4NFkYIdQJVuhU+8alBxjRFqf4v6RzXYJBsLFb7jk7IX8wXipi6rOZGba5bTo4h5a2GUwZ3SN
ojsmqv5CSt4AvpCabWh9QFEr4gPTAo9Ks1e6RPRLSRpWGsVjnu3bt0ttTuszEg/aIFrY+aCDpKQx
efEdX7Kk4RLpDaXyF0EjNqatahngQLzZ/SvGGPch+Med6sGurnd3qV5daI8RKx3uV7ZcuIV+NW3b
YPTQyfH+Dh64jti8FdhKCOy/eJF4X8+hAyPBWD8rSA2F9bBKhbk42Gwy3eyeQ3+OjL0HgXpgYnDP
1+5nBL938gRYwzX0AaMFQ6mBJdYmaqfnD6xvSx1u4W3NGFLeiStaz4zzBnrQz92dXR5yxOPr092c
tSWgXTeBUjzq/rdvEsslNx92jyb+JIpLD3bYu9Hyn9M0iuOJrWnEsZHmkhkM6yyarsFcYCgcbplL
d/2ZdxLmnVyPn5L9PdbOKaPY2HMBzbMkZkvLazxOWXj6cagJmud0LT+s6dbwQcW5ODSknz/hxJ1j
6dB7acA06b0Gknfi6GJFrb3ni55vLbjKW0QKexz4QocLTYjljpIsL4BDRotx5HRaOv1si34XquVa
mN2c45fJAMmCizNJs9T1Yrq3nq7GFmiKvMOk4YPjbAfUg50wqJ3PqtvyxumHLREamIjZndS84f4t
+lQBG7JlM773ERcLkyTxArpeYcHOE8+B4lCcFpM5vszHOZr06i8Ugk/WQV6VUPrryPirNuxUw7Nb
ocwCCS7i0BulWF1SAmZgLL0Fg9VbIQllmR5L1sYa9uIEn1JjAmj8YA60DK/ltdITpltUEhJRNTc4
a33H+vb3SSeFiRAXcKJQCtaRTaxrvNxUDHwHRytbH+CHYKfhwqAUJenDk0SLJHrAk6vgpBMQ8qHG
gsxTgMJw6rLDjN6wW1hh9l90aat0yzpTH+minMKQvDVdXHvQqSUcVPMaRqqQhZw2roNS/jKqTyC6
9Y0xrSBo5z2gbM284tp7/k3OfSmSA1y1fv1p/kn6XBTbJTUbpd4bu7L6bPmeAczhuTMztUpWxr5r
vbN1gAd05x0feEXLsofefSOtT4WbmL/VsNr/ocT8IGoDg7I3+l9gbjHoxl38paiDCxPsW+d8girP
gch5NXEGlPWsRaOo6WU3/eVIM6IoVf32ie2IFYxuBosOdDtkZ+oLwTmU7roZADT9/4js+mKFFJyM
WsyOGSfQTPDNbQgxlsbSrBuopUEv8PRxfPyAObv0wxO5cisaOSJDHYlz/m3OadZbqt4K6Yb5mJRJ
tZ446nLRJomFHrdANp8uMYICkmSIOSpGbD2QHfC1gUY4TTmWbFDPHAXQ47mQaoPa86ehx4W8PIyY
HOc6JOUaLTEWXGZ5w1m+sT2dfQcEj2hU/o2Vp42nvcvCFwSxvg+010OOUPDozsiJ/uaOaLk4H0GQ
M5VloonFfJqnksKlaFtgg7PAy2J+KGe7LhZ3ny1+aJ5kZT3QH97mz2dNHknWE7adjU3sVUeOn8JY
M5kkaRnaRLmjGr9ygk+Wkk7FvMlC3EVC+wethBfjEj+eqrjM8VzTN0/tJeOdSMUI4AwLrvENK5KA
+8tNew2Qo4og5OlVrnzYdGLBTznio78KBd2rzKgcHTrTVmHEL3tLXmji3lM689xTQU9RhHxGhgF4
GsHHZ7t0WZ4BXuhpPIV2plrMqXoVOIwqdrNf8llhGWrcJDPX2k54tUO54SfSUIVmEqqK8wVRIAx4
VxX58vUxAOvWziBDUJSLx5GT9f9ueBYjj6xVSM9rdyN3BZMmXdhqUgb0dwACTMyJnylsL/ygdfuJ
F9vBUHilybPtRO/fJp9k0LTyBnk3iI+MuOtl3WX98/0hQEIrqVljlcQkK6ZevvwL9QRjtmix2e9m
j3Wh7fepYoly+dbKifY421l5S4t2TmkhEi4HAJFHEwyeIFS0f/FYsNjggnembacWW8eg83CK1xXq
PHPFFqSYvDrsrvL98SikcNxBP/QucvPfvXqstI4ddas9NfvOeOtg48ynkBDeDGqNxLWem28tgm8a
muokVIdyut4ZS0qLfVX89q6UVT9VB8zymvpZpdcEWPezw80J4XWs3XenW/j221yvAFIeHSgNf+lN
y/nZBL7yzdGG7MnfHLok/Pw44g4O+x2V4qs3/jlRpsdb1GEjgMVckrNxSREWrJbnmk1QDeG6KxNi
S3cYkXhqlztkNpm3UmSRuY+0wqQaVupNF0t8Z08a+wxR1uQgCrAF9CCJbJjkq9iSEkqSPGYRzqWC
D8A8nlgZx6VrM+rkAxUNpqHUqArLK0dZJy+5KsFcYNW9pEAgs4d4uN2HJlXqhyFFXB5v9XkOtcIW
EFJa5/cuv5YjqIew/TZuDwv7lH+DaEam8PjD2Oh2+xiCnXH+snyxGr6CP+H/FNEaJsJ9sOq/ZPI9
rID8Ub+OubjV2iHcJotR0Ksu2SqwcYGUHyGUmkpqGzI8ZnrwxdFJc8DFJjLT19Fh7nS1otRSobvs
IY6NTSOmgK7UdpONv6BaHPDaFkhlEK0F9DWuO1UiDyMipLER0NOA1PWSqih5f0aQi3xeB9UYWd8f
mH5odlW+vcmDsvNhkUigOhBDBNL3eDI9Mw2kj/yiNP5KRFbM/jv8AzLI8GhpbIJqAjso0MWO9kL7
t3CrGDKZSrYYhiJ6Vd4/VZ8+bBXgaDt5/f2gF0P7x7PMNZla79fSXQKbcu+Tdi5jbDW1MDMWYBg2
feX2GvhmmJLVlg+yX6nPqiUWNr5MU+zPccOdK8ZWsdmaUylnRt3lkOGNoQ9J2g7wMqLifMOaPL57
fi+x2B3zNYBeUSxf47pT9Eui7bDxq9ij3MWGBxs2womKY0Yim33VtMzBtLJ2zcIfnkjaaynEZ70d
DySQ6DrLlv78yse5Wt5entA4bekzg6WfMWDWwfjRrbko+vhtEDDWXJ121Zzb+cJt90PMDYsIpm/J
11fchRrO4giwg+jw0MWDEJfBEuWq2TqYlQ8hhklVVnvI4+2cYAGUNG2Fj9h5ZjkfQn0ToTZrUNe3
VKm4+6JjiEx0Nhso3DrZPapmqje+vmy2QnY/j+d8d2T9j7NgyWk2gHJfKgZZLuDnQglFp6T4BMxF
jAuslqc1uWJgWSf5iXSupiuOrnOG4CkpkvX/Iy/RtnYIRsRw9gj8S1RNE164Ji0md+wVe26DwKE+
kTtcbowwZ2ZukN52jfEl35FKC7PUr4YvHkRx/PNlFUxJRJODNODeB4eJHBR9dPSX6E2j5xyKFVXf
3c7amBPUqVMQbJWTOVPeZDFj81+HogTxAKWsgCZIpZHteavu8D+4WnGD2s06nO6ZAPlP9cjpvqP0
ZytiVPKGxv+41mkAdt+5Yyo9jkVBnKDOplbo4px6zZqSIENrxHKsdvnp4UXsN0FY9rGtCE0lxC/R
JEgeEdd53vwcnEmfZZDXUqzH1e+01OIi4X17gnvIm3gPYOCyKmk4mzl+UWhqfxFRizXISz3T4SNa
qIWgwO3Y+ftAKelCXD/tOsi8dBo3lp/GU1XwCotzdKKNdZATYJl1IjaJCByO7d8IMfxMTeRWjHdN
mmAzDaT38wmzrtuPn3uZ6Xt8AEoGM5glX2/eywMdihMcMSV1g0s92yh8zd82HQ3cs7LVdlPBS51c
7LP1YX9sl+hc3cWUEpFNtC9q3VpXPhQDeKcAxGksnvgyQuKYXmBSoPbfRIKLRjIkfOUZqadcpWkV
7wF51c4dvAx+AbNksfQ0KKigM0SJkbFkYRf7+5L4UxJYPnFIwX713LxUXUY9GwIsrMd2XOvgOiv5
J1BZ/G3dIGzXc7OGn1M60WrfaizFzbvWYOKQ7nIlLKzUiMVFHCllEKEX6F6PKhhxU0WPYkj5XOfS
CA8v1vP6MVAi1uYw3xQ0TPU4qawRnzq0LaBhOsa8awArltoMTBpQx4stZVruthMtFPiTyzDB6TzD
dUP+NgckgjUZ4og4Z9VwpledVYM/sC+lFAE7gPtqtUnIfB7ysc2xf2JQg88txYVd5elMqspB9bHL
79ucOVLrd8+iz6vqbU+XYeHNMNLdSzUJG/tLtqYscr6XvnN0QmwetjBf816o9u/pqGLnQDVCVY1M
7SQ6QGt/fcQn+TDM9JUHMck8liyEUbCCuNxL3pGLHLSWQRv2Tyz1K1tNoiDTiq89bxHlPy//cLlr
TFLqz+2UuxS2tsQ8e1LW3lrxjXsBGWEKjyULIi2a8cU8vflCUfbh/HFU9l+lx2onkSW3S98Lstz4
aVhmB9uCjiHlWrX2XzPJIUhopoAM9RYcNK/DNm1TWr76+UHlNl2FcuCJHe+6nXQVhkGxPMuHAWF6
VX9DRkTglodM7A3XzdUoP61HzbsU38wCyHJ2IZILM6sZjGgAa1iedC6r457zqbTkZsEoap2t3yEB
O8xprKOhd/Qey5FqYLXSngX5wOmg7PpfCTb/1o/yOFRILcTcSMLecJUPynmdv/KWhU57YJkCl5SA
9ulIAHsgpayaJ77H4X4YC0UXBFF7r/RgQBLMCi2hyoq+5AIuVUUHKE41XJhwdel0O3Ws8/AAn00u
F+951EDpNurFYnIdSRlfsfDuXrhk55kK/2BxNBd5Ks49f1ox2a9a1H5T3xbhqjxCFpTcuH1TMhH7
ym51ouPnwuRPORSr6FCIwRZ1NFspUiw5Q3HAzu5DrJZpmXS5yiLAjHXFtWj2ax8Ai3E2kVuht4Uk
DA9w2+B5242sPCB9cfVnTwXS7ldQtCwdbSE/s5FPeWWuaSR04KarMgDl8QbkVHGn3xKu9MofMff9
uRCOBRlei5nR5KlU7JW/+d6P0e4iZGGxG0i9+CbghvLSkg9JGDdmjxehUkQK6q+L4pR5Fi5TF5W6
IR01QJiSV3WGPV4/6+OcqO3WbmzhWGUdDW4GWI7PJLwPPpAp31/XwgBBU7JpP/xBWFFm7mVPd56f
iTfQjiqWrEOxFjlHtrgei01hx9Ruf/WgOrV9mJRyD5fHoSBYyN7AjpE/+xALOjbot8N1X63vvKRn
znnzshd+Uedx1TuUa3cGPJb3eAOjbLaqLWpCZmdJE8wbVMNc7eTZ3Mlxo6tGulOHs1vGfyddyk9P
8qFvgfKodItOy0uEazL1spPet+Wqly8fl7DhNzMMpHAxYg7FuDYWvr7mbCT7TLPp2vkxcWUEAz2K
21Ws34MxBMAr6Tz0hWaB/dA3Sl72/Q7oJWKzm5kejFuHTUeGz4ycBF+KaUTPFyxJZ3UJmrRF8Ey1
8E3RoGNvRkPZsvGAALELeuDaL2twm1RE1bOcWF2KKSB8WiyxWgmvFfXBL4q2MAbpNegRewWWzxUT
O+VMW2+fhhIOnhIBO8y6XXpAsLBPlErUlbohGYrh3RVcSkpL1JAHGU41K/NMC0poGEw6K4bSwmx9
bIBg7submTRnP7Hm0WzRBORT3CN5jxU0AAc4/QT2M2GnWzRKpL5ahJG5ewha+4LOjnBYzjLOCsw/
7B9cZpGcMkkb7YLQrFbahQEO5tI21l4gF5OsQBP7Ecuya4GIvgtPe81Ng+XRoyyc05AX31ozh3T1
bNmva3E39YN2UHe6kURhPgyxgYrW/rvkKKFLlMjLcH7ML3lX1DyD+uJO6cXSjS6DBPld0ak2g6cd
RqSqTUv9HhZRh0sJ1Sb5BGm9984KfCs478Mojkm8EhmaQmHvwdNi+WIEQLZFkTQQgKIvJlSgToq/
H3rl/Y88Ss5hdmNFBVAdJQ2ongCNX6qt0oYud/GqoMlfO/5MQad4Zh3ZiHPhg6NBftr3Y8T+XTKS
e5wWh5hHjpMuIxjfvV57/H41u/q8/Bu6gen78TtyT74uY3zV8tzx3YP/fEe0pm6I7poUKTMFjm4q
CqzQpmhRJ4tYsgddBe8ytriWG4FfhKEo++OuZBCn1czPOF4Rilu4d+qJfurtJby4Cotbx+3Wcb2B
CsjORMvTE7WGCPDTGnCkgtaGYZBZA0FzxupSftBlfa2J0FtstG9hNM0OsVZR/sZFfElCL8Bwnn0M
HFpofbjDBlE9Vz/gbIjEXlEZZlDE5pGAr6Sf9vWDdVoT+Of67Wn+5KFabOFYYaUKbo2NuI9Nq0Hm
QBj0Hg983PqdKem75wJF1iDNwgoWK9LZKnRdpZ8RjwaPcuf+3x+bjoE8nsUyOuXkRb68aEnRgnZU
DoJGFIHc3TzMDgwvbQ1F9uKGDS16dVFrx9Ez6Uz5jZkhVPfSYjabzrL4YekprAKReZwuvQvk1za+
9xgBkPWRpwm4XMo8g9xCMzU03ZFc+MIEKmSgw7ebzAscCf6GfzeJcJNdaSVNrcbTJpnimIHrfddz
Ib34O7bXxDMtiu9cGaUHrV4GrLi5jgzXksZ8Scq1hk7NiNwyXdTCme6rA+PtDNhYLOvHpLEqSQMJ
11YjOUwKn7c0hk3KaqoMjeins7I62mztT/y4kvy7t0wEHZNaZw98h7Phshj4z97BXxag0GBwJi6T
JcWd/H+nGXS+TxbmT+nI8TPecAaG+D3tZHL6uzrgB2zJmd6ZSS+B0Rz9hZVyMWnNjP+zvMSqkUay
TEsGynk6rjxTsM4ygRRqPJRF2060B4bhIaP0IxebrbWK8Op3/QpxUA8YBoizo3rf+7C2qZs8h7qj
IyKP9gm9jSADP9YlGiuMSJxT5odn21+MEJT0jdaAKFXOoFU7LDPG1HPW40qcNcJFpjpWjaHvxBBK
M2XrrdcvLIT1JHbPHDiVyLWIharaB2AL6wc9PXvgH9WxbJ9gknnyDLnnx+pyGSuacAOko+td3mcD
ed1Q6FtOK2QiEJk0oQxzoHzkSZLH4doXeHwr9ZpwsNwlJnW8YtXKS1LYe+jY9qMUW2Txey1qal28
nu4iIHJoBPOvdcQ/bQQIRQoR8E8MqGPFSzRtSwVIsMT1M0f3c0ISxgFfEnqD/aKhag7JHA8bc3cW
Uptl3MvuncUcEXNaiP/+s2r+6/k/h1hkQTmAkdcMduJCQ23AkkfLE2JAFe4ZYuBC/9lDEdC5A19l
uC2dDbQRJY07GW6iFplZgM4Lf7tr+EVZs9BfEzBYWEloN65+B73plPwvdLcBZIMN4PU4A/0h4X39
W7giGItjL3drYFrOLO/4YYGb4dTrCnj+lgu393QKgcsFWgHzE48DS67tVyhAyto30sGG6z44lqRT
Ys76cGOYwAdQBSVGqDJClbADiXwbGYyK1yYuA/r0WGVMO2YGztLqeWkXvssTINnpJJhpCY9O0E0R
KE0wn6bWFwVNdYDXG0OH+PfJQOUKkAZHp2VoaQUWJYMv6HpNk7VXoNriF4cnCC8kUaQbMx4xYjAG
baVhdvkWO6dD3EHxS5LSGQhobRTvHjIjZdtP/XQ2awSVoYXCCXSayKiXPZKgaSLoN25mBPcA4/Nw
geDUokkjFyrjyNIQRmuM4+28UksPnKviDIToxRB7Y4UA2/zV70JHA76JwDeOGBfVN4vj4qKcM140
liIeXxKCNqLsrPv+tEBIsK88UwTqgtZ6oWbcLhTNO4+BEW4JhN6Vl+YmIK0hd9ETmE7TaxGlodge
1tCXGM/BEZZizWjzinDz+L0EXkFia560xxF2yHVYl47Fv4oInm6H7CqS5UxByboiDgCaJyP9J7rs
Tg5ZATbX0yH3lScsuPBnxiMSPaEZppzMfMkKmNlDifiiOl3EZKFA9Z6kRDrR78gdg38qrNC0AvLw
2j2/tCa7omPFCdav/yR4p/xHKSRu36WoAIiJ7cG7w2LX7+rXN5866qsf54qIxTnKcJa9qr+poP/U
EDxYfD8CCIQkbKyWHu65eGRURl8wq1pGC1tGZRFZG3eaXMkDAjb/SDkmdcm1kIxWczOdm4lR+8QO
gxtL/KQmVytnrte/mDjEMwxbR14d9WV6StAMB01Vh3m0ibkJedZLDSzQUIg50ULeBgRUoHxKVW4a
nMNPlEhMEj3emzAdwdddx55Lvhbo6u0d9grWK7eCjOVWGVpJtypm/BbrrtqUqT5arDg5h6X3RsdF
HiiLGrEWArVrxLuU3C5c7pimBwGfyijuIINbCKEaFaNfEfMhI9RA7QPeqGv4JlXx85U23P1rJ5Bd
BzwBQFESOoJArmZ5k1NV5t1USMqkpSXghxC8FfpQjn8oN918HRp/LP9o1ZFv5gZlN87qOMPfeF90
NdzZ14WeEq1QZHruNlDND99iN2kBZoh51aHGqrf5yLxhn2Yumr3g8t6tfv4bgiMCMtvugCgrOgoK
DqXLakBESMVqH7tId0KTHfzxwk9jrFay7mYsjxT/0mdcOda6OFXyXbr4cGX7IXTxpWqrbYTg+knw
hnVQ85KMa94b7A7rawQI7spHQoEdKbNp4GSKK8UfNTFuur1l4kQvcO8oToXIn2xsHqJK5nVdgnVb
rCCdrvjzvvFZD43fVZ1cMZwTydN04HJTkOjLMvUG2JJM7t3tz022XyibZX882nef4IX9TwfiWiyn
CN6/mOLPp+1B4KRVqKnu+JqDO7M0GaH13J3OPUfGjAN+x1z4tMJ4DR81fFWKIFJ5nOkE6RXxFehC
HwGSTCjjOrI0k7YGSOvORvqODtURwpSQX0BFh65OEGhdHhMNINRXQX+Cuj0cTgXo/zpYODX/3FPX
Zentve/WRd/w+yXrQVbZ8OI5z53rTlgpwdxy8+jsBixWXD3BgJbAGE182Rpif9eDKXNhIODo9pPW
gA0LLOW7ENcEmOfbw2Xut0kg4oOHmmQOE4VDo+Nx2JB6/tY+Gzx1WadihxX26xB2xzPOFZdOKt1v
hr9KEkQQd/q/VIes5SqiaP+ykkzwmKwHMNXTeZVLtlp5V3HQCRey/0SzIYaGMj3UbC0jdvWAIgOO
l0RQoM79sNPJHLb0CvNAAA6MWbDtS2kX2Fn+FobtLunO2FtnNacKIGJ7CRx8wQdOaqfiujfawfIQ
EFkk1tQJ2kKYid8/nYjlNXZgoSoe5FRkfymj2FkU4aUD6RLquby3CNAirbYjSd2Ma7lU4b32czVC
BRB9A/YaeFSq1BxOhvfy2J5ZmdgErSbEVPl5m4Zclry/P1KBW0eLhsA2G7q2t/FJcAhX1ziuygfL
EDjgjqW0mMXJl7njryT3YxlAB8vVwwgJF6FQE+FpHijn3YfAIU+uoBRajXUeEs6nneePzZFfckF0
vryyETYeyEp52VkpTDDshcgx9Dmpy+1y/6XRKAgsUEybH2wUiwHixQ0M+W1wWGeYQ8Tq8X3hNv4q
1cwe4/QKv6KQkReiBRyUNG7gUWW9+Spnf1SomRMOyOslnMUsWTuyv2BUok6z4iDe9NBvKJvR1sAt
IjFxKmbQxO5Ur3dVXBwUjhDyswjgutVq5Nl35BnKxY+7E2Q2gbFyeB0eugiZjqIm3pqL53FtIkI4
H98S06ABmp6OZtHZsSg4vPhpPxFaazCsHqtB2UsKsu5E9RIHOyxcBhmXP7wad0GZMTInfwKdKIij
f6rUWePz+8IGutl+7tM/8ONMh5mwfGQ7jEhEgV8ZK6DGRTmRgDPq4trVxe0mEn9Wd9/cMd1HF4N1
qRWMA6jwLfZ/2C6tT0PBufAdAL/1iLqO4HKKWUAKGVHV1XT3QoHR//Zj6888B0hvsc8Ul9ZkyeM1
ZjRcluk6A+VYnAvlvJuTIM4FaPRzEPZMCkOjtElmhJ08trU8yJxTQznzaNaUqBAmpdyaxfRxWuMT
MUifYpkSMQKwSghzU0J3HDL0a45yTSsaKB9NWVTkQRvYSqTod6BcJo0TTGHzrYG2xPoyMyWNFmwU
q6m1pxB/t4oTIP4MYDHqJs9WsJwBSlyw34vc5nTESe+eK5Pa0nKlGa4lojf66AvJXikKSMBRJFYg
n4noI6tvyYboBikTXxjFqP+8NhCrWe0ngeBxYmW2GzKwjoIZ+HkMKA72scCmMRFVDSTyebH46aEA
8uqVGpLkt4TosKJ4cxx4GvC5Am7amglKx9+zMiV6hQk582ET/vRz5WjWwXTIp2/ajRONMMBWfLuX
HRqujZ7f+w4lb6bL1WOAhAm1P/VRnLTEokA5OkOy9gB85Xp2BxvlwHaex2W68F3eOvEapgbxCuQi
iB5IrAfC1yU/SdjeJvVIqFfyDYFsA5VFZfHXKwOgYo/VErAN/G7G1eRSfDCka2w1u9sQU0hclyfj
PHuPJsSm8rkS0oYzY5Tp6McN3uZ5rUMQ+62iZm6cSjJ1EykuJl2ZwjAxXUaRNpj9UPfl4Kxputar
YRSPnnBcuYXzII5AFbo+wTPGdTCLHr6fqbktOAe7xnNRIYj9ifx18soNu2rzj9Vjnd4dweNJPg+/
LduvAdaD/HHImWsT+plGtSffdI/g9tGYz3MHeLGGmvIfwDNk3qT+af81K40ASqtRBlu7XVPYi2v5
MFnWeQkywmyjLPyIMma123TeWorZOue6EjiHVqx2tGn6hXV+9HWvwR/hoalnknQn6Cmld+BB4E2m
N+1pviIlJp75UaAP6S+f697olACMSFfoUPLvcIXWVUN6LDUIydRSmE6CvJi4JJPl/G1ILByBa1x2
JlfQRH2jvt7JUpqB5L5WEyUjnx77M0c6ufHslTJ1tVyHEhOjTWgMK5U9yaMEU/W+G0psAXWvXcGE
pRyiub1SgZa2kiLhcC8qe8asVLEqptVhfukHMv8QMZPMyfLPiIyzzFju6fRuB5MGtfn6DkaEtRNN
MDThMxObCHoB+aHIWpfSEA2mGWL/n76g+3uTLNwwLB0Ox24RKD7DBzrTXbmSJxppEqVjHIreCx9g
K1FigrF85yb1qSaOR5eB7P/b/5QXfbafpjaSMR3rOUwH/ZbJwxf0cKdeFXwhO0CDYDrbyWr5tQqR
/FaqrO6I/4Dsh2KuMXT3qKc+jNr3fDoj96cQqb2M4KEzr1Uet/rtamZ96vwedsNEMpHMcQe8QT9q
nHt3YcmNUOcibfLM5ygFI8Agasgts7TWKdHM+Si6YGhynziJ11Dk3GRPylfmJ/zt7/0m708Mxlg4
SQmce6EjOgIxhnISlO1BGm3YDI2qOrL8Ja/oyHvHWIZiEBiMw+TKNqY5zvkyXW70lTitiEDLb9+Z
eon0vCF+55bZxQ5j3M6k3UjvhQuM92ITJ6qj8twLOLY3k568iij9aQ7EMmr+tUfT3ZiRAjmtbp08
Td7BeSf6cTriR8GYHozFxqYhuLXkk18KzUz/wG/2xIheHiAUT8r6i1GlHNZHmH1pehY1QMz7UWoq
mCM+xrk2TC2Nut0OyRgtVVPXuwsyHtUfcImIkAk89pxmU4/QvZxSZy7n7epWmEukrD5cOihjOvNA
Ac3rt52syYGDyV2qcNYQRPE5b4pEPeCML04oj1qNzXJHvyAAd5HFBgI2gJvTxNAL+j2Jm4y8j40t
ioyLO9AYClHKPG090rjgDBCPpmpO80TbE/1rhBwXkD5huGmqDoThPTv74ClZQVQYesKOSJeVvNto
NS8UydSWN90lRsY+zYii6N7NK6O+7QZhOi5HI2RoyrCfkg2F5G0M5vF0/Bp7W5Am5BL8IR7vRs16
lsyoRba/ns3FKezYeNwhsFkeqGxV7VIJgvIXNR9SrS5OMTx6uD9BE7rHLx/YIZUiG6GblUwYn7fc
lxWb2cew5m9nPPc6SGP+jgBN3PXFW58Cdkt65Lv14brO4Z0QZKrAtHTT3ala+KiJWgVDTpnwHTTZ
hKgW5I9rNka23Ahp9w8ug4/Qq1RQVK+Mb7iXSsNIfmczrF4z8zBDckj/lgiEJ6WBDAvKRTCjq8Dg
DXWeQmyqH1M98tZyjtiap8KLMAzc0uHrwjQS8g67rT8DfC9XNPyKwN6f/Sh+FKZVyaYS81KN+hmj
gHUdLSuP+2Sr5E0EjVM0wxMaYTeJyrcU+TrN3LoH0T+mErsknFPhA4BY8x832E/jAEV1E0gZTtoq
g5JyRC5oR3/Q3GPPeEgEWiF01nzuhneAx/SdIGXB0ZMLEV+nK0ljvg32wx9kTkVeXP3meFqE5DHN
9GIzxs5a4ca6PCACdeFEH2lTb9B57RXlv6bRGonIyYlJBhzTSgThf3YSOVCGjCbRDA7W9t/0jxut
r+lsykPSABlz5CdzJvnOrQ18DyLpB8BYWX3J30acNdYLr4WvIfSVOQM6eJkqTIRaICTDoaaznQqw
gJpAvJw6/I0qII37WVPiMEsJbKUa9fPMYk5F8bmS8HIfIoxHrpsUaoBJvfv2XPJyOjRcomxP3/28
Y1xkPrAB95t4O0zdaMp6SKbv+TGLG9zUwFr9300KS+GiZqkvZbB6UtBcyTWxJy9+TwK/8TdLVXF6
5Bprgl4IIeE9PIyQ3kXtrtKdLfl13+6CxQrmY9uQ/gmhGkWv228SdjogzYGcy7HQ4h46DinbvSLp
BxKZ93eSOVfxbteORs9Q+muDZVEmAnRiIr9kC/CSuiletwGxdmRXNfhsf3mWCw9gGFbnEEmBCBEy
RjXKK7BHdeSlG2fZgWk9LuYBtiK82Ds4jq0BAtFk9jMzh2fa/AxFxwKUNYoyZMMHCL+0fMzbPePV
FyTpxZnyzDVoTnx29JIPM3DnymDP8QCBiMKOn7kaskbWiPtRL0A9igdPb7985qyvrPDE1KObAjKi
cAhC4k9xDs+kWloiQ8K+XmtFtNF9/7tyPSsA/cYh0/SVeRwGlwXNJKubHPYT6ByI2m6cnYEmadN7
hrqNgIFRj0HggJ5m68aTW3vCUnNlW8aBIjtFD39Ci55bQkqwDpnY1gQBTBUb4A5L+vuwnY7tPco0
fGI9YMnuCtqFA/oBjq48FxFsYl4XF0YX62UUYYw2mVWAD47rOTNGS+6U1sQQuDVlBoxDs+MrtmcF
wZ95MorBQJmoIb00wALS2vL1VYc9FknoPy4A49X41VLoiEbLsg6U1pl4/3hQxEyfJqrh8wT/Rq0X
yVIhQ/rd9QQCETdp1QvWZ7X8Qn0YBxnOOE52DbH40qZVK4a34plYRhS6YC6sLq9I+gbx6qplfQXQ
M5w4VSj/Y27PzsHr9CK2FkdsYWvuTreYxJsyPJW3XwdS31sv0BcDjoG6eIcX+PAQjULdoumDLSzY
zDUpv4BijRek/EqcAO6An2UG6LFwbPqQC541XrEhAmnQX0Z8StdnZXYVt8o5Py587r+2dq/nIs7c
IO85L7O0QDsZVX+gTdZkqHgNsNXcVDBqEJjh5NO2XvD1V9xbkpeb6K8tgNc96mO9UmQFkddE8pY0
Uk9OJ09lQLi2gJ02B6DPSB3a90xErxJ+odCcv4/jwtMM/brnyRBzlGf0aYOwYMuT8jZ59wMA1qzq
OOfVmCuQ8mJK9zxCHiXnIwbPfVg2X1kUBBO7aGPw73ljTTXTA9WAJDnbWUMekzGmyW151fi8ff43
ObXv27YujPaYlWp0NeGukwuCaS3yfHFuwAKd8PFSSOXlb5lgBjIze7PPHe23/NN+r8CPkotFc6OV
gdJ832l17nc2H9xrnsGOCKuvakwaUzFkadY5c3vNDqQpiBNe8dO3dlPatCaiSns4xaMLPmBoRsbM
wPSXiwsFIOqpGs4Sf1ookfF5XTmc21bkJNrEDNK4DXiHIbvXse3ZaF9NbyDBKWKXeRNtvQJEiMT1
OZ6V5r6pkw+FVZcId858rmpqlgRW7f9z0Q+Vo1z54twMrDoVYhduNPu8hR9aAMfVX0PK5u3Y4zmR
gmKpPu7R3OWzrJCwvCCAReanxnZWXeIeA85mBKhRV2M5EML1kUCoGEIwLNEgotc4v5rXQqYxdKCA
HK3Hcz98iUgdq84da5zdp7pu/4hjPpqQYTW7FfV7jAGJ2iKChHuvzgMIXaJyYM28XrrfjRV1LszY
cGH5s6ulj5SJ0oxAjHqRjQPqo06VapxxQj10PB3oxbZF5aUcvaaXexBxdQKo5LK2KmfQJh6BH8Bj
hHDX21+Hhi4S3NEm3AvzLgtF2agDUKm4phIRs4vCwKWmwI8kIpedr47Pk4i7iB2g1U2G6YNPUxhb
UzmiaID4He/yQvQs1ABHTHppTTvDgGzoI7UW7+3F/zTAiuOPJUfaG1fk7MrHf+EPeVJgdC9fdPKM
52qAe0MEruOmg7maTNwDX4w9DKhFXdLMLiqfSr+1Tog0pxzoj9qbzMhBITMqKiizRV0LOcx/GuAN
/RMuGmUGf7PUHlEfWzHg8OvNbPKOiLJVB89Wo4V14RLH7OcOAbeP1mUGnOVSIJckuqdbqzDqo4iE
urCovfDmC+csyTvaKim2eZ0ya1lFSlqrzr92aHt1XpYO1QrEzWmzy9cX6SfeJl1javRF2NdBQNlK
FazF5nkF0sOPj8PKCxPnxAesZfzIvHY8LcfWBfdlRLM3NxzoMG5xgHLkRmfjWRuIdbYBi6SyLk2a
1uP/wEjsQx/OE3gXQqUD1XRbeHwtgoipS26FdQRszbcOq2YdKrGo5kTqxEFvcZLkOGQJexW6K1YV
cTeNwIQOQOEQ2TCoiEgxvD/3d8C9jjZ43CYl+jS55t8Ubxn/2KDDZ5Tts9nyReeLf+2hwSfGn8yi
bGKLZGU8ikRNZ5kXHGdeoZG52ud38e4eSSy5MLg8VNUXnjhBaxutHT2eMRifJ6ATkog33ezezx9g
ulpiP3qdcB25rGydGKFDl3t/P4/NZRBPMTQk7aeV/JA9j+nPyA2ShuPR7oNfZBX9buzxyaVtWo8o
+ki3fpRQS73kbA0mtdQuRlmrGuKC/DzJSqAlX/nOnTJUOS/2elp13HVTojVrEsYrjlVluanadhMv
71UhGsauADnI+fbet3OdT8BQfRLAGK6WJQSt0eIuogfY5cKgVSdFDYxTQtnQSgePQciShoI+pERf
Wp8O1rFo4sIOiX9dmyAELey8ou7VEqa9mzhyIVVGR4sEjjJhh0oV/Vf3aaoWb8S67lVKPpVNlQPi
aYUaG0MZfJJA1lFqq+kG+qQTeUvEDfQ7X4vNCYnUqnWtnOZyJlaiXc1Nu1MZkkB3ytjn9FzZDLZ7
O8tXQagBCyAG+R+p67hECl7XmmzL7hbw/dJIkWutsCFgyT60IYHtS+CgeJIOJJanxEFgIQ6V+BCc
ABpGGbpXCimTDIuoYuYFAMbo74X61OqdlVvFyfRerbL/iE/bGTRwce5/PEGUOQHB8zxHglt/1/UN
loYOVCdsLI611dV+s6aN86BixCsqOanv4r8Bw/vsIHGJbzcXzmcz6uApM3FAPQLG66zZ2nd7TsAx
q4+prahJEl6+8CcpgSetBAWbMXdSdnE2Zt5AozVV2mCwitGg0mrRYDZhrJB9OcHn3cZ1DwckJek2
Xs/zWFqXtQgUFNh0aGoTAdvxf3f6rhLjFYRm4BJw3VYLmzK4K7TOHoS31sSo6Tl8390C6B+FlWh+
Uda3XTYVZ/GhwbS+1f1qHPSFp96cpvVjFDSJaICBOn9IgrtVVoWZV7SQrpkONjZKU+f+PXspfZWq
cf31/RUiCzTqL3Iz7vFvxWwpYekhABK5M/pIoGGH1zod3AZ24sV6+jutUgM0sNsMBXlUwNaiR4Mn
kAaG8bXj4/3XmS/1OH0RMBldfPJs1Ovjk1xanTNbu3fGCTCHBVEboS5RgLEE352ARv2ahJ8rqn3X
YXvaBZSngRmjf9Nrv8zcfHVhpPZZ9BBMhKbI71EawgWjp2qgkKwSD5OccPgD0As02QMMPhC+Msa8
WYQeqOZRX+3gm7LgY24SBP3aGISZxU++JWKAEixCOShk5S1e8RxI22Lh9M/R5OpXRco17ejFW/+f
gku8yQhPdNTIU9e7J6OJTwmAy5vQwk+gXeDLzxq+PU5fTY1nMsC6NCUf3RXXz7XaSdVInGURPcWu
saSteLvLRB5t29i8ekc/hM0zxEWXc6wku9jMpWa9pa91TPrSBi6VRknxum1pK9Qt96EgLeT2kr6r
XLooEE7Oavy/nFXgsKwk6c6wepIJBCU2f4ACVLg3iXqhlNpPjPWMRH42VXPp10Tatyb0Cz8aMsAa
n196yZlFBgSv6XOEoPjztpG5MvKHhehdxtIMg3i7Ua/Hw3n15QZdVouNfuOJNw+ZusyQtgsUhtkr
EwAJRqwJ+uZskOSXxPZRYk5RsopG5McYvJf/qh4GUdp4bZ2VCrz5o2YpuxlCL+atfWefNPS4PDuX
6vQgJgQZeSxr1WKRuMIKt9IJ6R6jupYh4gFJtg50MFUultcXM/oFE4y+aLW9EAROESeCXrZzTUqU
bETSpCTdqQsN285DO2ys//zioNepxRKLY2UzXVlJshPfKTAKVEKpuxNjlopgfveBFH/LiAR7tHfr
aY8zblWC3TY8j/UPSdjll6SWK+TEEQ/SEV2Xh4IvO5EY4Ymw1b4dXy2R4Q0EPYqf5JX3d1Bpcb12
+HU0OW6i5tsDu/o5SK+WNi9xohYwDGm6jV7lFp2LT//RwRRdWHXTOvxVSvJJVIbvBb7pw02NH+te
acbHGH0Yd3ZcRjZXaYUzNkCFXK3zCKriayUKWHGQJDIIt3fx3oJiTR6sBJr8rJWwiGrd3v43vhKY
Vn4pgOwQ7bCVQ9d0I3OyEU50IG3BJDkSXjh8vSlFiG/4i0rZFR4odNExGEc1zsvoGxv6GDd7wl8E
KWaMnmVgghB73ERB0I/yP6upnvbC7k3oi4u8n11mEB7c7LFPhsO7GnzzJpIdjV9OJ6mPyaW5YIKC
uI40wlRIbJXAOOLcdgLqXSINKa31uee5qt9S4YNS+MZcQm0MW63aL/gmsEZXBRBJNN6Xxt/J36H6
3LUJwS0y5yO6yEAYigRppDtVokMxGBD1vxfCubu7nhcyeCsW8En4/Z7PeIkJpr23bDdbaQHexT3M
ts94rXxOilgwwbNwj1aOjWkk0sWXVkA0JM/wMx8dXY9pBkwNxjmyn8RaqtJNt00M4y2/r8RqSmmZ
K2vik6Gpg/ZHQ5U/jyspedaPNbEc7JSGhFyUlAuSRxxGJk0t7khokrXHvDfyMTRPUIsOxtDCtmDx
HHQ8yKOpaC4AJwwZKZoBRObXsvvWRK9dVStqrrr80OngrTGW++5nb9DspkEDHSfx+eIPpvGaq5Mr
1coYXioKoXtUQdaLexx3WnfEDs8D/jbbe7+VnX/sO96EEgL38iBPeUrPENszF6SfNTQ48Gx1vauY
OuvTz771FIk3jWuI7YtmsneB60gKV8a6LSuTWjLbVjjlwzhfr/WFaauUo6kSrHjBjtSJNELzq5iP
/7yrSGFl56jaHawHrZnboSGrsjuNDIWjl/VVgyNvdPy/1YbPg0l4z3Eeqv7ElttPgVpd8OxOsvnl
utgCxxmuoEJ7yj4dpIqp1BG7OkVAaEGl6qRCdTa19tUSor7ASBX6ixf+R4DaXgmwUOXDUfS5tC90
uHgPQp/2K1GV/14J9z+bM9Ln0Cdz8av7yJjbLst4YS0zham3M2zVh9/+Qp51GMf0rsvX2n3Is+FA
F2YaWcqhVWa5HXlmgbwD5hnzUVnbacET9AxMGgMjVg2LlDB5xIHYOjkwqiLeb3Xr8BggoLrBIADa
bVRo6MBL2IZxIVIyrpti0VrcwBlrGkEl6ekk2e4LxQSNlLRhAq7Gc5QOiP32ffBE1+3kZxybfuD5
fOHDIsSZAoCy8dnW+c4VGSJiH6cPO2ktZgmERXhIdlPJCGg92/7UDg/1IkzdSIW2w8J7CAeTXXne
DLqUOwqbXowZpqppJhm4NHVreMCg7T8RFzQW6GJPpGGjLYw+MHyXKxkqKmQaWvrePBu0suM6AhLZ
JjHBCy1wZh65c8Pc96N2diLz6jyl86eeIndpA+EUDM4MKbcK05xQ/tdPYTcpVdxKatYZMTRMFY5+
/vPxf8j48cEsgBu7+iGEXGEmG5CF6lACCPpPIkSD7pJHouy/LysT8G53zYd9ipmFLiixK7a02te1
OhgPYbyrc9xIF0KYOCKYu+APwg0Xp7vVwdPpIxTnsTfCuDFky+5cdMcS0CGrJuwBt4fetM6GT2FH
rsEjmaJFHMgrPoXs0gOk0YJudkeSs9nnumAhyh1PEqC7mYYuuvR0A1wsWE2EKtcxdShUG6GBxcpv
PKIwVRJ3kPH/sYM+Z41gsVHFK7EgKkgrrFPGix3vzIrfXIvmi9yFI3NOGyDh8zk8c1byX8NlSEX3
uMhypw2S/BZdROm8lqLc08C/iGDHIGME2xIOuI4M3E3UY+Jm4aPzjY/mBUj3vRh4bhugi8issTYS
tgt9T/tgXP5IFp61dBBnpWKroaOH7B1cgRRxh0eWL62o5WQQoqpsoZ0h/LoktK+SmyAxpXRr58au
rRWJna0yuSEOhlb/FLXSkfVaTnqCznBSGIzi4vLsE4zF2NkJWxlbuPmWQqvQeqXpngWA/xpiZZL/
7wRMqyeJ09HnBnHjf76JVBBKLU2wdIcOTKdx0efnYim2pld+D9517/EJKnrF1tkJv5gTWFXqr4Fw
Yei20manr8yjGmOruyIGK5l2pVqve9yzE3jzy8O9pGEL1WHScn9RDjymlIY9lnrlzcjGwnJzCFJd
f2lF4RGUHH08oWACkBGgy/WH2SqfEWYreS9FrtXTdF55X86pBabjgqC+CxRmXVDUGO84LAHSNK1r
zphN7fZFABA71wL/uM2VMBRXCjMedUyjUkwWSZsmQQxdFiMF46BAskISWAHWY/hTVeHIi9gKhf0M
lKWzdBEXliFZXpInzidkbe7r7ZaXVJbTQW9MG1sHq4m5yHQuUN+sYrOXk79toEoY1S50o2O7cGlO
BFTWdyDYGj7CC/WqGeGLZU+KY2SphOpjo3u/n5cTdWNNfqBYJxB0i9HAAqRzS/BSdqr5kmOwqOFc
SZ9OlbrIxa2Kd/3RX2hhDtMeS0djBhSvNQ8paZMhACc4qUakSCQKa4DI1aBUyKTwBppgcF1ZN2Th
Q07n7W6oqIaO6Q1ppo3D3i8GX0tk01XdDHH7l2iVPr4v8slVrpGSyceeQfxwT2+NUIC7rJjnNiPh
P4kCObVlvKDH3A2qNq5m2Fenbs+2e6HP/ZoMWnrt3nD6cYWcgXD6uK6DjC5yjvIEMuw0mZ5ZuO72
ImPKQVKSX6y7JkArzYZ8LZiaNXqwpWyC9aDPQkA3IIxkOBYXVJ156TQ6zgQaASvGLublIUoA1cdQ
6DlCHRfcTNZLoV6iqkAl3ffKOCm0dbjtf5h6nmkxUwrSUOY3KoPqyhJ5yilrpI2MBtEShz8TSNmp
L8/cyGuMBtPsViKOMXqokMrwMwxRwR6Ft71gSGoNOlchsJNQ2paB+tdcz8RYu2XuZ9LjmMOBPlib
UFLl/vAjET/R8zUcFc8UcIpjGzKwJARopunnMpeoauJxtugCHDipC9g0w7K9Ky7eZVpWHo3Z+5x2
cpsCIegs/eywQZ8Y8XhSAtJlEC623NfX1N5K92aXAW9MqtpIDXChjjTCGLHW8vDtq1p3nwzkbCH0
e2lb1nUiZ3S4Dg5IBNS4NC7x5yiWnjbPLpquMGThSEziSaV0mDgd+haNQrLgCsaUeoenTXpQ52SF
PsH/dqT0AA1NGekArWKErUSapzf1hzLtXWBn8O6616KciwqtrbWfyOLKskQcZEDZQlEmpRx1NXYR
pzm6j8/irEA0MsVDcD6KBJrRyymPmrCAS8MNMas5LHrq8cTty7VTB1836ZIZurXchgk0yfl9RCMA
3mpsvvJtilEkIc9/tmz4qQ5zO5rnkL5BhPGwbrtNy4idW7YSrfipZ59UmmMrWCu3akc3GJO3jct+
UCpMBnq41n4vHgCsqbyk5ZxYQI0Ud/rhu7rL8b48WrecrQ+VRhzJulPnc+Pt3RSfam4jOt16D7cq
p9+HUQXH+W9YkqH/1UTLsO6b6Mba7aPljFdT/6iWNZXQa5WTcJ6l5H2Lxw6prp4TZNKnAs4EZ8n7
Px26sEmLnaJobRYzCaAUBxwJSejnQcPFNOB5/yIRomoViGi/iCX1DEQzCwZDoH10T0dRhz+v5hRs
EeVh3TFw5fkBJScak9pzTlrN2PAyiZvGF5RE7dCIgiupDeBDberzbKd2wdNm54dRDdeapwh+UaIB
r7/9/jask40v3Y3e4f/2tyTygEhIsMKGPZe8q6lbmnwCiVGJFVIQbqhEDLOdfkN2Ing1XDj5uqS+
58FwYIyhfjPBX86cSAFcNu6McJqa7AAbW4WAZFXxss760O5MqBD44s3ZKCI3FFyuR/T1zuIlSlo7
omZ50GXRLsJ4xaGZ5lJHx0H0+tS3wh7dPdro0XUJDnBI3zb3cOm0ighwBht9VHhdii93zpZ1+U4y
KaI9/hCOI58q9Jd2YXtxK2DADdUZJHMknRdKhqrnAXphvu1rAV8/1HZZIFkpcNbnwQPbMWHnriUQ
aJzW4nBUFReRQvQgDYY5xKjRbIo92YiVdO3C7pD9D3WH3DPBN/B/WQ7m81im66InAiCX4BePcrGb
9AHkkJCNzyAYyR/pUrUUA0PMkvJBmlB4Y4bmheKYkGDqRwP7nCYu+/5NvAHpbEm7OuasBvMt/csy
JvdS6v9TIstqBgyAGL+C2p5Bd/r42TlkX60VaX2bccxU7qcTIrh8HSVVRlIBAXJKjcZzY8KU5uIT
7Vc3JL5IE/f9PSiGHc1ydAmF2ZQJSXsQ2ptna/biRaz5lztCI9wljKaq8fW0a3D08sgQUSyopqzI
6CyaRTtEvunp4IgZRuQJPkwW4j4txDsnoJVwzLLKwjVggAH4fUjNXxwd5aamZZDuzPIoBxB+CIy+
9jKcmqt7JVKDAGvgttpfw26l1l5/DTv3B0xLbDV4hgFQTFPx706WCzEh0cBi7W/L8n6Jx2mWcgVu
jGPxh+MtAEDHJO/sh7DxrxzPiXjozXiv2bdoOe/3anGeq5wrExIw69jc9qdViqvli1y4u5AuILbr
d1JHcK+p3U91RmzhqW/Gv/I3Xy223piOHxXuWTXbvOxSGemzkodgzggqoqax1DEIz0sM+4DsEzIe
2QNVo1yY7ZdNiJjSvjkGlgZcBFJHIvDN1v6OWOUwvVVoeQ1zo80SCt2M6XD3Viiml1FjTa/ERXva
DoNyjUiTdMINaZWzlrDZHI0/shuv1nbfWSP9u4STBTayYRZcFW+8PlfQOls+xnpAf5fr2Bi7/LEg
PdChFBxW2CboFAAaBYNTIv6cUV3LAC/b7M5Pg3rYb45NaPWQ2y9efoJRRm0p6lcVmdoDuQqP1kSD
s1R6A/HSzV/BrO9Qp0rKpFmBXnNM9/XGJqYo0/XJfynfhgYYeYUIISE3Q0uwptj/OIO4JgJ10/is
AP53VOtnDYeSOUaGkRWbjNkovra0b4ZWt3QmHhTQFeyN+yB8yOugPp8uGFdW2dEEb4vDH9wdHSuS
H49Joq9XQ6LGioIylWx0doUt/kF0mpZAtMidsvjy8YmSjRXD1MObeh83CecdMkOHDz5dgiIJ8VXN
l4cGSRHsKoCRWf0dTDdKG+tdO0UVn4WO6BCMBS4uoItmqpjd1tjQUcgKygAZa70KiwORvgnPwNYz
D1U7walLVFjhul0fQiReMxvAs3TSw2RO1zlcyOe4VExVK+2sy4ZgDTMWCIdnf8Fea/2UjixqLCkr
gko0Ko7saAvzanRPOLdLisqBMEf3Mg48nxBu7PR++gdLZxlYH0ngtjtdv4UvMsaC2A/0ftLfrtJi
AtKukgkWq+BjYrvP4Baa3G/kaJD0dttx4oMw52IK8j9CJyo4VtaAWhc75mb5AyKiWaqwEQK4mHPF
eVoiRu4qvHdXu3EFpIkTjULJoVoEde5wuoWImIYbPiG8Mfr6k4aVkDqndiM+yN4Y2S4J14JhaH2h
rAmcwB5XMBKFCJOD7SAqMXeXqpwak4/dSaD+Xuou/ZqqMigb0YJjfwCi31rTtjvj+L0qQ/dHUjA8
f0lhY2iJv5JsNCrBdN65ItyV+TmWGqp28q/poGNWZFheejiGVooSr3jDJ8qdqmgwj0EKOIAJ9Y13
eb0QdlnNbdNTJpsFcrmsILmLaAwtsrPvQ1OTJhliZP693BFfP9bhLXN4y9+6eDsaFpJ7sExEzTVu
4CPquCbY34OMvKaVKEnQuOAqi8tTx/Rpn3a7bP5z56fXr4YmtiWO/tC3n2PSVmZec2nWhfM68o5M
AkY4t5nYTXSKHqwecqSSVc040G6auDEOoWQogDan77JX4xeH8uDNNMcQHZAEOZl8upXTV1HTTbkZ
VUIeo3k99JD/oLTM0OgwLYjcuXM7mgD6UcbgBNvmmhf0x59T5hiA6BpxJf6Vv4QXAnv1cgBkTPrv
UO/NCmgUfANqLsplPXKkg9Lzj8aQRQVb/pGnA47WSzSXa5z5hPXIc3JYGJzQW0II0GndR6nn1GYZ
MCwrR7vrDAyzxSwtkMewOuCDXiVaGjdaAMogLzLxKB+Qj84qbQMvcEjS9JDYlbQ746j5NDVL5E3Z
y5MbzWuUnCHiqpK4VtFGFsho7crZr+IApfAhPyotzdec81vUkehHy7duikQIJZObtyCGiVi6wPmM
tsKps4FoHw8HDDUSoQTu61QJ1ZiyLXt+4FYbiBIDaMLvX/qV/aM8ywVJ1aO07kcjchpqAnrcIKQF
v+EECGQyNqRU35zimZjBfwBe7FXW/LO7CkutT3I819HXHcufS6SD/9lzTfQQ0yrN/OntZxtOOKD6
L72G9j+NXydS07+KqJ+fRCF0sbYzk3r6aXy2YkbOx1MMdBnuOBXcJZNNWfBnECUwOgs2iqhQoryC
fJvLLw4ZDWGaWxEq718rYNLdyzJCd5YmkuCkEUB5UtR0wekfwzqMxTSjiONq7KbEYPDegecSfOBG
uCxjef78GkcAQXpbMqio7prnCDg8qTT2C3Sdgs4jA5WLG3vlZIV5yL4s7MLi1ycMKWJgpegl9pMp
wDE19csUreNxdRxe9SBGn3rjBK8EAdFfBGha9WfHhFzpLGFZ24ddUkuI9bIbMZ9Mc/wkR/0dSOEj
f5/KZu+vkSgVr9dfvJPPNbgZWscmpqbutgLzJGT9bbC9NdwtN6s+v/EU/3VArWmUPGgAoEgDK1u6
CvHI0ErVycdWHmx9QjlxDir9uzG+tLwZVJMlZ1ap9ZrTeKuBMgHlr9uM8Ux5KLU0CVSpvO+tSbQ5
QdLU4XTkPaX4oz/hBRJ9VLgw9pGvHwJuQ7/tCApiHLE1X9baNjHtEKUDm2K59swWo/cFhGueNie+
1F/eZEu6SOMsRzB78tIG10e3xK32/9TymhFwP7tlQ2tO+M14uP3/DWMXI3Xl3BWPMFuPZAJN8qkr
+Q6xuiNAJCCZIg7RqcLE29utNEClBenISF9PYrVlnZJVD2Hr67O1N/ylEJKiOYoUh3h60Tlul30W
dTIq/akQ8mdfUeVgosLgFv+VS8oQb9n9te/wR0fkKMVJyyYy1kVrlEVa/vSip4kvuFgLcj34DsIY
0BNPSmFgbXA0S7FFAU8VYy/1PIJ18DBZRWRfB0QCSBtDsivgxwUGJmF1iP8VeRJQi1/imafu4lKg
VAEe4NN5hltuUKLD8YiYSgxWyTdpCkmXPkGGPMagpnvpdZl2JpQo6Ri2Dm+5iqWUhllr0LfOF6TE
hpDIRshNylJSPG93oaQDYLEzF5TqfWr4OD/E0KcfIRqDg9Zc6MTMI+NrHnGtGbr2uMENQEaRA3cF
a1dtXessHBA77nx8MunKrXq0IczkYT/7YtgWkOWPjSRhKEzw/VywTcnUts2pHE/WHkz+USapYUmz
jiCx3wvFxP9x7QKH+YiFzeXn8I1guSuyDpBpOUnwxjELC13fIsLPMzfXjnk71B2XKlY7iKh33S1o
m1JMlXKwHAetG75QNIAIdsWZJAZwt5WvMzMQAvq+mxEL4ZmwKoyIAZmsX9vmTd+kliQj1Je3GYJH
VNdK+pboRQYFc/vhlkwkfv6jl7ZVac1HUwaaKyDFtfy5FziBtdbKGSvXpjtsvhJl8FNMKaxYMN1l
Nq0zOGmcwe90oihjaO3EeWne7ZiFupc1b9tP2KOdjoZ7LAghSnibjKZyPFyaLAY0Pa53NP25vZtW
P13rD+ljhHKy5M91tijLxngRsos8QLyrNUvlo/2ioKCK7KQKaIT55D8n8nxin6OSyW1gnqdF2KVa
jBgICaiqc7TT9MZy2P0LVbxbUADE+2fZKW5iY1hO05aSyT8N6ZnHZ/hZueODygTU2x0JVESfoyGV
LE84J87be+vFqpz1uHpMVV/n503lpXuBviabLoxJ/lh+azihUW2Kd/Uu1nbNH1Ihqb3eydC+6hBE
HmsyecHojhQoSkEdG0DpNRpxuOK7o0NHF9AqINivdEQGtFzy8Dfg86RYrUiUvAE0K5Ph1lpVnoWP
r7iPE49FoCBfyqQP3B61nWcMv/UitSKifcJePN81MAA4+RmBQA1iyAEXuBQoknchbU5oN5Z1M4A3
tW4LsPHkVkPwX9Le1sbkusWvbuVw2BZPZuo/8VETMlWngLAzctSoCeYqgXPCk4eWEp8CXP2Facav
FhJ8njA5isHJ4V9OHQVOa6IWSY9pTXvd6lv6PxGbPIs013HT/o0B1TWaLGQ2VmPrwBOxFE+Clzno
rJwgGu/0bAAhRwob2bYMEjMPXYsj1I8oAR9IVd5ENLpT1/JXAjWoWfGj+bmhdwBSAx35OIxvdoG7
9r5+WZ+yMnQJ1mo2hrcvHa/vHIn5rEk2KEHKe7bR9thKRUk+6DfpMejA60Ym6vdHccnmoEPNekj/
DwuTjjYjXtHo6PUH/7Byl123s1Qd73yETzlK1jpmNLn/8OR+A/9PRDvxfCKmcE1r1GzlRPWgtGdw
d6XpN9Gkr4Sco5I9NGDblBhBF0ru8+1NM4u89Yi8HRYuAU5S8ZVsGHNgjpV2cw9Odkj+LkfJSVoU
pzYj5mtqVOgx/aR45KRHaYTqZTUlcBAf6J8YZEeCHjsrH1ZC2TPeu/T5J37zZOEh4mFSVA792aWT
xBL+yV1UkC65MquZTXxRCvim3vTbaixFjfYXy6Wdv3VFu0Muu9zQ8qMVgecXMG+GTZ1nYKWBoNsB
5SnAGOImiidct6a4t0rhbMWs35OlM3aIY3Yi0vfyvsu4L698k1NT2v+P+i39Rz41vqz2vk4rgtlK
2+ElThVLTpaQ71iszxcJ639+55OnXiwK46NbuJISAZrSNoQW2F2vxYcgsg1WxlXNkGHW8UKC7I5+
x1mX2s+CV+hwnEceiqh2dtXFgEZWp+xLJ6Su8RSfbJVLjjsrRi1qgvueauPkH8gOuUviVgoiU4xz
cTtODitbT4OwF6XemU+yVbLjCubND3qweykT+Kbga/ApaQD3MqHOmiEX3ur3aNDedsMp3w4aCY7v
LwlijP7kDJJTwdJdUVwTTPtxgduL46mZ6MMDYO9LtwDgOzwYLjmf2n+qB1rIuNMtx0xPKNpLuD0A
bpZhSudNJfBe6z6sCNYDUOSVP49SEb5RNPbnD4Oeaqs0oBlOwVwl7iFmrak/KgqcopPQuoC5D2bs
Y+WYNUjSIZeNriVzyu2M/LGCEt1w0uVvLvm78eb+G2pTbbiXwCgakMmShbfRPBmspl/4XO2YbUUk
DDfbirvC/H+4URrr3gKqq7Nll4ibKzmMCYHdb4VNkEpUJNx0p5NSil1KbHFLRW/32v4DQnwslIZE
b7E0UU3IS6O5HJryF2Lihx/8vlfB1fmDYAFkS5AWxyu9EiWm7D7wyZV5ZkPVxNFFs2d/LInrNprk
YaITNto4LNItCz8YBc32Oxk1s0X5byMf9y+foq0Gh0hD7gaX7xGY4oVuOsXPk6yQat63eJ1/hWoI
T+hd1M2uABwHjLi75qSZ/5Z8u6ue40fkAiAOHObaYPGqpbUp2DKaOTpRWRKq+lPh5f1gCNunyWTJ
xSgeyKE/1lRjkJ3xpgL6HXWibxLEe5R+6uOMxmWhxvR/At87pKGcr0pOM8BRg6TMCQ/abmsm0oo6
yEPLRT792PuH7ThzTPrm8fxt123IThYuRBdOeEltYwC79Hi0TqQXiDc5jk4h12iG0/N4yEyxpJqj
TAKP/ngHxkvT6fXyvYKSWls6qKm3kB4VdRpzV/2VoDhrXRnSdCwXmJ83jqfQiX++9bd++euAFHqn
BnGjcoUbMfqNVh4VDdzj+UhIkHthNcrJkCtVTJroCYkXDxsAxZAG9F80vjyw2caTauHWKSn3dqQu
K5sLWD3NvG0H5cdrnQqSzEKY9ZPlZGQUhad5GVzXCDCB/Z/76yeitU205iHafhXCifWyUnWsiE8j
TMYdlWTlrjEtAYML8CgnMm9YkhQiVZYVh6IIRUt5tCrrLGVSlfDOGc9mZ0Suv+7NjKK6kwcIOh5e
UuAYbuaTokMAeqzheygxRtKt7RJHGbVYQbZBAtMkdhosij2IoBlJZjjHc+o+331lejR29YkyD70A
1NlI/O3EQoa6TIHMhwXwJlRxXDmNM65DXCkka0cstRWE+gorgR5OQfg9aO05yv+hENEjAOnDtbvU
6x+ha0z9nzV5cwi5pq1I/msKYS7DFipmx4JmvMTtEhb/kjxi9p5WBFuNkz5BmLZ6HKvllwjsapKY
ztjk9xXO66tFT7HfXoZ5BIVateqPVXPtD5r0TA1LzjznKS1MdMqPBRGWVizmsSgCaXZD1koskOcF
zEP6WBIZ3MXZPvQwcjBHkJY3cMCYKjJxRpbHLINDHJ7FQ8483+HF+YkwEeVquvWRfK7hFosNT4Aj
c7xzb7WuXXcgHh3oyiKeh4rmGEAc4slZvOlY25Vl0ZUBBtuMr0qqLO/smz6+GZp2r3bjmd2zuN+5
thT9moghxRzfUNWlALPmwOZdKBWYS665llahPsB90N5gdFB4FVTkV+qo/oUCh4SU7u6pXib7+mG5
T4mgMj6yH/zYXAwclKgxu93NSAvLPnDz4+KGthiOhmp8bYBiaykVnwzymNu4222JbWv2RsaLPV1W
06fTrMrS0fijYpWc5wIBgB5aIi7JKSua/YPr6J5p8zYDwCd+jEihb5p2pINdtUNVAmetxikZ1n8Y
qa9b+qVvIQXJS90rPEMQHtds580/S3TPP/GI+uzsIfL0WMme/9t/sBTH8OBFCC6i12Jm7Gx65pnq
uusqlhGLNFz3metRgbSAs4wsi3iFH7pjYUSlFs5aKrRzi/LgJ1Zjh0YCsvvmjWC3Ubr7Eh7/gTPo
w0tFWJdVmRwFSYgT/O+oO6GKPktR9F3rnSj/yc5BDxLHGMwH/9ccJTFwOzQ2MIo9XHhKHvoqe/h+
f6WQFVUR54abxSNgmJtA0fi+cu5g4qOQYL8zDFL8fkinXyQU8it3htZEZ8NI2KpFw+SXMPTzms9I
i1vIluoc/8rNmDF6rgq/x7S03xEfF9LzthuaiNHoQcHwgIm1SahUg6ML+qTkX+78PgDokguBJR/M
dO1NpnH9CipWyD2Hv2imWrd2/+MVNnF0490K3KbVRK6Emp94i+liTxhdCmmsRpaGGC6s/iP6kgnW
d2KPD22c2EAZndMovVTIFM99Z7ytRB8ZJrDraSfsHfHfluMDMba4vNb5a2h63vE4p8bDvPXgtHrK
fXEhNpRwOyfl9uQeuBhVFUeUz3xVin+5Fyt1ijktgpdzShqmBuUmANo9kyiBdPm4vzcKeBpX1CMu
Eo5xup6F2oVEbbRIP6fVX4gKwRlt+yTXLbUnJs9uysEaSFUAnSvS2EjEJExFehZgKTHvhx23FDGU
IRQBhy3Mb/emNBdDTTvF6NuPrAMpGiJhWrnpijIzDSk+dIUz7PEeyB114LnXj0tWtaPD8ftP+wyW
EzKlgQx6W0ypFfZNEURKWsAmY/FINYuLj8w6OGVrGGszQK5r2iVUiFnN5VZ03YfZKRtrTWljoKoy
PY4Qtzf9Aeg89OUCG/Se/ZzyickZc0jPvvTdfUhNuAg2Exw0OowO7+w37eXjRwiVJDO0ILd5VYNt
kWaeTglcL6WVwjy1G48vPlDBzs/bL5Qb0uFNlBjwoDm2dYSnPHUFpDI5amsVec6fQnRk2eOlqlf/
SUUl3bqyifMkGZMMbeBFWd5j0JHDztDnxNcEAHYji5Yr+TXpsBHJqmFtenLtYis+5QDQ2kwpYUJ1
a7hUwJtwvDjtcC0OBrSgGl0yGY0ZxNrk724C6h6luv9nj1d4eHSklNgNMpiZ49EGgGU7mdzPKq5t
PeOaGbWi88BwzbDhlG/97rsOuHw2qJCl6TNhyCHPc4a6aIABFCYIAyII1soRvYqPErAN071ZlFYx
xiLDelLrxG2ssUAqYj0ZZUXvpZ5mt8PZsenD+GDUchZHnyvBU9RkGz9d7Nfs0vwnwlTz+RIKHYyI
R4uOeyoD+ZgNgw0QbDdcJ5/cJRqqfEPClD16AI5kXAYnV49cmPgoDYANW6bdIPDAlh8kSes2EDfw
qCxlyOH0sEbqrOuA/df6HJQ8v1oSjUttsPfq9b0EWfnfm7I/gEEiy5FSse32m/9iovkWnvKFYHI8
GTlTUBBW0gtyG9trcUptgSGHPo+07yrejQX/VcJdqWFZnvtTVI0YKbEhIdSmWuV2avHvKC9+kv/3
l1kt8c5v14wnjk32/sIEBiCyjHWnbKkQekfMTTq/f0ROvXrjUUF9W7lzxPx1hP4Z4NLW2285g83I
9ueww1jNO0NRt7wPp9lX4stIYn4f2SDRJ8DfYZgma3x6/VsPxoeD+jfMagwPpT2EEhtDBoTi5YVz
f+bsdjwFtBaIi3K6uvtPd601ej/V5I4Zy0DzIWXXwMgLUDi2jBkXMGjKnfrduXgwLukOeXIf7eDo
5vhSE5QvVtNoYZHKHH1flzuYVLK1Rg14FGHfY8oNh9t4U+lEARpsn59GAMcnOCj2L98rlX+sHMp0
+kfgmrsI2bdscW8W+8S3ivv1YDX1Lbp0c+KKMdGfGCsjBb4V/jHtsXOz8Xr+ZZakG0XZY2W2tkhj
eyPOj+yvG+TkrJbgAm/flnHxGSNX8hCQG41cCWkr8kNOGBI+XjpkJ3WJSts8psdG8VzygvUIb98o
ttNeRPidT/vyyVi80JObn3XfJWMGCQV4p6pUMaxZButHcvK7pmm3/FHvCjokbjJhBA9Mj4rqvyAD
Q2DYcdeGE4htktwhUUDbaRBtV2HE0dOVRfyt8WWiHe+B3xVFb/wbKRqDy54Bied/xwFZXb74qdGP
XWTDRrVs3kt/f5XN33isRIHDmlQstQqi04uHGFQuCRn6dMtjrfpspywHoPlTUo28lhjLREn8LNmJ
tvkDcw+RQYRFKqu2pEnwtrGF7O4CIGJJTrs9Az/kSkKdQ341KC3NIVVfgGmmoKW5NrQoCD5OhQ7g
RQXH9bNt19sdASBYJ10yMFWzojy94Obwv2PQ6W2drH4mBzZm6olAAG7VulKj80nruo4OK92wdi0X
UxpNoa+ARmiPkd/XRFHi4HA5SCxh8yPVOytYPzZVOJe31f3debng9yU+P+AVxCRbxkR/eydtzjj5
Ogv3EqwWIUcFX6mPpKFacnkQ7Zcc7zQvY7mEuHmhsVk6h/zPCkThXg47VJCyl4O0z3ppFikbMtoT
5y9WSZf5P4jOJHqmrHl+R1f++GFtvVknESHpRoITzMhuVCBOiqTnN6/vZgDkVqh98Cz+7OwN9YV0
gBIsDAVMn4Vioc44gF5Leezf3l4zKpjo5FkTgbxGqZDyeLz5HCAl5szQFwOCa+y6p+l4hs5qb9FB
xgBwkbXH6L73jazb8vYwyCLacp/8GLXsqTHVhdKYgKuGvS4uCq7B5daJ1THhD2xFWbX2aSD7iFek
9nNFT3DeCLHLKABE9jLmHkzRKmkNry3wITTTtZ2GDgt6egq5D/p9FdPvmk6KNuQmHDC6oV/Ht/kF
e9jf92p9qht7eDyI29AXxijVEoD4QKeg2h5k530ojFRz6hN6BhvuhQOY2h4BFmmvhcZFpj6IZ7LA
BacLcrV7ZAQBESp2pj8JL6yBCluD7JHv7qOPVNxATDCG+vHk3HSMCJRIvaKBJ4YMNNrJUJCeMVjG
D7wMHktmDU3xHxQGEAVX5/sVLCWKxK/Oe1Qc9wwmiFJqRP4MwN/AFsiAaV0oQ6MTZdAWUXG9HaQ8
iQra1JcAS1moWFP8MZDHgiRJ3ECdDBA+kG/hMlFzWnZ+uTlsbblHldcp7l7HyVkbhmRqgVOu1aOq
rb2LM4E6XvhM0L5WjdBoY3Qglv9T1eoGh9P/RQgUDqxUuh2a/aL9+P9QiAAFxNQNpoK54sQBM4LC
R/Ib3XA+rwsgGJOAPiz29G7SxoLJsZwMOnKziRDeQBMaSGxRER0IihDR/fNzKq7er/dFov6LdOQu
n78GIPlAtYXFxLEiOSeuGC9/ChipnmlbbxluZW+jd4MqOx/8NqGaEs3npYsRaPbTRK111trI7xjX
zNpFbfZDu6FSouAXj2lckRg0IGU+VoJeeUGd8AH5Q86qq/DowK/4+0F+APSh5Fgll7sz9/QSgsBL
IWie7XQnUfvxNBBPCSULnWjudsStWbOsgAgTFblAKtkPJvoCbCyeRt/a09tPUodXyoTszLaxrxZ2
HvjyxToHPxb7rAoOnKznAzgIhZLtYQcoi5B4v/DYCiZkaA3AHN4Y0oP8XJdAgSt+mY6SOF3nkOFK
2s/oOB+WgW4UxGa80Nb98JYWY2///AEOMGoalDFg6yUzIbr2TAboV9uTkRtaPG67B1l0QFzFS3gB
kapbU8WNIBgLRKNW6YnsdZQUAF1v22xwSFik/jOrOU4dqd+w52ekjKuSg8AuPPWCMynidd3j6lnO
ZZDpcGCtDJsl98NqsC3lWza9OOZgmo8gi0NF7tMOFlPeI59RT38T5IK9fcJ1bY5aTnQjvCje1T84
Tk4buGeTGQBGr+SmBxa56TJM3m6JMTkApu49S4peUcQEJ/Yn2IEs2CYDwG46x6L7ZZ2VtgtA/z0A
CY4q9e5g+2Xr7IXFe8/SQfKPGPT7gMa1DoCL0tuEqyEgqcrgtaYAXA52UoPyHF1RXYXxhzogUx+A
iFBZHfNtqi6onpCUh10ubNagV2AJo3Ij7xslkSEchozTREUi0dMC905jiEyT61YDuTb/F6Qe4hl/
Gjl71D90NLzk9vROAYGZX0grAFk5se8DPyc8Sbhb6f+RhIdjWAK7VaC2AGsTNKLhbd9UBFRdZxeV
D4mfToBbCT2EsVP59wHIxVS3MUdeir/U1BkOwZZ0XtiO2aWIm1UfSpciZWvys7Laf4+YQ1vZW779
yHauKo729O0D+hy/VW4DXucB1ssa7ufIg+txHPjU3szo+sghBNjl1963AafZGY+yZPDoqjK+d1rf
UblxhPsWnWwdrwU+FVXX2Escw17gYGnQWAK4v4bCGjfrX+hRRxx8ysnERUPfeA3G8vc+J7kmfOEt
hpbZU/V7yZOJlj/lTH/4Soxs12gMGMCcDds1FRmHGk1if4HOUxin73zjZGSh/HUFzJl+PVGEEFY1
RTK5HaBbfbKNtolEb+6wQ53kVb52jILRv4EvpTUViARofRVDkSrxIkGDCED17oNMUAmQ8wzI+2qb
QUPMc9ajlsUebkuQlcewndjw/DhqkxOjaZdMCDeyh7IIc83PxQ4zu0BBfOM/Z0EcfvadCaaFzsFb
7ayV6P3zIeHauRerEvZSgYEcby5URiixVTbvB3qLpXSSjiiD0Lp2jr7UYpPidOVIyoCM9Fv8UZWG
JdAF+CYiXFj+dpvWjcrwqPAr0Oi1/ZPz1+Y/akaCJBbQ8Re2opHqOcWsjyYM7ukZwSb/udPu2pGi
DQpxe0inAeTlZFJCvv3cNF+vbtPTEwWwT8ql00dZIqJkot3mqhHUKHEfZUM7yVLIBk/d3QwOYrLG
XJgVMif/L3PsxmuaDaaNeU4AxVnsgswBw/H9oJ1fh4pgN+pe7S+zzGWk0OurDn/5wvZjb8MK0jMJ
YhTFdwkPCAmTPbUCYrB/QkR6ihgLgIF79AuO4TurZq81HrLb+0NISLBArPiShNGPBK1fP5dVHDPI
VGJj3pS0mYM8yk93PCYdF5qhX91JCIB9IHSXuvBUoLZm2BkeVX56ozppYgl53KD9UoKXSi3BSE27
MWNrMHiC99zhB1WAcifaTUZTGGIYWGOGBLQQNsr5wqBTwqjQ2ogjs+9BJcnLcfCqiTJ8fx3RRbf1
AeowMrGbgU2SAjuUCSkzNuzAjgb+w0LUuM4DYV8aS8ssmVxfwrgzKl8epsicUNJNpwNRUdIZwVeP
UKikjKObw8kz0P8cXT2uFlXT1WGZbqMt8eJ/Y7pyCB1DAjZ5/YLbqf9cvF8mfmPcvvEaoXAAixtQ
8Xe2VwXMKztXNSpc25JBJmGuRY8Tjs463OkM55sx/Rm8xU/1hxVkSZs3i8Z0CaX/7BHcTlqNzt2W
63zI+bj2QmUxuW706ltyKJCwiC8QtZhqyZ32cbH7Qr7nvYxLPkAs7MNdDYiAYz476DdZ38XkDtVD
eaNKR7NegtKpsIjeQDD/bC+r12w+mRkOCHMKh8hK2tIYJ4IkpEFcuRzjDUyAuQrXEbpq0BzZewMq
DbQCB3D1aASbtmnXh04ZRorIZPppTuYu1wzeg3jeIBpVjEOKOgIiAmqG3Zf5/cFMKhYZ3iOAhc7L
aT9rRY/k7u3jsKDsXdAanA5/5q0uuB+J1oixkNN80T75P+3xcR41nU4BwhewMCE1HCppLUloc7c3
GAowbaVByfKG37N/2p7BFx0gpEy6m9wMnuiZ3Jv9jRnRDtgBftRjgphITNMJrR6u4aTRDOTDXkdn
ZMf0zTBxIU+jIuE3gvjutbii97z+fkkUrWRBGVt3Vj0Vhp8jjcNLwhx86swmbw73NObSdfpjcqYS
U9j7OmhQHUNlIwZMmXeo0ha7g4UyH6oUVQ9uB0KmyGZPbmCTB4KA8AFKJfl0favSWDMWcJfZixS+
Io9IIikOp3ojcXcZ7bH4AybXeVhXiSGKb5qPvUSW3oTwT7QJOqmZSomiPaxwFje0wnBmVsCqvphC
dvabYXTD9qbqTje9H8bHA+qHCkGSAjXBfUU3RTaYyVH3mggvVO7Z0wa/J7rWWDBdj3FPoeh6YVXG
l3g9Y7cacEbtsDurWSm65bfcMxd1Jc6GH7kwtruvsNThMNV6WmWlvW76V4LgSdBR8WVg4Js14LvC
/czdvOz97ZwYdDGUX3tVdWPbHYpQ/BudgkIVC+RgqKyqZy9myEilrCz6wW4xO958qM0owUzzkzz0
aE+7ifCChTxYEwm5kzinfmnLO/5v5SBvkKQOINA5/IaxitCHvEA84jdjOdU7LUATygdQM/xHvKow
/TFzvIfkjm2OW48xBc4aQ6+1Bpb8AgxQaQr/5KH6sPeUe01dEKCI1UKznS5+j9TKWztpGMRj50RR
GAjvvL0fmm5AMEK1OZzw/FTfs9R/AEV6yuGu81wjCQs4nYPrBQ/GsZktIegZ/mmf7PO7F0jl0QBt
kuWHjLWPogaNfP+fmk4+ENL6lh0caSJeYfohfHsksUZpKGW5B1ZiInFB2PbOqPcHZ/HkgM54P2XK
le1ilAQZuWHkUMyuYHDKmMGThhuqWTcd1pZ6Qy5b+4nCxDddlGsuAkd7e5pFXXU88uHPNFLhlW/e
DF33DuE67PlJjj+Gi18ix3tlkec2+iTkMTn295PN2F7TAgUlhpikJO9VsP24mrlVHuQBN09DmfR9
ygURrn5DGdmMpQ9pr+IHYP/0h0RPBOleKudAB4Td/vJRelxjX4FUqYxr/+jtZH/Qv4dz9e4El9VL
uSx1Oq19wT53QvLNPCZOwuqwFeeR1hZuwbXSr4wZUGjKlXXtdG4g8gnZdebA1aPLAdfggufHqnE3
zi0ylzev/ukfWNogiV57HOhaTZ4TljnbU1quMYBNb3b80OInKQmW1oMmEPXGXMNFqO3g23/CHz6D
P2PNSeH3WT1mhZkNQA8yms9hAMKVXqStqoQ7jElNOaeSz2LISiJdPJXCZoW5PH4gsgSYLmPJoLqo
+YNoZQbQaRFpA59+bZNWTkzd9dMGuZUgEeDT8nUOoTE5zyPlAEsOPYuURsVd9BFTVaJhDk2V/Su0
hU8Ke+wwAgiUrvsJQoqELeJCbzQ2vfi89a/ppnlv0rj4bdSQvYa52RE6JKrcFhd9elTuIPOCUdfp
mNEMvHmF3XXiSZsr0acmlejke8o3yKBaSBvEThpPrcxsEwQrm9gjxW5iSeQeZJEovCX6+kSDrSK2
JYSTI+PJloFN6q9zgR9Vc00LDg7E2I26k9QeQkJrHzhPKZ3bbUK8aPPXcqj59oI+dVt6xPVEVINC
qymJ8RLc+6wEUzReqeUhN3XQ4qO+T99cBSFkxCGA6L3egn1m00sXDcOTt8pT6HA56Xqnw3/ij/NU
Wfe5yBLptXXZ4Ed2VAzV9SGZ+Lx5Eja1qcq0T5KDHG3o19Dr2cM3X/vnKHM0KMfywABCvF9HWqdF
IMMd8wysXHMpl/2TjEueY4RkttzZKjzQ5c/XMHGKyGturfVzBaQkPugsHd9MFqtI3/ioyXadMEmy
3VQU9RtsLjLXnDHRxBHIO/p31uWuigpulXM6p32V4yuJijrnD+GgN2LbnJr6xjyQBqtraOmjMZ1a
456d+vVf/Ww9zEq7kpqNR3iavFeOTeois7VorgvdKBFoXIJCrTuuG862UOcnnBbqUA88OBdJJFyL
bm0vvle5mrqAzDG6jQCr20Lb1Fw+FioxR0jytlfI/tLMrl0Ds7eJw2NKLoHPZlGdjFpBafjkOUM3
/iXLZjvAI7XfeoAaIXCtkMdis4gAuSrA01TRiObozixytCk/yFNfi35BSJ+fAZ/MZSMNJwuq1GF+
7qxpGEzk8k7Xkk436bUBbHXoQ4PJWN6XT/KCsTghPK1EM5+Bezfxejc2VVBToa1NxQ22RHzYJ4vP
nGMl2RDvVxi/+DfFHDi3t6a1DjsINciQa7iBJGcrWFsHV8bfWzxe2wCmPZfGGoT8W86ZXkARynzv
+XMhjYWHT52f0G8Jk7tlZFDJpm/7MjqrupJ12AJXHVVhL1+3ovv1wU2piwkuyAR4Q6Tp/eoR9WZp
0Jd2EzbYLG+RpZ8wUd2UPdolC7BSIA87jHIfDxqepxFjzpA+3GOS+ZWf+SqlNZTsXNk7/6DHaAvX
Lr1nJCO5s8U2yeDzbO75/ID8KdmVF58Jiyhu11bIII14paf3JKHKoxSzxN+sr3pi3kmWJqY4UnWM
NIyeSIymBaYXNx4kYEptrNC8/j3tb6GOuBExAIizghTAYKpa4Ut9JkJJPxfJdHi4H9Z9SETaFLY4
eAzjg1jH3hGhZM8ypHR2SrsrmmvDm3TGcJszE8sP+KSd5UCfQT2/TVOdz0OXzXDtmsgTuNS9Paw4
pwNdMkEdlCCnd2Xm3BtHCGQAjk4JctKI/28BJOV64w/F4VvZQ/dn4q8USxcX1to+raXBErL3snNn
f8fjCyLLbhHXPbv7ZaOLQRmJ2A7NE3nmjEuI/4MxWQsANIMlHN1+gbZjitzBkRuugeyWxKtn5M/a
ySLnRyPnMkFu2KmsIvIwhsKDfDuR/zxa7kxhGC1zhXJ2WU+M2d2Qgjymb/UgwEZJTWTkRUEOn9vq
DTVjA7sfHHaybxZCa8ZBQCFqTgGQFlfGRBh0xQTjxeQj7VMsoLwv/CUdoQXp0LO0q01YbeUCWzTp
60nAdY9wGRndc04ryn61duUV5yhvj67teqSD2U19LwDD6sg6Ym3Ybt3NRIETPjfA0Ashb0IRF2Nj
IEKMkM2BsCbk3V8Obm8JkYAXLcTanHjbALcPVnERoW2rX2ZIL1OhNYaTmCA/t6AZBJEcdpaQuhG/
K+OCBmh3WnDd2dYoRDeVXHj16TL4Gb1lumoyc7AXiqQTsCEuRceQVnD6Bjo4UqyO7PLXTEEdfg8I
UQ1ulNN7hJiOSFOmcNXqyPIrazEruguxeoCtiQHUfE/0C8H3z2DWuk5x7bDFOC4GAy/f8LfXeQQ0
3hWULrTb3PJt+nYeU31FOt3WZgSnPwHkzySi9nKAdDcoJ/Dswjn86m6QhKStHS4j/NrMYvN9iGc6
BT5VVXbrlXF/3Gh+ADaqJgQGrgXH7IrCE7gLaYM79DIxodkiysYK6BPPll+iAwdCRVEbQXQZ2rn2
TbS56huY/Zr835ChLQM7+7S4oVh/206ypEH1CnrCQYE3Tj26BofoH30P6u4JEOxNm13Ml1OgfrnF
ATKGhlXz5PiWW3lPvX51GgUUQ4B17WIN3Wckbh3wxOpTTPb3ret/w0JQPzUgGbUUep550gWHAUyo
8b5Tpt0goWHLYmGxJP7KwC4FUEeUO0uZfoYP7nIThdUwlwM+GUHYRpOIZjJSPmbyQ/wtyYCqidce
11icGdEYl+ujdUT4xvDzTpjslALbRohMPubMQyG8hdP2se/w7jrwSv2vurW9hmNn+sQ+WfpDdHjF
kphnTZ32OoeYScdbE8vXTjFgVNkEZRzWJyicjsfaoShUN44xiVFl/AfQRqG44xbhX4gvtDYl5Udm
ftlbBf2Wgxf4r6VNvHTly75MhahoAjQENi73Tzt/9CZpabnlTE3qEDGbpaYPlhsBIIfBhbsOlPWT
Qa3rZgfOJ5MOCWcfXN+mLw8E9yFcNYW9AME0PzlhgVcn4OJQZEVYStdpUElxFkFoO4LvytsoTQ7g
O8IeJvO92/qDOOn3ILWg2O1UQhHARRUAPBXSYcaTfHAwEMusDfEmCTCXicGdZ3JtbM3mU4q1I4ue
bHBLOHMwadJii6fA7QvS3jI0enHrp15EkQRBbyczd6v4+wuKzMO0CGw99OtlIZWX06g0FR2Kig6L
0Xpm1JYZNpc0jPM86zjbXeVvf+p1oSOaeSTL/0Bee5nU7aDrVE5eVlCdWMzsGpAFEr5n9JcNhy0q
4vHKGD3rM3zztScr5IdZDM+nO7UmszaBPC+L0o49zDDDH1Odk37pb3XgBEbo2Fv+0BYuc280TeQ/
E+ZVmihbXucfm4ELQv6iHrn3srZKlCKScwpiO4Uqfwt7C8m2/b2I4NW/1LbTw5uptDjPbHKti4QP
1jU6WfhM+AJDku3zOzee9cM/Grg5eJzC1tq+Wz5OWZ32jzFF8vcvg1TlAtkJMVpZcvy9/Ijh04QM
CMAAQB5CPYNO0k13LIW94sGDUlglXvZu63DEen+zSOeUxCYG6bEf+l9F21Vvg51GTV/FLExl8FNh
6M1hPOPWME1Kb5LPPX7D8qhUlJfb+p3UVI7d+SVW1anUA10aIcB1OuiroYAstEFDHlfXRb81yzlV
REPZEoofmLqDjlNpeRk95JYYQYYY3gRfon0dCuDtSx1o0gokf8aDbkXCz29liwxVmplEIoXtHc4G
c6muIzimwLNYdtLSCjhQp1+CeD7xkqawEes/LADS7ifRiAAgAEjlqx6yhj389dXxj7fbBpr5LEd7
cYNF2631XeKEXoyimK39CRJg2lmtIXcv3nHgItVkZ9TaleD9DsQTpGBlrSsYnGyssSJRMFRHGfmL
owWYWLervsxXFMCJm/MZLz9haj1tyYVCurh/vKNbjNVKPApthp8YkpI7c0hUZQRXLU4zHQJbbTME
8mA9w+rR2JW2poynjQqK7PEArvx6CQvkY09Ui+pdQyzN5IVU5WpUu3+vEhAFdUV3sS4n0q1rmzcj
xzFeZqeKrT+xE2TILKXLXHFPPtR2UMK2RICG8vpvUmyX/VOiSPGH6JI025+1YP/cAbmyVHmnwbcE
F6CfEGdGL7Ns1wTbpVJxRvDugw8wrjLWIx+odxljWUOPnK64iww6bLRgJgyCr8R8hmsdNcmgZ7Fh
Hf71rfdJgb29LoeIAggMJQRKUTkHV4KH1WkXvlZFNe/YLky16IN0HthqkuZfXsZlbSmmDLYOfXwm
wDP7CfVdYKa7zYmIeaWOVKBR6+7PXDsG1AHQ66CGHX1MI6YIfE8mRTZeARVUfibRZSo56Wl+qMnD
0D8YdH70KV5ia/YQ3TYuW7GA4H+LGuH9Rc3Pg8GwG0EraDssNaO5FsRXSlVuUDQoJWTwNJ50j0rY
3Y3SypI2zS5gCzclLkdXSHc5JjuzH2mVW/1+9bYSks80I4b/R4FhHomoBsZNu1gMYoxdu5KoODH3
Kak4gQOJI7hT0pdAoQMvVxNgEEiytaxoMSEDamn+QjyheZ6rKzs1O769mE45nTXup3Z/AujIiQby
u2ZpPtEbNnfgMmRkDCSMsnDxum8KSzmS0SQoOO828P9k+wsnYYGfaoio5LPKngSpxsFPlfY8N8Tt
Osjs4J2cKyyKRjJouqcTXO2SfxsGqwFqH1T4w1EogYZoR6ia/sa/PlITBycTt8enVWBQf2hS6xmo
Ng5YnXgtTQxIY/jenujBBrrWlN7d9nk/VN6yCPjddjqpOzOMDtkHDAEMtlGLR/MYc9kM4/0V32fQ
Dzhw5hpP9rEtOF7ZbfpygMce3AkGjcoGLbrwiSwo8SFNGuTw2MapQIdgGLM/RqiTzBcqtIMEI6dz
SBxm+aKHvJg3xEAcg2E69GRhJhvqPAyaLOByEAfeu9MUr2O/JGB1ibGr+zDbD5eKA0YR1Dy1DZvs
PnYFVu7gTsniE12rRLkJs9qqLmgKcjq+8YiEzvjX5p8z2JbWV08lCGvtaNAStrF0MBtogx61yGnZ
vUhkWd+uzB4U649UII2RKFiQzKfYuSbgobd3BHluFmmGuwCIdiuKC00BKK+QbRt8y3QEDxuVkeGN
r5hqycfETwBlRhbhf4gZRJQ6E/ev/zKa0KUeDGAULWITfLWoKlGUf/dncR2fBbGX/LbTjx/CokOl
+OD8VWAXZjoDVQwqBvizZ8Z8pPEwY2jLe3lZzj7XlF8OLytAaNHUGKUVq3qYJ7pD7vXp2CL1FMn2
4q569hrxL/YAvtagw9LQ/3TEOWaVryLZslJSZ2t826krCtgpuyzJjq5LO/zaIw5eaxwFwAcV4cmk
lIdRrgPg8dSalcwtxg8SnS9yckkiBe9MiS8MvkmAmLCRCxfhxahYQQ+jD+vFS4jmbtHYQkgi7ivv
4W4gu53ljWpVsu74PD1axZiRX9ZYXzfhAS9CB8SMiwqpMMPAedEd0Jfw5ggzIYu27LERSMobUE2D
n4alh9VSwjuHrcFWlhvWS/rb9JaDM4OQGqpgpiruE022EGOxqeH5BhRq0kIwRRTWtRaEATKFGu/W
d3LE9hbz134WTOxo74mIpOnPp7U0iJaIZBI7SehYSn5u4w6DY0k4sSfXf0WjqpbXE7A5dvCSaU5D
kzmcnzR5WVkjwEblK7TqPbBXN4A6ssu5dMj+ci9QZ+tiO7izL722n4zzd+sq92WE7wr/hrKAWDu1
cIOivx5Qe7uUfT5eb3fmyeAQX42LbxHVZjW0rCcZC2LRqtw5lv41XPQWGZx5C0gqjpYCicXn3dDV
atfdeeYsjh6AYj/xD34k3CriwQBQ6fPBFvkx/O8iZdDI/zL3Sh9XBajUjh2f4tFTSEODUPM68f2z
Ebc0NU89jIZBfYYE6biFYViONf2lJoXE5AxWr1IklyEY3CU7p30VqJylu4lo1bZtqvqzlnZ57Lbt
He4IXhneycEUcrXMHOxfTzIywUdJp1Ktwy/aek4vySfYnOvvjKrWcsVBU513OINUPPxAlbJRzDW0
Nn4fwAkW7bd5CKhZN3CjPONQQZzRNzCrkRCq6LfHSHUe/FscW6K+xZiFA4sn2V+zvvyR8N49gwfs
UQoOKaaH62UE8ifIdbujja9VF7smLWmg2Zw6bKjDhvfCz8Qk3PaPpERkd0zaEbZJjEgJnMLXJUd/
9genPbXTqGllaisBUB/c1Mi1avexWrBpxEEZrs1fv0oDwUululjk0LTMQu8ejpD+Ry3f9MGC0FED
jAFDkQIYdvN/7PDQ2SAhz36bMyrrTrFR3v+klD1BcHOCwKtIhe70ewX8MyOjqmWFq41CvSOSgSzm
ay+hNhBkkKbR4SdvSPjQKbiCpPpXryMDjlZU3GUBdz2Wwzk7/wD1Q4si5SNLCAP0I0PAR/e7WkpA
ksKgGJVtUDqURVKXFBwGJAms5UH60WrKeUCGl0XTnTP0ru9SFchv/5L+qpK1OV2DJL038LAzbMlj
bB+UrkLbx9hLF/S80sTpTH7Xhy5edwVVC1TXIUtZnsVHIr+MkYFDq2MwsJIGuROBPrBFJDA2IFdU
H/PZjPXZqBwda04HceWm5LWafFWb6ywPte5KDHDYhsSq0TCnzD9EZZOYue5vnkNYNfZsq7ZNeXHf
W9pxtOQBGKYiGKW1xhxJ1kvZl14BKzLTbtYXdxllL0Ah/LoGfn2OdvqMYA/cEYGxkEdHLhCac8cm
XEqtGwkhR/Xj8dOq78K++iRb+TSWF4YrEFXrNF8rrMzuZmLrg/p+BcS+ETENU2eV8G/ApDktp+il
ZTh5MfN5aj8Qcvn3mRqTptd/9AtmOhipp4iJm+4CHsiPeTF8oN+6nNymw8YOBvQSBCLm0KoY8qn+
qUOfjLeEs07dSPUdFrzwlfgmRqUdW60m1u2vh322kr42VbMhdcbW47DgvrASbn8D6M9k2Cfmx/1Y
x31jikwmBCSqK7cROisWG35yfzi9BSu48FmvNUMoT19AsqvsYAjmHc+vWqaFJB1Wtt8MALu7dZgf
gJfpTnjazMFNUdo6uPtXTtQBCf0GpAqakjnSa40a+ez3PyiElBfObxlr4u7gj0GClI8hBvt23VJ4
R/veNQF7xqGburZ2qYNZnWS646A/W5WOK72W1O7JpIm9lMIbvC0MxFpVn3a+vaMUu6AnvgGcmA5I
1fd+tuXL6i2WvSb8cV4ZmYsaflPdaILd9gGJ5KvrgLNrpcbmVFDEgKLlLepuqSXmLkVIIUB3vdOr
8SzYFMn6fDCBV4+8ZtWwtcD++QfIWANNJk/+pDzuYQP+4JwEVpRS68JrTNs6bsFTVECUDjCt9vA/
bAt9JM3Xn/NMhdzTsQU1j2b0um6KrA9mWYX8rFEvBz1+1hbuyS3Yd2s9AKawdSbkpHq4jERqRWLr
UnMMQ+Skfzzk1ke7mkqRqQ4YbqSACWOFMAQVSpjirzSAnx3z7NkmxS/pp3KglXF4UWE/JJkpyQ3w
dto2jNH/MwT8NMcF+UeixJB7VnVsZ/U4X+QoV9nwbUWYAHThYBqt+ATpsronOUMGxl3kFmkwhmrl
uzQe5Y992DK42GPw8vyNwu7nn7NPbXy7nfcJN7N5a4Df4+ZKKVrtKTOttCJUAkjG4k9jgCik1pfK
CDGSi/1BP8q9lebMmgOn9eNdmMkTm3u3o4uw8Yw9Uj9XNoea0pMryJOV05ur432BUDVJZo597Dwk
p+dyEHyr1h8Ul6bM1FJ0eKbabPKEQgh7A2ZGJrd5vpME5u868RW7l7gwOcdNZ41NMuMvBuTDbpvK
OOSH0oWKpkHJkZ7f6JEZYs+Tzy9dNhcmHv2pMtSdpLGBRfpgPE/7tU71kUiOU6bQ5Jg6U4rdWVsr
U9tU1ODXtoyDF2x58Dc6DAzj0HUlMF5g0hEkEtvvvsWzIV+enGjO+E9hHiTvy/OP7MbsGmWkGSom
GCRDOCeTtEGg9UBU1e+Tcar2gNh3+95/QLrOCCDGOs95AFi1PnLOS2qVky4eZQanMTDUTzyT4BMj
r9QhKnuCl/i8HEVxUtPcyiRLMRU4wnHPZxpOqdzsRuwRCG0cjCwMhoyt/S5bL4xU/EhQZUqnNQ8a
NV7yvaYJ3mXJpj1DHSyuyR8aM3+r6gjhUg1RSj6gcjFVQEGGeRP2NktCq481fHxJPnsn5bV/owHS
iQiQz4TNAhbXWBNC6KCVYbjLAmNKzGIelGV5E79tO7AeTHZKUDLwSmEWzfrmM13Dwx8+GLt0xFMl
dPadybfcVZ2XOn3AQC0yecF6LL5MzdJFE81Ebj0IX5IYvyN6pqedRvoRnlV0mlpQuGKyc3Zuq3wp
ubpir4P5UV7ThtiFP0e+xQjMi+x5ua+o6AopnSLoCVW+jAxGXBsOMgx/LcnbKhkHuLR404EL0ob/
++D+u0hBUGT6uGmmdfQbtW0wwwCM6jQXChPbfUlCO25FpuSFhoSQkG1vu8o/P0oc8B5WAV8C7YjB
fY+BMtfpllqR3/lNoYDFqkdGwvZYF93+g4DTP4wAAzeoHqejdDSL6fFg0AZYL48xRAzcOgALUozn
eoW80qfycGCkWt4ZHIKDlkJc76JvEPktheZVWUWFCuQTB7lCgWjU3viuDJbwPuIbH+B7oRQsBp0x
Rscn+2OmzUtzC2V6rZdBIgqaHc1chmLuiAXPjaen+kLHHz6KWBhn8p/lGqbPDTDJ+/P3q6Zk8dnX
XVhPonzhZsI8k0un6H1iPU7dO6owinnhLcUp3rzV4WbdXcAOJ2k3hBgDJw49gr1wKVYPmskjTiCk
T9ZOr6W2cRyVKmLa0gkdyUuZbINleLnmkUce2bwCcuJCWebw6n2RP2ZfzpN+FhTDq4OJAjOqDBBo
EIFlZ0zhiMaZw9KZK+h50Ds4CRxKBt25B8bfCZc4vgnbiZQ1uY0L8yawigFWt3Md5LxcRNblkS2l
wZw5za6g3JbZSylC1xeRMLaIA6ys8XSoDxS6E2Vt/+Nr2PKkur8YPRa/wPBGP45hr01Gh2TofKeq
6Mf/T/yNx98lqgPDzo4ghHAvBxSl4bQiE4Xezp7zraVo7N9HETMVorK23V1vG/mnqO6kimrKyVQt
vY3yvAiuvYTV9HlkyK77lPWW01u9gEONZVebAlSSnLTuVFTi5jVKWyMViNJqHc0idzfgTEnJadtN
vNgM/x2w5deguyzrFoeMjXMx7BswN5/OmY0AgbkzT3DdV2k3Uz2eutnY2Rb+WQM9Toh7EJmw32Vx
Waq76CuA1VxD7d0HzJ7l01CU5Nh+mgVT99dh/P9NKd/sanlZ0mCpjtR+aF/SYsn4dCB2sEJn7Vdu
p9wwCbINaSbGBHLcxxwA8Ckc+tiJy7Zx1xzJtd5O5wxFvkQhX6XyZzZwiXwcridfl80/NG1ccIKa
SMUJo8pX5X+Dl+oXYdHoR7QhNmsaqbhC6LcUdt6Fyn1XlA7rBJ2TbrDJmxBrjlKUZmpVypAyeAvl
ba7QdiMtPohnMx0spH32862sIlpvjsa4KJUoVDNSwsB6vpnTvj8JJong2ow201DEOdR4dplznhoE
35lLBjdYqw5X4rinN4redqf1o76rpO7cbXbtJElfpE1MlMDBPZsw8PuLHcW5Nj1dPfxWalQ9Y7MV
tJMD7ZwbJjO0hFtKjRD4Z1+bo0V1uWvuqKFABQOpKwKBUhMmioL7ivPHXCqyzMf6TvHuC/cahKjm
WG8r+RmJ4amSk48NBSjAlE/dvD6FhuUVr31YPJUs8ZK0O1QfuJc61JLaPPyhx9fYcJF10BSCrxC+
ZcjYy8gDOsHrWa5SdUSyFQ4wmfMpHbp43/snuSziP6Kmhx8iG6lno1eSsSi3btVZi2H8+tTwCHzr
6d1I9wY5o+geAWwim+pJDnjqTWt+ODV4TViq3tphBlu7xTIvj0d1Pffnu5IBF/u0TswT7KfxkkQs
Ce045tEHOBL1bn5NaaPvtUHlXWaiWENe5XUfXh8VtWIi/BjEY6ZMao85pjgDpBRUPGKfQwNMBG3Z
sVg9pXeD32+RFEoXtU9jc7HG0NKCWhuT/DCzbb4DvFOqc0EJC5wa6DO1U6bLfVGLFf2WfSoTrhPv
jwbGVSY2dxm5LVgJ3V/l7s92DWGWmiqbz5FpEf3KKLZm9Kbva8xb4/tybipXofdqSGeAVi4J1TPI
BeAdQ7j7jA8/BOtKJE33oQ9sr0DkIKc3LQWV0j7WbqbXyt4Sb4shmGg20+yV2i0SEWJU4Sa86N8H
w+I2EEI9nAmWqpldw4y12Lqsg/Oc/U2IPttktiLRGuOqGYLQEbvk/cKJFx41v8mdFCISJYAjrpdT
G2F0H+VdlpWqnTzsDTYEt74bKiXtXCwZzmzZ0+HoCQDxPGl1FB8GggNgkohtZMiv6Yuv2CWZTxr+
vCb2GREtXk2XEFZBO48DWG+CLEsfkF5avHVNuiZ+1HdkBHubWL4Vgp/6JhIbPyiSE76YDTtYjgGb
LlFXYp1wQ/Qkhmq6mN3NsFd8rzSe1shewuK0aCWGb4CFLAMXC9uzrEByPH0IM98AIKKQv7r8dRcQ
RlxJH3KDioiOHf0V+ihgcpLGna6UrZo/pCr/MXNDtL8t1bead9hnQpROZjD8Kqd19KZDIkHhDXsy
NpvxqDG9wexyUAcZvlCpy/XogqUiq8DVmzbOMj/jEXGUF6CPGxWvcM28B/aGkXJgSNupt+/+5YGe
Sx4ndDsSdxYH6TxtrpmOJeSIZ1g48OfSg8EH6r88ZSGsdgPpCFxTqn3MBIcABN6Y3y5M1Y3fS7hd
hRj7tnyUNZJb0R4vgjBfIPQ5PerPR1QKnrDmcsYmpvNfQel37QeXj4WCGAZB6texi4QCwOQXZWXC
1uTteaQr0cZEFeIECZf6BrCA+JPcQq9UlSd1Rmv72/XxP+vmZUgWl/1oZ7TaRCkZdFWrmPQIgZhF
DTayG7V3gOZrHzGNI2c181os3bXcxvmaS9VZR/ITwq2u8guTYUxJiqE8VHChpU9uAiNX9fjY2SAJ
FMpd9y7paa5zWh8Xiz4ANSfRoL7rc2cEYxZhQ9HwnXJMzzUs+vk7OdCOGek05Tjr6Q4X6DqdvZDU
UFpsJJP/Q2W2TJWospGW6nzWc64g0dLhwGzMmVdlhCPPVYFiMy2URgbGVC+NscgOwU9Ml8c8a3Eq
Qen2+hZVAgw16AyPvpviOmZo8da9jTp/BfkRGhQdclJnFt8XDIE1xU1Jxs1e1ucVArPiObhAcB/6
saOrO6E7Bqv9vVIB5SkxAQHWvN8M/f2g/X4tXqcl9RiBhIEDV7c9MF5l9uNWPmmv5h83X4hXOLiD
WOoTvFppE7RR09tD5mJ6ZLMbEuf93hoU9WMjMz+lYD8v8etjd9UyCbrEcvJBSUMH4lm18GycrrI7
6MPHorpJKYbhqidtzEZJgyg7jzN1AMf6XBlDmWaW+GoH4ClZftuvwA4VJ2LuCGpOQXwZf35s7VES
9HmnhktDcI4RXG3M1a5RMKV4sfjZPz8b3tS40r7F2/HJ3H4E+VV4HArwpI6MYNed969MbQLicrhh
wQMq5U2EIg5t6kC7vF4PoBSypsdABDUMG+poqRBp5UFEPG5U7NBbMCZOE5CGOPWaElO8esK2OjjE
z1VVsD7bt08n3hKng0fWxvg+zYZpgiNVecdachprtVIUgOg1T1HSp557+Lt4B8q3m8jdTE62Uk/Q
4+AOPY0fO/o9wUdO1Hz1T9GDNArIuegOGeko0QL/6ODAXJoVoD8QW4vETBxvt53dmhSaf13N9Q4Y
+XpqsYIWzqE1yqX8pHN9/s0GxieU+HR/i0tdNippTtIiTGtoHt4NRueDbAwbDO529KeoQni89Yv9
EzaeqTm27qVsCPnKQnHQlze5qGRsk6eftqay5wSARv+68NUF4k0AxX1qMdVDysF0VbJiFOXPt8De
icFIsjNfGY57prfO45r0dgTFmjomzGxizzlbkoJYdl8pSL1hAcGkanM3aawU2IA9Hi+dalGBn/lo
0j/lNUS1mcI0rJOCKIxxJcAp+sYPlhWEoFELqPRQ9Sj4TlgVGfz+RgXmXsxarrRg02Sa5nw6xgrw
iDPeSUnpPzMSatrnbac/O9TclVM2Rf9CnYD0+1/Y3irN4mH2BGBqa7Elq5f0DwCgyBhyRDbpur8b
dSGkf36yAiFCR/2G7KZkeWiLQoHORG2/3pXc3StkuqfXuxuqb7jwA7LBNwTRYIduB8MQGRDJ56xL
Ioa6ThYl4pviSbhN9yPzf2A+ptqMsgtLZ7kSZgsWAtGtLZtS+yut0UCN6CPRuyNnXIoue34VdV71
xxp+QwsTuML5eLcrMb7QiArgAXdW32i7uJ+Fn2Q2RUmlG1CT0gtq3WLuLmC4Ss6DQnVyY2+CvjRh
AalTPB4/fpcHWTXQkX6HY5MQuB8ZdYWSYdT7phNcFfAJAJGnQTvEZczGxVoxSMlGi4RwL5k6gO6c
pGM6S/Xp7VAj9R7Cwv24Dp60+N+Y2w5Vshwuj/Wx3lkDJihBq9uzJ+1MPQo1ntrUfvSx778i0tnX
x1B5Ew59LRvK8ARvE0SIV6tL5SDF+MMYAlapINp+nXccgGNWCA6JbGIUH+H1DwSwKjPAUFmuO8B5
zYmbiWLEoIxCpDeprfgFdE6ccRFJQU8wYstD9tp0mABhIt4pTtNCS5TuM5e6TEQnOyRn6UOMNUOH
8+JNuT+2gk3h5p9Gdp561JMRekofpnWKA4fSNgWgd6wez46PGrrpJcxQiS9ZQ6kkA6rO8msAfA33
FY7uD+OJc8agIYpGmoHL8n3wh6vPEMgBIAsVVBwq9bQ8Wr2pS9tbPX6gYZil8QIEGjToX7hLFv0x
V+tmo7H/6UiOPGA4mfOmS4k7P2xsHPUDEVgW9xowQy2iD0dz9c1lLdj0mGevhkikvNuIzTT4gcU/
vC5FKzR1nkw58foj/8vIs9dK2umivg0DcbSnnD5WMd4BAryGxbgLb2EOfKxwyDU69Ba/Nja/9PdM
xqWA1Yb9bdVyXl6/4XvsoSBDqjQ5nYSMf/FHUsOCY69vZVXhhZHMYpWKQiJ8fuPbFlSsYF/rMMjQ
8J2AJckLk4cs56X8Y/wwWYGm35T+XkwmNeYP+fX99Cmgm5vt+vFiueRE/A4SYdHHiNK/wrsPe6KN
4pL9+qcRHskC5m6iuJjSkh5smhpnJAX/cfEFAkslvWVZeAikXBjAwtmVqJPMdsNouC+/WIL7tab9
4teZqCJ3msMgZk3TjkuBA379bWYIYntFL51i+s2Z5H42GeIALlyoa5dhnc/nV/0g8sn3CW/4onqt
x0xXhalc5pLpFCR5dzIoUpfuNH0Wn+i7oSdqnBqPEz793f0cSz9JMpWtQVvp8PPQ6LIaN5RlPjns
D2L+5247kmK/7n2uYLnYBxiydfTa1ABtseFpj8whRrL2/BH63ErtFrs7nyZ6wJUmChsIv6IE8S6g
6L03TnBUFZJqREIQdBi9yoFw/CzYDNL3JQMGVr9gICWPPtA/xzFlGQNPceQi8dUlJCwzV9lRlVBo
lABFpzuwD2q2L9EncQhFip4Zm++g20iApnqnWksbGzJ9akHjsILNRGJEA9NdtN/+JY9XgupFexJo
sa7k1aAb1GQSbT2s6zrVScztofh1wlxYru4X1WpX7QBWrejQ5faBiS3cBYXbyuDSP+a5kQEcrTZB
EZFzuzpP/HGcZ5SPCn0xUDnbXdTSyi7Y/bHFI82Ot6s3CnUn+jzvCozdTMtcJtA//jIenaZO2c0I
nsnB/4tqe85qf+/fPVGB2AbN00tNWMlFwZgFb5Hk0xi9gnBMO/AUqWJreLfLbUYbltzTYs3i9fon
fGNYnRrU/hoZfzlcmd+D/INSmFA8qg2xGaIT2ARKHHKMhzIFJq/AfP3GTn6zxaq0klZQZfX14h3J
fkQKVS9ahQEfzpJviVjUcHVNkdJsVnRUkES0/cA7PHyMJX/J8YpSanxiapeyLdkUksed7H1eQqaC
Xh6ZT9ky+JodUDvjlXEFus3umgLx0ZjDM1KtAJLnjjsDM1AYjp0H+MWfgs2XxvxHGIxiY7lateJT
p8ncVGdGrZflDfsqQo00iDScoaeX4OfuUmwnUNKynuEKd5c8nH6KOtYJPGnzhpmmI08QKSjhzbJy
N0ce0jD9zKSTBCr9e29JxPPbE99qdtpOUkCiZyWwIa3ECmKLqLbAh1/olbX759sEhDw2tX+KGMWC
QZ12OFy0Nk78PDuhbqaG4NV360mJr8kJPKN3ahiDzK0c5vUlcO8H0AXR8XaBsXRrcchkn0C+kuJs
OKaavraZ+KTTERC4Z7BORzVhOXG2Q3rcCydOLumPptZa4UPuLZlTMUaAm9mQrRVA6UFlT3oYzAeI
F0SE969nykm5wbL5yQI/G8Y9gTT2D3Bcv9wDVGePp0Ahmc8Kt7wwS3G5xOPYhAbvqhZV4z4YG5Q8
nbyyq2SbvyvnuCP+yTgJXBSn98aH8Tesookpgr0sQamGwJXyR5K2aKAg61YDrAmNgHoe8V6ZfrCR
PIIatcRdrUnK3gI9t3U/cbESD0qDBThf6OyFZ1sCwhj+X764VwicCZ8lOZri/yq3v8ztLoHokzCK
wM91wtg7odhM/LzkHmjGNTj+iiLVU95jrfU0Wh8Gxs9LqYizZlGGSDqdUh8aLZk9Mb5ab//SqjvX
/MbOzAmVdJVi1g65Svgi7E+egBwwxQyCC+64HD3Jm+Jb4BJDB3EYb9K49ieGJZc16bJAZkRC1neZ
UQ/UPUAjEJP5S8bSl/2EF7U1G9Tiz1guLClwT5PXJyZ6eJ6IMQvHp+GhCTvOcBRcWTv332N7GoO4
nYT6a7LoMEbAAzWJarNu2pi2UoUiY5cDRHRCHRr70Us30QMXjBMX+m4sKg1ILL5vCptAQxfyWCk/
8rDLmis7uABEW7Exd6glKSEeIReT7/xKNMiMh8Y8mAUAFAafwcXHQvhlu/Q6JHSImVwfP0aGhzmz
+XlI3bMrBBrgL0Yh+5Qrv+ddYHUEBmDtuXsfhELiOP41hnyLIry1aViLaX5dnOGSYDWHzYZJJCuJ
VeKB2Sr/DtTXsfFTk2VmB33Cen0CaMaZ6wUVrQS5MvrvL5O8baUOfyTJIREXMYeJTZyLtIMcVMPQ
n8dX8LXNvmJoV3GFSg87cbe//axYYTj3LrMdw+pDhTaeHLjtp8IhEUj1d4gmlBcKIdUO6+vhZu3Y
wT/HZMQFo0Tj3ovuPoTDZyxI6dBc1CyxL8mvWo+iEBbwU3W2nNSVqUpvFmXCtW24DdrnkYumKN3B
eRwR/AjLzfuGnglBUn3kfT9l2/pbYQyfxbv16Yrq4kVXXce12PWfCPFXFLVV6coprgLMLQX1ToMw
DdA8ibz+DLQfV/PTsRng0gzDzuXAS86o6RMnGgWSD8y+HyfcaeloDIyhBXJsqerLEayHmOBfQMjA
BVXxQhi7LwOJL3q065dQrDr2fAsuKvrnW5wl5GJO9l1/wcln4jS1dKWsDtQX9ZTmlfSWxBzMxLG4
zpX36KVxRqic0gVqhth37XcVarWlfDYi30Gz/A0QqcBO1Qa1XH9dHPy0PdIqsDngjbHvETp8PFMg
3ii5eXPA+MixyiohYnYaL+f4VYdv5Uypl8bukzlXLzfVRn8ORn7tbRvUGaU9NuqMS05eTupvatD4
SI7uooywjylRpbGvsqjQLubNHdipQ/8/5z+dGhxhOgtA06MCdcy2ZK0w4W70CqjN4Cxev101SGlO
jj7lv1u25uvjk4SEBKuJiBndLhFuTj4e6u+waPXraRqoAZos6LcF6DUlmuQ4X+RvrM3Jf5Mr+zWr
XoDuTxaOYJTwuQZJGIXAHfZBXlVpXJASwdNy/+KrwnCwYI8/sOKrWvsFti/16E/81puhxMwN1EKo
HKH1tS9HyMNaVh8pin4WrRAJQY2Mv4/60AQkBvBuv1Pllc9VpYOSG+RD/prHJu3WZOPtVzhdYk60
pFZjWdPU8R6ypog4eGrsfqCRbbJuN4U5TGCKW/AXQymfcJEb7EZESWyoA5btZ+HUNeHvKCHriVqe
ohT+Q6GS6kVu97xD184moq7xzpm46/7ZuZr8YJjhFSkrDUhaEEU17I8YDfoVvdfJaqR2dSQnRVZO
p+RFEjCGdTRAZUPxumbQMZByxyXMONSx0vBCc/UAEAkTooJpch3C1HFh+brfp+c05jmIG/0CVhaK
CyGt2Y1s+g+ssGSs1fvjih7CBg9GVXWU+YapVghLs1mA0UeYBZsinT/hB9InEbNQBWmbAFlumMVT
l00Y1TtTjSHjjBOh9W2IQmlRt8bQSMovcHasNibic2y/077teZBCCYrSiDFoRzYkAkp1+17642KF
tfyXkAPa6uAf3wVpM+qgshb9LNWr+pdC1TBnfW2bT9j0ZGazsoKDcCNqCbWWGOq1gP86bHLZRcWT
ZOQ3os1DduVFc74x9Kp+MiSsmIrGhhguePvCfgHWkIH4dZjItjyX+Y/Mu2eEhPzP5wCYtswFSB9t
WO6lSASHbBRzmTEK7NwCx0Wqrse7k25XPkFsbccFG7LmXtWyqo/qQ2SX9gKIY0sK8LchjcvEQsGA
xTzKhdgdrUYYBu4JZ9ZfRsW82a2ZHQSjHkEfscudeBgv1r4xJpba6eOcDlSx14B+gm+5RtMAiiWc
uY1YxQWXpK6TZn9Weqbto3Y13jrEGpxwQpT/LeUUb0EKCqNvBYEP8HXMxDEswFEzEdh3v8EHhK5u
cMSa+ngayymPh6PVGVcexhEEoDptY1ug4N1czEeC6rVPskMh8JgzD5ItP394IraCUrsmFDM0slZx
PuHWXXDxsoasg5VlwGGZawFqDZi0IIdm95CroRCTE8PqJjNGKpqtcWwL7S3cXSKkusMZYyD0jM1f
rYGt2Vq8Jbw2C8A/J9F6uiJyt4mv6zYaROlVcmhjfNfYbSv4ikdA1OhwcKRSJgYMj7a5VSXlFfVE
TQwMsxYWP+RzEhU9Z0UuaorUMiqwunIUVbHJ2OCyudZ8SkYNOfyWVNO9L1CJ/EncMG39FvbKvSMz
+RU34eGIwut204cbc/p1DcaE6Px/iB0LyyZ7U9bCaZjHVO49w5T1nVmZP5TEISoen5zWMVD4yB85
D4bdnV4jhFOOBbhxYx+1GifrUfNu+JorgMgDoiVUXz18SGFdeXMWYKWt0ULaEgEME0i9kozRmwlw
h6nXt9KKAkQ9oZnZsZXAoR3ZpdRsV+/CO7E3w5AqvqcPXJmTAsUZS1o4nvQmx1ums/CZFJUoPvc4
7Pe0xbgFH/oFBM0jN2aibbVaDhbHs0jEMWP3fY0B6a4oueVVqDqXNdxW4WR7wwWTCzJf82RetfnK
O18+AyZSax5EMxOWHYp6tl96jp3b3kNgIcB32P4NXCeeABp8rvfpKaQVszKUL/5DqxGLDAYnjOoB
zJsPJLuIrT1JzSsgp0GX+4LfM3xMj4USH5DFsdBRg+pUsrfL6qOkvCKOT1LHtpPR/WhKocL/ePJv
qXeieYa9XKEreHNa5H16HAMtitDDgLeLPd6DxlaweQ39huB3OpqXyLWwX5q5QRq6qfxpgrrDYUzM
fNSA4ZmCp71BvwRtTWxiD84r+bEcaKfrCG0lelumhmHwiQ4JxtWqAZIWBCvvk453EuK/GA/Mn3hO
W6ODu0/FpWBoOs3W9pIkAkWuVdDXa2ZHd9BZA0X3S8x7UNL6X4QIIKf8AQDQuM+vivs9/lMVn2x8
7pXNbpEMM0zq3a3S3axa3W6BAdrP4V5GUEp/JRmaESCFAns1bUjFdEin03gdPn/4ZDPh/CoL2faG
M7Cep5x4rjlcJhJO7wG7XWvUKQy1NgTTGaOuBeVgDrcFErT2lDqBOyO/zIajOSTHhO910p7Uzy6J
kUdU1fjw+/AG0+2ZYyJaLtNZzc4Shr+McXMAYYnysK811FW4zbTTU69OXs2BB150u9JmMz8wONyG
sHHFYdeDFeiNxT2sSYD+W+cHzVJ9ZlM7JmmGuLHIMViPJFiffYkspnG6n1LtbCoWXHNiMOVvm1iQ
4yHAT7rtgT5Rja+i4ZjkxOpqb6WmBFmMabK2TYSSfWsVMyVf6fQbZC8g+qexmR6TYKBeun+QvwvE
iumW82NGCFffGZcE+rxRaWA60aA/jWncuqKno92oymhg6+JpLt80uZB8+qnKanghaASAcUvcmS7F
M0bcGjjRhGy5c95WQHcsKVKQ5obw7ACXw7JeQV2EAqqcURSLNoz0MTUZ0V8rEB8yvYoLEsM+BlJg
WuGfVTZ0ELc0Jf3GtXlnNYL36+RN8etG3KJm6tSUoeAo5Pw6pDlGpFlDSv3raO/XFW+idUizxWE6
52S65BZ+HBp+3q/3qpn9epNsAO+D0+7EPedW02gyRQxFnoMUj0evzjIyyron1LbgWOeG8sDZMdC/
97uwBT+yRf8bM1v5AtPONYFe7wSMYdJgPxti+rmDBm7dKqLi8nSct0D5LabwHxPeRQQmstdUTgpE
Q6jT9mFsiJXwzVLKWM2ZvQ+wK6V2k/K90ceVY07KDphbS11fVPIBvok6hWL/HDzaJVgKB0Exnl0D
9YMWhVNrTSp4NVilNHsAVunz6gH4JZQOjQktDffjorL7Gp9CVgM6N6P1yixPGPLyM14zoSoMXoB2
5KjIZD5pXTiK+OHJQQ/vtquhTqsk0s7L/61flSNzgqplC8QamVI5RNgcRTFlAIzbTDSTX4ZTCdV6
FOrqBfZp/BjvTflUHDUhfBZoZI1QuHt0DPQ6Pv5NH2v7qt6czG5A/jqtlNth/AaNSearsLw5d1v9
z5uOYEHf7rKBSCbi7h/KJN2wBFdJnDknXvFkkVw5dmcn90C9Xvdzgl2Fcqp2oBQCZKbK3MTixvJD
hWhE8hiskimh9P2uQdmFxh2xGgKzLuRMCqXlLz0GIiaJR1CvzNlvILalMqCgBfUGD3F8ab71YE1c
s+i9YMIX2uGIcixUWBwh0lTfuyyCNwY1DdAMZcu0x9149P8BnS2Gr/EpmXbZHYKedNoT8NLnx6Kw
1CtKAAitM5yWrHApHo9GTHx057t4ZqVFXQr/cbWaeqknBJy6OhUogVAd+uvs72NuxE/CiHjtpdZd
jrgtie9HfHw71qTu643Pzych7tqQ8BOzII5tSQIHOIzJfPcYm+sEOBJ6JaDuQnLO3li+I6fMaQj/
vzyY4cosJaetX7B9rJNZkKFkq0waGBkhCwMS5hYLuXVKwJ9E0EuGloJbzdzHFw+vUZ1WAyjTXEx0
xl50Jjqfhx36uKQDm0kOTfkRIudPlqpl1GzVfB2x/NHTW0K10wP8MNe1wA5quvVC7x8GgVVjcvoy
jy+MqgzfFsyx4HFG3w2UpYb3ZCluyNsgDRsstGsW53gdhEaomVwmjhtuZJ3f6sSM+h7Ynv6Iy1vD
diz6xzQE8VWfxe6pU84mCoUXTTwVQM7kGCXJ3q4AOY13IhoZFgqoYn4B4aEnIP83u1/LiKtpuhsW
Al7vChV9+bwHTWRbiW2ugBnk1w5WJBx6K2TzY7I41mU5AfHkZOfPItUKWLsHKxE9muMecjk4BVMa
CTT5PPjNZ1S3aTnZ8QzUzrs4R/3Dc/yM+S84R312tI2tRzjl2G+13tioQCOcu8ftuuovkFM2ulYQ
HA7BVDwBqa/tHuhl9f9oPwdmyCh68L3ryghde6Eowy9HBT9mt43fOViX4qqpiuSN06P0TuaASsWm
QA+NOejaKgjRVXnsmF0jCG+pRK8g44cWE6SMTWHU5lryOdPtEBhDcM1XHSGPLCgHm1/SWBHJLzVk
tfRCR+A7AswIto5IVhQ0+OqWq2E2zWdsGuON8/o/fq8DBUVLazqPdXwESZmk4++zuvjXYCWLfDGQ
ySPgLL8sftFsQtRda5z9HEpV9BZmHoM3O+BNRqXyErymCwM4VYkZnPlcGRKgGbNc3GQucMU4tIPs
9MaZFOl3lreEDfikDQ4FtnjMeTNlUmiz6dwhUPn7kSX9gXnxMVmq+XxBSqQxt27Bv12jXdCCJ8VR
vncl4Saj8fTL9tqaXV+t97gJMamqPgdsIEkMxWoUj6rQbS/vSX4WMBxJ6iBBMviXXJXvkbOOkqqq
+bKhWXsGFE37P2Ecs6ETpGCWQz0yw0nRtTHnFLiUHzQZZ8z3itfyL3vYoeFq6j6wP+p5KI+hEuwi
X4snCvmeOlASOihg4AbVNM1YNfqhOHxyQONHr9csG2jbdUs6NnRHhDgPi61zeh7qWBmQe3F/bZ1h
Nn98d5RLc+J2gZxZ1AOYUhnHnT41fEsKtGVWPRNaQyKmpWWPEj6VhmPKbYc0kTSW+QUOtqz3gxbw
Ng7EqJbSWtDBeSPrGRBby1D56/Zs902PUEsRY4Tj6en6Dfh6QXqd4bOhG1sSt1wRgGBxa86/5LA5
Q6uadzYM7QZUtfju3K7sgWSWt0Ujo1CRsADXVQA4R+T4RmFm2x/IC3T+CP870o7vv4gDIjV2xaPs
2qhTPef8nfdbfww5dI/+BgYv63DFEcRo2FwgINBeDBfJ8biz3dEGrmj8HIo45MAU6wfEhVDa5ZKw
mk8gft8tgf2XrbKEH8026/NQZDqvmERWWrLq2IVPrrJyTM2waDFjJ3hVRhk3p7gVXLHJ3Bw+rB5W
y+m5t1935RF4kxvJXmQ5tlqBqYksyuX2guHwoDZK1z4Bm9T49ikJhUjmcyz3F5phsSM6onU9/VOh
zWJrT+NSOn9PM777y06funrWZiQUgGnjtZm5wZ38mPyHpsPcKZp7t78JVLkAU43Y6bPOltbWX9aI
2CSCI1TbJk9G47Irz9t810JOqqPVgKhoeJ6uVl15lg2xRN5GL227+C085sjdG3XLfj1TMKjQofCh
7DqC2aM8Ie/8pw2uEoFHpdUJwf5kUPDg4j2Ui2TVnESDqEMRsdSdVugHmJFyVCnQY8BsE7wpSL1y
US7V8NThxSGxCC416wswAusG14H5ZWeVenHg4rXENYJcoDsTQuPIxE5xyIRJuKIf7yD6IgWzPT2Z
nJQZXgV/DykHsK+ImQPnI13tXhJx7A/05XrMfm9DvV0WAAta5gbBmcsjmzr853uW7hyb67PnorW7
haNhL2GWUybBYspfKvvx7yhCzBujOKmsjWqRZi7bq3pzviEBVuaYE9H2t04hGhBOOEj7bcCvyuHh
ZzZM4AhyirMwMddV/ooh+yoIZNlTlAxAF6xM2eyL+N4l5nG5B20Bxvyr8Xvlh9nkflNFcN6Uetwo
/GQkqc5paAKxFZDcgNP7iF7V4ky/8ZWN63NrsdLVY8E97+gjoMfsyValbO3UZ1rokb1evIBkeSOt
KlOhvpnxjT3ISBDRQNsm3/k374OLM3vt+D3jo5G1Ccr6cOn6BhtBWCYn5dilcWsc8GQX2rxyU2aE
q7xfUA58eZ8X3Bi430XRBOeEZVruvHO5L7n1LKlq+pP2kZpGeJmWZhE2369V8AfWO4to7ribPpjf
Q60LBbb8io2OQTzRYfkUDJspD/PFqwndDpCTuSPxRsPRrq3XEGsO/6hfviQ5yw+h2opLwACW0iS3
lnVz6njWDKYcGfYCTshP6IDebPHZLExMCpCaU4noKuIfiDmFJ5+9kdcKsY16yQ+XIYr8zc4eOlzv
19lYomQ6NSpEpujs4ySExDGrcdMmKLRbbMm4fgNi0sZARX3LPgX6dyTjbhzzBJ8BTQbNizC4a1gG
ojR1QxIR36jK3sRQFyLLc7i6nWmCsfTt1lZWJ/WTuYxwLojJ36K1L7AgIqjY8EHJik8ecTan3wur
VhoAm5I/cWAoIa/wanPPY9Mpm/bbzvFP0iVRxOlOUPN+xm+5v8CzKT4/lKZqeP2XdGl2Fe3MjSat
byUd8HlyBLbg2gUPnLWLJDB7Cr9wYd0IPuLr6F0Z2Z8h8YgPOHKANeQez4EPHPWQQjPJeVv9ZfdF
BbDdlkVx+Mk1zt9sb1Ef2zb8x5ezclkipISxHZWonKNBHty7J/ri0btuJo3bGRpKRb7Vpk4veQFi
BwircDAJ/eMM2lCqkteZilGTo77l3Ezbu05HOem4AROsETvFzUktWKlMFa6qePaer9grCNjgE74P
WjJkVz5pGWFfdEuuEl6wCxD2LX+sVgkR4QML4YttC7Vp75Fab8guuy1NUl5Xl1voK+LzK7Kh9kZ9
ASjiRND7W+7my6cNH+lNmgQ3RLai3LFDBVqQtSNv6ZEG3rwq0pM77QgOMuzzT4qJI8icHwovhtH5
3mRx65k6N18abxzv/OjRbXUq9S2yTq7nyMbR3o4aE0pqVebC05KaHsTFvUgh+e8dJvaGnBNcdBaO
vx2/sIu+RkHVTne4BhZl44vwS6NDr82YPtbNhj42iX7M4w6wO9z+ykKk2uZyPLl3yz1oncsKzL5G
J/YkMo6RpHjh9J5X4MXbPz4IcKn/QjEYqRa8Dm8/qsXzHEN70fLYyII/IjDuO53i8TKYehJVu0iA
T9RRjS+zRXiHDTElthnqB7KxpUxvWC6GaV7ops0KW1zZ2QtgTWVdggAyrBD83q0N6kHNj+/teBfI
dYHLF0pDbZgdAsOA8C33NCxCxD/rZIJ+s16RL5uY4j8KMvTQqXGxnkMutetCXRNXlbs1bIB9OFxF
Rgo8Y6M7RHUThGqjcH/bnrCTiuvZxh11E8b3vSgmCN4mukOuwYQ0ddwSuO1bZCU+PKEko+jmPj/s
6twXTDia8HxCpmLX91rjsj7QwbiizGPFP8rLZFqP4+YgT5uWXxb03+eNtVGcKPc0FLNKTVjCGfyY
Vd8D0NHjnuT9kJe5V2OubBjNLVE95cSg7cs4BCC9Y5Otyb84ZCO/LZy7XurhMLOTihy968WOylGA
69HvkFoi55Gn4g/4vUiptlmK1RaQp7ALZMk8SH80egn41SmGO8aBy8Vl9lzgI3unojgp6Zgv8iqs
yJiep7uqrddIuOqZlwlFycMbJ7dp0gvIWny/GpXhRwVN+eKscwlLsFTmaOnkF8AWUbjpHTxRZKH4
Kr/T1x0XwHqlNWKzxDcivTubYOA99sM2A0UV/WNLiM78E/xJLi9EBrqjt6641QF2MOnjZjBJkTqB
qQP92iuP6g/ihgexouiQtqV/vLI4WKvDIBrQp/5PaDJUDd6nioi2ZH8pqxLHLEx+M0OKSSwswHsQ
oSxc7/vMOjpfkfXVv6PCUw4pEqQl0rWllkJwKIQvIee3Y08V5aqj6xgW2M/6vCYIT9l+v/LMzpOI
Gs2uKwao+mYum1V+DvexbHiJ/tYFGbo6cOrYPx3Vl8LGsmrjGbFaQMZjcimbjqv2S0ECFBSbz9+P
Liec6gq4+dxgqNP13NPzGLRp3z+etzf0WdJ99l34HSoNGOZaM7ZdUlDW4fXPUKOtyVpNvZ23+Aa/
LqDtIu8hI9n/MZSpuFhuvOhi1Yfnr2f6WjbaKcIm44aGIY//BeI4lBktOG0BpDKK9sj2u9XnDW5L
elumMAtJ5Lan8bGN40asMivICC3VeIv9HlBraTg2uVXNh4M+Js2+9QYGP1yLzKEH9kAlmZYt4pzt
6r6Y0h/sH1wYuEuEZRHorxA+DdMt06RJtO2xI9zF0Av4fDIcvR3TZM3mBwzc2R/Ki3EgbLzQusKg
5Fkacl5LLxtif6nrtVoPOSoIRmz7CjDVmr6LAoOhlp6ptCd/lMXjhIqGxFXLrt1q4FpTO75rrQzX
txXeBm+z2Ail9Qr9pe2/fasR4ARF+v8Bvt9AZ/trbWZI/a2SL/WcPY8fEImnYJqCDPnvRx0idoYb
jLT/TjViVtkB0DwVQLkdPl0aEZsXnyzBicnTXTPklnUj7VOuMBFKqANiRJlTGL2YIs8Owi42GkNn
7LgtcpCQxuMSS3BmWxZWK72dppbQN10g48gh+vMrmrVCPZaFVrmHbBWPiJgbJDGYuwDuBqfQRNpL
C3OmdQCpk+TUPrvEA4F37etxzwH6tf6V+P9xrNWPKcTuBAmRmwi+6CBxWd6Ys7w531aiImFEfDXy
GxirtPEZX95BZMmDSC9mhWT2jqNE0zcEaqtWrbZa8wzw7ZGMYrza4UaUId1pLdTsqEwYljc/Nw0J
1GbXnAbAi+2oqFlROiW8Iy+ut2a0VJG+6UhvVXQUC2xtmAnN//ELsIcQrYKrN+RfEmOJVjR0qRDw
BZEFzBB5JpcF10RE67yvw8t8BTDI9HyrVxXhyKr/2gyCNsrkWIJNnFIG7AT7cRMVdLZae0T99SIf
1WqyT5sBqzkUZjVL8kI+b086olaiDKGMg0of5RJ2fxhw4K+MNwDG0xlcrXkGGTvn/jjhQuYwJCEp
54XHtFkJRmK4wUwdsFkGenF4UX8OMKrMKWbCRVdbOeKnYP4VJ6P01qRTDde9L8OhbM1p4icdulTJ
xR1T6A6qiJ8ICGTYt5DZ/CJRZzw++PAUIJa/lAT+vw3hbVcqUGfk+TFXif3e/u7Y+L12h3tRlwpw
1YPuE3H2pWAgISSx48sEtEft1ob1SWp09i69Rn77o/wzUlikgG5GKCaD2NZPr2wcYZHKvlQ9SnOk
mOWQqSyd/zs4i39s58Q9g6IUAo/1bEMWv8m+eWqpmeRc08E3Wrdm8Hp35SGTCBJDOZ15NM+6t9B6
7mbSJTUKZEkKtqLkaNGECNLUln2lEh7N0Oy1CpYRDR0FP1g7/Gp1raRMpkGbwQBOPmf//lazu6ei
936Ndhl5Tx/XV3COjUVLSo8FNUMrVyJBsOy6N6MlEDWmrHi0WNEjI/6GAZBzHs5AOtpEsYt7LNCQ
JRuVZCYsvK03kRFO9nPPLp6ZE9nFaVDV4AgJLIwJYic+kL9lrGYu+d7Ignr/mO8PQB52rfzFvyuu
bSNN2Omd2bDKYwODA5XyFrYxZ/6jubZx65wO5sdLUDk9Dcv3aEEKysrqi9XPDS8SL2P0i6d4tY11
qnQYfbGQ8T40KFwOWKhcJ0hxQbZ0cV27HxtDt6l3K5uELINEmDIb19b0+MilN+f69Zoj3XbvR1ib
FYXufywzhIDNjZP6RWP6hLe20EuYhjPJ0sBT1YK/9+ZWCOcVg5TCKh5HQNvRtwjHSf1l1qdfRf7W
6IlN2fuUbHpKT6D5Xhr6QIBqguwfortpqRtZjZpKkZF/pI50yZjt+HA9BKaWszSAumc9/CGuZSaH
3woWpOaMzE8fcHL+Wjwq6r9jEA1eVo0YMaS8f08RRyoRDUL3ymIccutx9vcT2fq1c7MVG29UM/hi
fCwDT4TBH1PzptmBJZud0WRt4HD0hNnvM3uI6iBQn6T4tx4epzq8n0joJY1UaU526Sh9vmor7tul
IbAP89iSmparuWNwpAHjLGz8gM1r7m52VQf7IAsyHtyiP4MIEGAyqDojvLh1+3cU78D7shNgehyi
x3yI2JQFYkgHIqyxIKcb5fm9yY1PSs1buHvusv9JrAgX798VzIJY4d7IpCU4B+6hlJU59f8DRDI1
gPtn2QDKC18zdYhhVzaE2GPF3m6qcx6CNiwdu/SAcKLjGN6nXWZm8TR9aqw2IV1fEeUrEkLUb9sq
s+HaHN8kdjvzNrhoN8UQIQfxw6uvSD52OihMwRq8MKUNSwvbkDShRoOByz+CGofRliT0r1eHMj82
He8wTd4dy23+J2m8pPJ+Rb8cULNbpVonJZQsQf2xrQGTUpdm1DPh9JlJYYjJr2wLisMbVkWhqmuh
ZSYvejuqIaTywtH5peSZFfj5UY/TWQm3sDP//lUUxOhLwg54L40GLBSKExo4BuPZxAAduFHvj2OU
Yy0wvp3V6y5Z4MW0gE4TcoObH6L3X8qV5fDVgDaAw/a3//S2O9EuD/VXkztv6OtRtB4O4QGWN3kh
5n8AVkhIe5huL2e6G2mLzupB2ajpzr9t6rXq2M+tr33u70C8Jf++LJwTLDpYVrsEZt8KM+xUrHgR
N16UKcGxNtBc346HIR5TDT8AFXxcia7z+vzdIoHdhrRbwfBR52l/56aNs6au53a8csY/LSXEwXMJ
b183QuYJ6NcZuE1+pBNoF/QyRvZtzqhE6Kw1EHYiTkUUl7p4eL8pQEZxlyaqR66VZHGsq0VIdvO4
Z6NtCBsjcYMI1VCoSm2tB57ty8j8ebJCgeFyELXmDFbCkE+8aV5UL/wQT5gKnwX/wEZpVAJSPKSR
0dp79tbMAt1bQS0VmpDeWPfFFEphPNQxbXWdVa0v7K6MNkYYN6QuN2HWNJ9UBykOS55NMXNaMCJi
PfwdH9TIqBpF7iUAC3Zs++ltIJmUXgjW2JmIYU1tk0j5lvdDSMH7v2KqsB+5MUfgHQbyDdpIZk8d
oLZ2bI8RUFtT00orB5qr5orn9zgJhwtKm+gK6pZZNd3kxDjFwbvX3ckJPbnooMAo+alCVNnYiexU
CD/s8ank0HlggyXuUhJvUxhxRzNT7JAc8iECzohT0gtQ5GdLcd99M8G29EM1w01J+csAGEgOlf1V
XwQcWF/M65TqZTM/F20putPjrBAml5d07iTs3WISY7IpAJbF9b8LSeBB5VM+ceK2wsQCFvWcNyKj
r6qRNfOe4SdXmSbXr9oEmTr+H6HRc2Zc9J2hFpH3nbepMZO6CYNj5AQjOacGphJexbK4ZWhuz359
0N9w0+EcqOT3y2piV931LyxpgirjsO14YsQNxjuma54NyjlERMRrUeeSSiEA/CTdD2qRHDUZTWFk
OamjU/C1W3R60H/yiUEyY/upSMhTh7ZiANuolw+GsSwl40Mg3Rekqpb3b7MqG14yZfzc3CC5iO93
StSTRWMIiKTSRG52AM0w87J4tB6wFpqThtxsewxzAXofRxWFeDcLZ2oFRwo55/XcWPXKWNQYGdEI
TcHvm8cpxjyK4U8cdscKnaBXI39v6OEBu7kSZkV+8aC/oOb2REgPxeYVDWgHSwUa/2a6g1CoTg/x
+9dIgxW2Imjnv4pcDgCBFAYMGLHWI6o2xpNrzxpgiCWYyNk8i6xDtXfb0hASF7WHKWiKu/cQt8WI
yRJegbBDIXW6Pk5KFZJlnr9lYU6TmeXCRH/osTSZHsxQCdmvAuWE3W8NV1rLO3itMD4EdXKWwt7+
tmstJ5WHcbIVWIMcs3HYEqKSL15IZhvuKGMdRShX7Fkjy8ETWfiLOXjC345AdZhit6xfejr4NGoV
yRzq3I343OVjRP1Urp7Q46cKgY99NcEf6bl7DEgfqOdnzaavwB2B6dW4Uszsr0ASVtX1rg1KaXkj
ZCVf4P8o91BWXZEoH32rZLF6sTnbov2mCqWsCnpCAJ/8YXgfeL++6qXSOxUSd6CFE/nQoYQrTSJS
4/Popw9GUIm6dnnssu8M1I3W3px46riM931kGMcmxu8BzG01ChrjpMhn4c/02qOv0WBAEQafwIlC
SleLUFZLxdw4MP+F1uIxMRSJgO3qa76WAEOqmQOP5W1oxV51uVSXCnIsmOX5be0HeYlteYR9DoHW
GrDe1IEoRnwt0iPL+ccePwX6j2hBxxVlQ5KWrsdBabfwA2fnSs7qAjfcim3lHcjJ0Yqeik3+hJtf
qwDB/kWEm+WOC9aNw/f2ZG35SJZs/LMBvTVrlp7lskQ3GWH/BVfJKh4FnyGAc3jktu1p3oTgE0eO
jUf/D/6PHtC1JT9J8MuvW7nzI58qcnhbsIxclZOxY126svq3gZGr6K5UzZGxCVaevGos824ewhE1
iyriEecSehw1QBxRAUHPBM0pJtZc2kUnVyUJqQhsh5V9K3gqntSLUS1bAkuCk/aoBhxmbtut+TQj
AB/G5E6Krbkcw+90Bse1ft5f14h0EZ8bya+7n6427ZUmCSiLECJNCNWtaVQZi4eeDL4T6piHZcuD
pchT8BxGxYnN1ajSU/1hiGcs5mEAji+dQnErnN3gpavLPhbNqyytvyj+xYHw1btZvDqN/o8pkDTm
uaeDwKtYm64b6Qwyv38f4CDvJqh6phVmtDeu+BHWUagS6VSeHAs271Bewkemole2KsPmBrnFlBPm
/NVEmbww54LsWPnExjPHZ0yX8OTCVIt6alhL4A/k6W7BEjDW6sLoQU80oa94yhWytHA1V2KQjxH+
4RYGFK3rheAAot2Oy7ZQw2MJHu391n3IMxEK/UrBT4WcHhEKezZdXcLwC2Eab+mzbbVkMA7AYlR9
0yC4sdVsdvMgUBF8HVc0GrA0pYOsieGaD/tCzrsMZihdMqbkgXOXZRpHsCkQ6OeFDOcAim2+oKg9
3VqJOyGui1BzbT4We7nUR2Ia1+UAIYlhYQTssFopb9CsLfUVhWA08ITRpFJonWfBqgR6LPcbZBcD
V6lL88FBV12pvpDFgjtBJVNyb6nywUQEfjUPSrDMzUng0ym/EChxs/3qE/qtwDkvULR/9uuQIiuf
sDbESS/Diht1ofrL/U3XQjjh78QX/5KQ/q7+CR3x9qrd7o0yHoqeIDc5xgRX0F58I8AChr2z8BiT
HykdbfQGzcoGyQIUTYOAEPyVpw8qh2d2WCA00Wf9O7+wWe29lW4o9e4+IQKtRnHYOc8UMOJJhQvr
3kaeqyXKYlgDIsFl0vBKCNOKuwmQurs779fta9PR7RGy9xLVUX6FgewBWCVWgVz5sib0DIdX6eL/
O2DQK59tG21aOn5LqJeERMEMlbLAp2+UkA/s7laUPPxoQjs0asvEZxdpzgzAqr2iBEojoTKTrcQj
BlfCsQtwkc9vTIV9la2G1JmKHTtf7Lb2NdKkpDETDZHIIVyE70FflVYuJ8f5lIRREM2y1ETj4LlK
XZpufZv1ixEWZNPll6TCYNaTSG+8StetZmHJj07061mTzp0JE473rSEV7jQ3G29r2EiMqsI5/GHD
+FbI7tL0+4MGbhivKxQaAtW7iVmBbNSogX0gxof4QnOu+5MYW8fTKWla/gbmf8YglcWHqxQL9VQj
LXTBSA/q/qGOSVdxpleAIaiYTu1ngIMGgdTypKNlLb7WEciV6BZFow/sYsCgv0DokUDwi5EiOX9e
dtfVOa5Pp4IHl1ZUgDhFvB8DXu4+HBZpXttW6GVUceLnJzbJ3qeZAlMfZlqubophVDQl9i5EDon6
r0MnBiqIZ8kaTKCYM5gcHGezSb0n3ZtUV6mzLqP/0TMSWk2/DHr477I7qaZwS+xornDuZidhYP7G
+4Aj6kfWZbuJLf5SuMyiBz2WhFdwyPtNHr+lrAltN84QoJcJrIPmkTPiV2LTsCuIEqnHItUtjjFn
EDqzNeNYllAWPObyuSi+a55FtyrEbiJeIgl8yU/WjBcDS7XhbnZ+bqRiM2giwOYlIHmBKEF1uyhI
ya2EY0tSaPxb4z0GaVFhxKhww3aAsEJwioDkdCcOZRp6TKRvShcxHEgiJylHzeKwjHW03eNDi6QP
5tsCHUq8449L5mPhlQQa2LoBVgesvNg+Pa1Jq/ZL/s4vpCo7wDGt836VNeHaaE5LD7RWOqJL5aNz
aDUezqzcDuK92OF3LW06pIGJUALvGHOA6Y1ZtDRYJCDKatWqpZxO0o4pwddcBb+B3D6Awl8fdzab
nVnHQ6D4plBcxipP7qK6a37ivwjIYibEiXBjDZEegBfsYQTSjBbMiiFhhV17wTZjlc9nrZ4aA5Zz
HM1aPBDfVVzMIbMedenf1o0YWRG1CpBaHD9vkPq55Iu03MhdmBHnVabMJw1z+JrOkjQsTypXsDQ6
JV4IopEVj8QtUIYacNKh4zdpLA2NV9xeCOE0lWi3TBg9Kq2ZrbwSiwQsT3eCysuAWUJojC0gAi63
IzP8EZrevqX7Q9Rm8QGrRANhGySfO0K8J/5oELM0K4UISNR/x7mhvNL5IU2J/w9DNQZjAtLv8akm
KzrVvfy9sxABWB/zsTFr4BCOepn103xlNBsAZdAu8t5YnAy6sf+ORRII85Nh5M2+z3vOn94XdHfx
6VqHPdObjNbHMjiVfL6LtKeFCuDSVW3k6mcZirxDcZ5WUHeOT99O4+tah87Z1KG2/BRudDC0d1/2
lO0QKEeOOn5MpSdHzv1hnR08GYnyu4Sgg5eJ3wjHm6FyD7AZx+yGGJ2U67Zxes/HCdvrgCmXsnTT
UvMgfKa+InFcJm9VfCtNX9LKZSenO3dr1Xmtvze75GtIhgHJtDZyEjqFV947PoQEjbE0SwjdVNsR
M3/IH1JNOWpUOvC7r+g9ez2dLLX/5k8LEMiIqCS+9LxpUrGTgZo/8JGMM1HJB8CfAdLAvXUc0ceZ
U1oDTAPY+d4SP9BV89e7jjiPKkTw9G8E72CcOKHV1YxZKDmQjp+RlAg1x9QzAGdN2J7ey92erZ92
7mFylJuHpn9paZoslvKiH8Vv44OOq0uxg8Jz9vwwuKHagZEcV7IbaPxNX5copY5N2MAyLvnTVSaS
xBYerVUj2lXjNZIo1pUDAPSAY4eqhsG3sT0zSsrvAuxNTKOiBB8QWAaBJ/WE0q0HlnafmNxusE4o
TIX7kE8ywWhaWoB92Jxd2OCdXDQkSfTxOTc9OHyEk5jgwj375o7hpNsGQbAfI0GazyScWoP60WIK
kyB6248cEdosfkZp2/aRQ6uwkjyFxK6d1z/kpwYEFg/Db5gxli3CdhqQ+zOYWnGVqFeDIq2hVVyq
cL/OBDrq3OFR8TxNcWKjx2m1C/LIjp+K5iRnZJtYXdS/xGvkNxoFU07XmlWlVCtDEVzv2OowjEL2
HPJYd6FNhQnE/gV12oN9K+1IGsKRwT1QdlIRSLXRsZYnpD51xjUrt4YPjx6LjynOZsDdOU1eAIk9
xHdBcrHUdGiHYTgxEnzpz+83JVEyO8We2p9YiQWe0eVpL/DxWLdcdndor/80V1V1nrgZ+jY2bXIj
uo/mP6vsCaXK1oB4QMPip+EtUUfumkyOazsuDvFPugv8VE7b/e03WZomtvqAiCpLgk/xgxzXJUib
CdYDJ3IRsJXDEu7X2XTxQRRs55PfIK+oQdpOWl3SJqAJ6VlrvrePuh8Z6+QgMT8/KO/UqhZYTJEE
NBF/jqE4O1j0Zh2vYl2mKx6BZLHSqfEID485bPc/r6fOOf4oz7+3+OD6BL+w3M6FPFlSD8rzn7wF
1AlZStIYrYKTx8lzW1s80SbevrRe7y55AaFGjiqci2vpaLXJHQWV0A+Ps6B+6xj+4DrHimZLv+nI
hs+RiAnDee33IjajVBvhZuw8kxPK9zNM0qGVjm9x8S0NbPEENs1RFj6OQjTvIQqwHGMeGb7/iMgp
cRd95pUYN963I5B2zUWJTtHzfMCI5BPBDHRQdNPJHyVMPyfLLERP+r9kzYhROfoWFay9JOzw88Hn
OZV3T6hJ6Emu3dS9qOzQ6xml3brwP8LmpRcksGpTh8ehudEq/zC7eVQils5QoI49w30yAgWaaedA
DJPZ5scscG0KoNsA1prdavPGhqmvVbdWFmxJ8+CGWvV2Ftq/kHWkSlFRg7ZCStYOYO4KZqPV9U3B
wD9MFwyfvgviHOmDxw1/e5JZ+2oKLBeDsNKMyfsaih2ppvQlzn0FYkc8zgfJc9w1qv04u8BeIi64
/8RuECZHnegXavJ3jRPApzSy0Udnaky4Fbcg3UOyo+U00qdkJQ79+yKBV5JNJvO4L7yg7w+1sW2s
usmmz6mK2A4cTY3p93+af81ph9guk3x87mw0flAfT8lTcNYd14lMsT7TWiCGU2Q8gFAZ/er/jjAP
2mgVh/CHDVScLodguGSNKT9rXddAxUxbbbqGYCmnMPdSvDVEDVpDMDuLc1meyGVnfzfrbOif359Q
JDW0A5qRs0Wf8nofXECyLg+NTyaRAiBj+gyUqVD17xXMHogXYS+cvFd8bL6Zrpf3lrvkmscIbbU9
YGBNpONQfFz9YZKiiTG1lEyLSy3tJnRSrsM8xquTqOSKVHV6sVlUlC+IakasR7eNil+YySryNSIt
OwSUPsJFrjE7gEQeY7MAv3sVkJel8VieWSq1FJ0Cs93fdHu30EeM0HYjqDXK048TaaHR5MVqdBrc
MNkq+ag+TTl6uX7DGXYCM1HTJyLr6KFfQoshFsI+orZEsD6MHNH6/tAyzEwqp3MVLIKOkVOahX96
0Ftcq1IWKr9V6M34kEDFyZSRHsb3o5C684uVeSa21xM3xHHXP0FOimXuhmlnpP+0znASiMYxv6Mf
oBOEc6NeLqTjHwpmTrMdo+nEV7T9jdY1AvUUjw9eI0YBL9uULtbSlUz7j7sVeNqV9RoYfwE0EHTI
xJbXjHyiSRWON1bSpVswC/3VvzKNcLgPj9S9HAlWI8ms8IEhJnOf9VUKKIuLMJf2764L+6sifFkx
ZPb8wnYJGL0FZxrfiV6cc1ukgzaMuN3if2mmyeOJXs3JqEwXUVKbSnj3DAEK35Q+i8vs4FXkYaqT
UJwKhoFSx/BiMqQHfr2+/S52tei6ayx9owBeL0f3k2SsFV0qLykq7yKi4Fx7tiYBMxhi0VXakiZH
t6WJZl0jXf70bT0ZxMw9xcTqhBwv2cAzvjcMNWcbRDTRZSHa9SZnErZud54HrWTS6o4SEHsXRsmr
OUFuIr0+UEfy5sumzp4xEYjGmGQSOk9p/RXWGfu5+MCvEYgBe1ZB8z5c9TWIs3du8yc1M8EZLLyo
Z5ZMgI/nYFBP/40D43kdue84d5aiTpW3eLcMJBotU7t1ZZUxdQNwRhyFoom9HWSF8Dk0M6xDvUFh
09dpiO0ElxD4ijU+K6/y9rhZaNIOMHC2T8gMqVUnC8qGMGE7oH3LherRl/ElGn5O0FEVKYnGwfR7
U7nYyaVdxVnVVjgndZkbNe/SPuVkuXHhtFe1DjGuCQGQlYodcW+btpWFlvne4QeuwLmEd7DIJf9I
0NlBWDUsHqVdPinpNCJKBB9uhA2K5qUBgNQzzO3/U8JJrwl1WfmAB7qK6HYhdF5ESjw0TC9UCYNC
RARfvD4L3S459cBUnV0+SKETdpwJhDlQ0C4wG63dEogc5N8wqOx8QrtARXyRzQwHBIJsunMisc7+
uCjaAbHR2FgTaFaWjupYPqJluJ4fP09w+l7lzHKoKG/NeebrOsekp2Rp6XNpuphcYHoBRNil7lvC
O6YKR0NnWQodTGqM9qBvksY7iTolqrD7IhmI30XYJRwi55l3XQXo52fuM+TBi6ej3n7whTKKN6t7
LfCiG9a5k8tCRGLXng4GpoBk2J2GTlvNxT5o5X1xgPdSRZ6kFrRVrJ2CtcXvAx2PtY3O6SoKPX4T
PCu8qy6PuQJkI2bzOzuEZR5Ye6sD2tk/8LnG7e3LN+3ElIGJPyxKtx1FqJtNoHLCAnAEBTDGrKRr
T0azIRPvEvZkVDFYt2ThI+0aVLKG8MBcSd5EL1keBCybDdXZp3LZ/6XlSkZ+auckIELz8Qs85U6t
QWhm3GRCmX+erHwqcvUCI2tpw4EnEmCKIP5/TYC+BiZg+MHU9XKZdM2kZ7iqnzCVWm+1JWi6OKg0
j8ggi7VgMfQDiQZDjNNtGW4WGU8HAOVP5Lwe3clZdAv7a1AcEHjQuajYRLy4tazdd5xOj7K/S/7H
DAOZ4756RVYni6GeFPEG2EA4yK8x9VInHHJ9Q0PBK2SWICovWRA1Q2/Gl9xqRsaxReQjgmEtSekj
I3xiwcqOZmBpvxw/v+5M28LnqrbwOi+CmaqkBqlAbzfVGqamob4AwcNa9oLWUCAQaNOBHLtNYLCZ
r7OxwlptM0Tf8WfOf7WzcfXs4e9QG+lzD9iswLQ8sXWNHjyNaxaNCbe23ds4DtKreXvoj8wwhu2Q
yTl35pyuK34aGxNv8lB5qQz9qaGXmh7CC0W7nWywaAWHEOQomeRcGfa4UohcMm+ClAfNJYFcs+PN
yToiOAX2w17ehYzUUc6+FoagmGJgIRu01fWYXjmANkEmkahH0RLlmsOE5im0alwS5ckW8Hm/FlMw
RA9c/IBprtdiMvyhI8MSLkBpJJz9G9Jw188qTB5ptilZ4Di1yWVEr8qY45Ar5YT4BvKdfOcBJnA/
BMlv6vH6aGfN2Ajgsi2CwdcsyDW/DLZUz/5jpKtyg8k95rtLiMe1XByMV/R4cC850u2FdWjoAWxp
Wm229NTu9k+miCZdrghW//LfWvqrQHUYtkFmK4J/vXrP07x4TtgkRzTUVqB+V0ZE9uNpxM8R8P1u
XevgvMlIXJ4X4eAj5y5+8IOQcmSvM+gr6jIC9qdg6ybhiYiNwCHa8/lDltw51ariLZSrmZoa0wJt
fMpEtt45MlUj0UY9jjYIkHO2UMCbFh8Op4wOH7qn9aT6L5Ed3XjRJtPRzuakEW/q8CbL95TNKLnm
KsgTDsDTok+e3/jr/fpv89nFOYlNgyp5lUk4AL4pM6JdXFlu1qv+tARzuyQ6yNcqFc6v0RuiP2ha
C0rQraBacDtdbJRN629ocg9Q68oC7Mxx5CNoyzeG4XtxkcZQkaGLRD+YBCQ4LN72Hy03f29jycYF
CVGr08rN2p9Y0RONfdcvn5OkKGTs0Ta9a/PL+gb+Aslh7GoelF6etcBx8iPhT0Fm8FSA2TxG7kA6
1Byna1CWnqA0Fwoh7gCKIk4/pgJCkGy+kroAKSHbHJWM2/Y3s0d64QayKQ1x1j48IxYZ1VMiCoOB
mq3b8WSIc5sy70X7Qe5z//lFxuQz7aStk+lsdWnebXptaMdK4iCFcAJitD9tGzusleQj+wHB5iyC
umTAyhi1IJdT0mXp9mT349OGzAy7ujoK+kRXxaEu3JudA4LGcTRlpUmLHjOD8MIsq6I33F5EgB4q
OBvxoQsqoNc27fdnQwwbTix1UR2B9/mULLXGkjD54lIA6moc3UxuN/qlWzw512E2Fo2FDzFcBOZz
ETzLB2OphVoWWFBTQffrEz1B++O+3TCUN+sqRfXJ5YZpp+8p0knZna0z93S2j81zOKlJOjjAEzse
fz85GDilh3x333N/fljk6jDXCi2MHA52D89tNSURUHnTltmMkqvkq618EOJ8QaqAoNalaQaZeN4J
nJ0Es4LyiPUC2o14lz/BaDYIAvup/Vu8NgnCtjD8sMMOVdqS7AFdrI2p9NXmvP5zWyKHYf/3Lo1G
uos7+2marXBjWAQC8B35ubKm8PC8dxz/fsjSQZKtE7Yum3w2TSEUKweSrZHo9jfB8mIEJaTADX0z
ffMusA2b2rnMS/cWT1rVBT/AgKzfuCEBc0d3QM84zsxsrVwY9ytw8OqvAbcRtkhnu1G6X6YdCIqf
kj+zBBOcisZD8DntpJzXCKrj7+11tb2FR6hz3mCKKwn2qIfx5ZC4QR5JXBbwUGj9FnkoRiYzoHgT
LXLGw/FmFuOotHZAyma6SrQ0F8vUZPld7n6zMeeunVU8HSc4dgFkToas5PPeOs8W0uvJMbOYbFPV
+H9t7T6sCYqV7SwR8nJ4p5LFDzAGHpzikGy+H3RAsnLcDPzIW9rAv24fNB/Sn8hI51efry273t51
yoYeZNmTM7t1UgdAIgaup2uWA99oxMw+dhCXMWlzYJXxpVW8QUQ4tPP4xOJfygklwbEhG74YmjiR
5gRsdEmJI8xUIY/F1NliYBl/cLaIreRvfe9kpUYp5U/xZpCRubXzJGGlDk5qFdVNzdWGi7tuKjng
omx5B2HgDybqSQ5HVCIzQ5D+572XSmpPXijqjuc+3qsHAyAMu6TZNQQiE3zhlekBWQsBpEw/8JPA
JSWjOSgpcIvX/+qENNbIY4ODItvBxDQ5vWw4j3vy1I41XneBLLRGFbBwa9wpsYakijJMvy63f+Zq
v5P15gwK+vKbL/3dZCEdmBrYuc7S83Gm1ABmi9rFX0b2LQ3asFVK9kOejEvTxTl/2skwzw6VW0OI
gEzolYxvNTMi1HMOWJRoFqIP4lby75pX68E6Hr5MWY522YD8MjwRTcL7QGwSR1S/qcNmpvZWSkYs
mT6T2GwPWjJ+qe0EbSmqwFscCxgImxL8fqmLA8Av86OUsOjmw57lIWxRCDtnAV7gfMCkqI2xLvP2
09IzL46+H+QdTCybZLjsRphfkT4pqCZU8ef7cv0rizE/K0AJtxhOVkbD2/F+31Dl5ARgop5O0mOV
TjYmHT3HMmB5W902TQEQqxyitAVUUenbiWm8huZk2256IcNebhGtU+6grpG3oG8UVUziezgqGcbe
ALHMHUyWJuPll+8UAc5yEc5ruSZHVBFHLtlsCoyh3IODaBuBWM8s39fCeIvWI4mFz/mZkPIUFu4f
HSnRlUzohtGf6HRPhUDd4kyHf12siU/gJFxPPGy/IqekaJHEgfP0kVoUdDiCSDcjHQ1rtxAsJtGH
zxb+vcw2KREKw2S8fsb+3C0Dc2ldI+vGdmaB4GVSn0bbS2nmNTOk4RAVBY4DA+xhxbQHCbIS9GUe
quNVeflPrHJYc3/VkGAA3vn/yU3t20pnZolWmQ/A1m/9BpW38iH1Wzqh0VmHL9td7C4QEc/gkyfo
kkq8ilQgK/Vsc5ToR1FdtKy+k2j3dJhfyYLaRIc7VSN/LvGQmNMNZ1H3PhNVjVzJGJBRQUXyPBs7
EReOGdbe7Z4VfE7xQQ3QRkBQhRPwvTiR5W22C15vF/OWhuHRwFC9Kt8nj9hNTjjVId6bW6lKI2mT
aqADg2WLAGne4jbi0SrH47AGETwPboJdon/p3As8XCVx9AeeK9wMy4bg4Qt71ArJf2UAOy1pLkaF
H37hz1YLkau6uiyCMmS554CWhvvef6o6lHQCnaZhnRwPvnHksmr+frxjXeHLkQHOg3u6RKflG1vS
1DcT0Sy2sbVJoJLq1kf/RXhOJksHegigomfQZWdEHWS2AcjXwAeCTVQd6HzkhJuwcTp1i2cGJeQZ
te1JkJwQw4rhZ9XUfczq2xpWxEadrHVvG/davjbjixrA8gBU45LD6IkQSFWgLHCw2OLET0L8MEOw
2x13Md65GrP5x1ZbUbKExAt0IpfLLdc3vE++TQkO25ErdPvHk6Jn4tXyY8gTg1N4ZG96MxviV6nm
VTcn3b+0rRsEB+qUj2dKp/bMED06FU3tg8Y28ZJ9IAfGgiihl1rX91FqOb6/ng6MOVtZ8kqUurtt
9hhEZnw8q9McdwdTer0knJZFV/FaA0cXhRCIPhOfRCYJAJFaYkHp5yLiCB3PuUn7cgEk7Wymi/GM
gIBhdvkiC6IUtPY3iWIuQIwQbqbnR9mOHTeZfNQlR5Gmb0ezWXBhWyMKWmay4Cg+ZvdtqbAxBqFS
D63GyItMO6mqsWON/awuhqvZZpdPX0wUnnLVLovRcXdVRyZ86Z2LeKGcUhyBl8YWvikWVOh9sJAb
DFpXJ29rUr7V0a7LfaZgDK0mz2h7LAzmJQEM1oZeH/9arYglbb+CAMic6/rEWKvykM6cGByQ4SIV
9XzWiowD1m3Q/W1FiE5q4HXngYu5FSff9zpNQ24ihHcTBau3MrpM+PGyQQW53/6F0bVYQ6pwKLwt
TpnLWAAyEjTUzU+w2D6GrdOWZwvzGVDVfmRfVHqHTQx6YDMcmF5c37AHrTXRLi6UZhLEz2VNbW4u
DzMycYTsmYQpHyQGDG/6e0eM9scwOcdzd7aQ3l0oV5QcLUXOKjsfKeEjAELI0VHHYCT4Du6Vd9Tm
CkY5BlZDjmVTmd5AzYJ2KO0Mx9RurcYL5Pged6ylhcZtr2kH14FIkc61HK0gHjCND4SAb2e3zqXl
dVGems2S2WCcqh6aFRUA+B6Z7kXlfnNmYH36B34aa4m1qxSEv1UkHP6YfI4gvFU6Vekt/7GYQ8Nq
uZz6psksv5YDNxyvfqTojfMh8kbsEFN8KxJoslGEV1i6gDCLQBBfBE977TdfjC/kwAgz8cgRAW5V
1o98Hk+1zm1SYHqPh3zlPG1OOJV2cJ22Hnqa23J3bvZTrNvlkzODxlyodvmWLOEYI9okCkiAyeR6
aJrxcS07dlT6s7iyhMVHnLEx4gR1I0e77EKs1XYmb9vUvFWBeLK59zV4DYJWTWP47lIrnbRTVih9
13Am7BPl1BMMFo+vYBSNwHcyZxTJCtdI7U76om8qXef1mHlg/J6IGjgAjoTUyLOaKH/3kAxm8b6k
VbyqFF9YwAOi2T9GEKP/QkDusgUOeok9BbNPjpMvtGSMBT9BsSvD2zofRaC09fvKFNCRlN16VtRY
fpXFAqluxe1YR2vF2ijXYkd+HzcUkbB/L3/s/EstiT+JXVaC+65c+WIpvwc0OyOPW9Ygq+MjcDmg
8qnWX+uQT2osNQh+5+NWa9Dw7G0IjWdK+YMQGpiXLaf5dwnfXng26g/q14ascGT/F+hPrTgCSglp
6AGNxTY18k7nRN9Wtkjp/T/m4tWVDB3ng3TAuo0NWEwtFpOIKpLyh/b6ZAAtj1eFu1z+eIFpjoIB
Yvug3FIKX3INtULnb6xfcHLnpMpP7dDuVF0T0dr3YDBldk+90lYjLmVJ0eHVl8GaKPZyF29DJTsG
wR8kUIgwB26lR3FYjAWSKixWjwMchdLM/1eF6wP9CBQQc2FJQum5qr/GJUVzYG4GjXoa1CPgtkiZ
dhA9o35QFhPCvnDPpx2x8e6/7/BZCE8BHcr9lTS4i7K7xCeeVaqHqQTu5rtstESijakS1n7uaCgf
xmw8k00PkrnlppHDPYDQvtdyLnXo32ctuXZmDUZb3huSm/ayy2QMCthY6cVzN2xn5NiySnuj2tdO
WYufEpwiwkKR9yjqgV4y/dfCdvNc6qXo9JFVUU0v8n1ohle1xvr29PdITp65d3bOGZARc1UAtbpT
Y8E1Plw4vxZDpg1wNu8Sy5qBSYl6W9qhaNPGf8H+PDReIpvkzEGxredLKhhHQ4kIVoJ4wXFRxHCw
SuazIq0pksspcF0BYpY05NJqwhw7tXw8L40X3a4D3BmF3Lmtu3xosFYtUjn0VdH/+W7zKsnRzqt0
1yzKW3+xFKM/1+Ym8Vn7v7c3rDvDvtyKv715FdKnCYJxBcMHU6SBelqKttD7hyw+izeRVGRzbQEY
3m8FDtAKrtHsRH9dC3gnvHMUdYFB1ITz5JbrLqu3Jai+oZOQ94nJgX7dJfSeA2rg8u9nWpi4BnjD
wRmcdrfrOoRcQexRqY/l7yRaUd4V5PE0DxzcQGei7R1GRLgFhGuHOGd5Oef4MEF5c/pxbLPFd8m6
ijO1gWm/0moP/niiucYw+hOQN54tWFbOsfhY80AyvlNkxRBbfQbZtT4gMKMz0PEp8spwldLPmLQl
hC5j6iCP8z2BBdt/wzqWky2m33sePlgKfigdVGVaOueiEjC3IpC8ODTqRZAI2d3RipM7qKthO6vW
oi4se2qmOwYCip+psuB0RH/eZ0RSwlOVnSFSpRktlHNK34Pt+ieh2m+WKc7dTJT2iSirMNHsi+Ky
lGVCxsuttbWrGTgwsyxL841SOf2u1bEQA/xdCnQesj0wmeXdAaxn541dmRMwLkIvy5YpK3PJukqp
1JzgthLQVNFzTHhytEXwlwwelKJ+teBy4HC/TnBT7qCTbcE5jyPnJh4FIKBGx+ZGMjv/6vLP7e+J
0IZok+PPmTviIjKzwoZxouGjQitcG3ccpwKQXmpYeVgbak643NqvywHtQJwCV74spJT0FCujke+M
2Mn7yIEse6Au3c2PwiCNo/anjRfWEItKF6VhoBOzp+7o/FjYdSBMFkWLe0IbjI2kvwRHhtdyzqTw
HRJYHZNCU7dF0Ns+Fhm5CsT8dDUfnznWOsWNa6fN4w7V4/orh5R+mdAXNSYfKdPA2/ioVYldoHxE
uPRZxqYxnCO+wfD9qzLtsIV9os4euiEgKY0FzqUHFAuXWJutwGHZMPQCMyFmhlCY+XJLx2SiGLmw
LBv5AmLyi9B1dXWVsgu16FHVRm81Pi01galE9ie+dqqSGUQd9T48BZtq03KgVwNkcp0TVWztbj0o
rdis3WFh94oDrzxrPyktsDOSZrkoPhbSekk15nG0i22/MsSXmd7YhPeC0Ctj7C1iwaMpOE8WoYRq
NxBubSxF37SMQruVZZkgV3w7NVobEK7WKpnov/TkSYVdxipV2TXHlJ8uX3u3L4MV8aWhStrUQo1k
sCAa0ofUyBW1lwR5XEsaRRT4Je1C8xrOM2nxHDsrJ1xfOY9S4AmKaXmPL+dbJA7/IeqwZn11IIkd
yeZvrUCmwllz7BrEQq0bfqpszlxu9yUjfXOaaJAWgMeErRpGXUETWyn73K/4wwz+xoTuGETNpPwl
z7p0ovja5tCBVuyakloQUVSMVB647uLNoHx5eGt5BPfP5qBG9ASdA4l0UPrzoeL3ZhkPf8xkpd1D
USPBedLkTGN/CZpJED3SHQtLDITxL4YikwNvF+zdWBQYqjZzry2fTBbJF+DHbcJVaOZ3rjc4qZ69
udvl0hRrGh+4Eq8KkITB1fKmRtOF7eIKJFoeYz4Lypmsxhf+DBeU7NcQc59OoUx/j5NET0rTXi4q
pSChPtv6ueSqkB3PAzJhHEt/XiXGldqpptblHUFcIkr7y/VWs53rEoyEeJLAHuLbLRvuMMNcdYFG
6tNZAwJvSCQe1i2Lun6O+3PsNgmRJnArvG2gmlgR8hZphLdQ3thtZAhHf6miEMockeEqg6xWSBIK
wimnexh01IFnJA4HiQmF1/5d5wldpT+bhrGGid+bcqOJBoZQ0N9fp1ihpSQWxhmXBF7KLq3uxTs+
Tph0LL6VfVpWWPV6QxCRt0fgOL2Y0Ye6W/enK2BkTUuLANBoINV4SAOQSvHGkisGCIf3/Y/J6IMO
8mq53clc3FSGz6AjvWZ4mSHNgkeCqgj/JyoYSycRop9VggEt0RRWf4kn2SRKrmJS8Va1nxXX8xO3
ghIYbk+HfvW4B/TI99o9gq51zjsZatzndNs8TMqMPI7Z0de4WwqphqQeAhJ04gbPvf/JiaUcsAyQ
l5iNQmB0lHrot+wfDbUw96ABWsZFuYbIFrZilMPgvrLWUmb9Oh31AIC3+gGhvO/xVopVdwbvPR5b
O3abjLssJTlzsgqsnID6pw02vfz6SEQvy5vSPhbehrQSnG426ZnwrIQv8rIATA8ZFkFzaq59zapw
mGEyjPh1uaSlHI/HKm86moPkuCJDbrr12xueWMusGIddsFq1Uo/dn0mv00r/OrolanmPvy9zaiWO
HIES+3pxOROwOZCiDEr9bJZWgbaCYrw5gHMp4T//aiCZYwwkQwu65HIBWAYNmYp55sWCXgv0m7wE
6EQQvz+Hk+60jPT8Zzj6bqCxmoi/TQcDGz9FK/inz8t8D7sddrIlqTQP4Rmbh2dy7eozVUUkuj7D
ASem/oT4U6MoAD5SfuNipynGVpqBRpHBi5V5RbUlNhvowwoXbUKa1aMKB9L088PvPzWBVxRnVSRm
wpHTdW1Vt3z4IYR1l/ma6GlEPvZXQdoajdl3n2JTaFs1w4t/acSibmEA0uuNUMPnv+O2czHAHJs0
Duz4THCaI9k6875Jom+7fyGsH5IBYt00xCJOkrlJuPkUC38mMz11neiyx+LWQOg1LuIz04JLzxkN
1CHK/KJ306syBvGeurHN10Ca6g6nG1Jjrzk5uRwfYf9jwTwAzY92KQ3wACrY3ACK0eJPoGcsDU76
xCh/pUTofICGhKYrIFTtfuoUcOCuD1gihDQPkvVTfp07i1MFweMhyxfhj6xT5kKfWm3k+2G1RbtK
aePaAFr7YoqiwcOCePJDZ2L7D3Cugl3PK1mAK8MOJX8T5Xshn0iHIHWZKyFo8qqBSnCaaZSzhYjG
HuNuompWAuB7QW08BgBi8vgzXVa01FCaFVVdRa6j/StxSxykKa9QF1pLX6yzn7V3DdOGrz2U5VRl
jfUGEhk7i6MHSCHtcKOLy/tGjTJDA6AgbH/qE1LQ14bVqJvgQZzXKXBtHbAp+vNxKJPBUiIS4/L3
ID7Sl9IcIG2zV6PCsYZiCsJg7E3ABVmukcGl8WTF6S01pgJJr5SHIaNWQtHasOCHg0oqVEuXQR9b
68Zm7o1xyEOXB1sYR4qOfSBynNgiJATBZjQsM+1uLZRznhqThnBR3KBG599vUajvjOl6eYQPMzfR
VfuLSaAa8uDwkfBCa3L9VFVXBfrpVjDtENzTQD+Rs4t9DI8edgCfA/MeILAX2+o/zSjonKpGDsW6
mVkMcNO1l7E4RLrcGiPsb0OI3AUO72rriO8mwfBT4ggj4obShMminoV7PGAaEHrIRIAEeHuMY3KO
QxTiPe3YiWIHf7ka372quwNUrweHP67ZxVlovsCZA6K3RXKjhvOUiuRxgNyW9c5c65BRUo3Jsu+T
h6WmqXsS8pb/9zpreRoPfJ9zfMIhrJGTMje2ipSmoXkOFM/Mar0f+leAEC65tYsNkhHBxSB6FMtA
pAj4rLbVYfcQohTovDkbvWSW1yuu02Cr7X0HRwGuaDLDLm/NABGfSx0djtNM0k4nvLIVw2efq8lo
fGHgN0dyj4P3sNunNBw91YsRic/Xm+n9Y8uhDP6FZ4TSMov+gT2asBNHvCpz6narBTr2QUTt1e4N
1Hr5ENl3fPLo1LWqnRZoIEW7cD1b/D7OhcZQEo4+mDvzVRYcPDF02x0+Wg//YMaPhIOEBiaAeY5E
Oh0kqKA5Yw5OBEPchahME8AzgNfR93O+w+TXeJNUcxs35sbAsV+tELZgZB3xoRIm2l9THu8fxbIb
UTz2TD9J39LQF625bhDAc16u3v9GtEjX7voh9yZkjznoLTrHEFQYxi4g2G1CALmZR4yPz2oVddPp
Z/9A9lZ2k38LZesKmR2EpMvi3yhXZthAw24qkaaHmQBMJ0juCm+Zo4ghjMrWKrA2ojo6q0SmorIr
2QBKUrhoP5/BFx3tQapiHsJ6Wqn93qREWeVfN2G8HV15VvsY3CBiE9xSVNKWX00ywL97Z/+H356Z
nc8V02IUklFhz220/kfia7qJyN9PWGJ+e7VJysVv2n8PkSCOIdsECl+5ZjGb/kfJVGs5LqJkWkPV
P7ndkmdgVcnurOBn+k5zN0YBCznG5qCFxZLXYDhGlhdFQA28omNEaCAvZLlSVFasyDMYF1mAIZ3D
OZbZ6s1xFFuhDD+67FYKFtAjfHNM74WRed3o4yJptEq6COEB1Crp00zaoF920jVERZ/z7i3bUrIm
OqzwoynYGAsqJtxH/rukCTdl3Lf2Zhttvm6ryzyeMnv6hH79r8pIH+hPYlWLoD7/gUOt/qok0i5N
qaLvp1DLh0TE9KynDEZ1Kp3hmKUc/lx/Agq2T9OC9I3+x7SingZo99TzOTTpXNkILlT/IlMhByEo
TDmWqeO425w4vCDg5UN5lwUd5M6+ld/UgxxLPnSdqEFqp3lQsMl/UC9kaY0t7da/SxFVeKowzy/M
A02AfL98hYKbFV2fUb0vrDJazmFt/OTrhCfjUGjy6h2qd5iBiH2o8BQpqJWLFFEdpbPEkRdpSoiE
Wdmr8IJQQp4+AmV2txWY5W7ZJcjU0t72dacVm3WQJzwrCbAwwNZTWZCTuQcaIV6nTWTbGOI+iQVa
HsOp7P9SrESI5RxVKTGj1WXVOhXJRPa5dGyomr5AJVgIAx2IZaXn0VLzBuqTsMf3CCVkGc20L8BJ
U5KwJpCvDlUv2vE/ZcALs3kFxwfsGiEC/E8v3L+aW8tNL+fB91yUno/37Mr91IuJMzOmkrJap97K
JHZaBzzdcuAtFVbD9tFTfV0gbInErZhFa8n8Mwhb7tpsYMyqxoi5786555O9le+KR13NlHHTVxYl
dMlxVI93Bh5SMNzelD5dddeugAV5QywvFDPh2/118+6frX77Qe+EaqxJvRYg8YZEm6eD5WQXe7dw
0CLjXIUjdgVyaZkpXc3gzLy+jLazSdyAT8bsqTkXMS15Neme9vbcoF1B0+AgGXnkpw5dmRXZbA3J
SVN/sgXj9kOnzeTkuZNv1VRoPEDQwabBqNthaVjevVkluqyXEvfSOG6rRMy8DTJMRtNmNE9+b8Dy
8wPVMouuKsMOCO1HWt8nMBOr7c8pN+mwFfQDKEJzeO+KtbeSKnIirlJ/FOQGdKWwJgwQsqSROFY+
00jJ89yn8CnC4+f3GIOi6t8wt1Hqpk7m3qNmtBZy/SJTGnn3vJRdghW0CIoHHPsExwryfA6+HnLM
Px+QPyCE2KDNXoP4J+UNlWzNR2KW6Nr4FOXI0lqQde84lfmrxThWG9N4hntF3HzLoM4IUitBrOgf
Vqvo4ZgGsJl1cIfYePBKQn40Ph4WML0XUCEP6w/ViBrFaTb5mEn4vbEwicowRvW1ia4i8x9ORRG/
wUC4Es3vYqYY2c4qduvYvlSnv55Fm/Ipo//11Klm5TbQZU7uOH4HSAsBaP95Uh5uXM9MmgrVSKE4
HNgDy5tIjePzsphQz2c1cUviNQX/uFBM2TjWwF0QPZek3m53DAj5rgKV7DFCalbbNh9V1rWlCTsn
j77ouTtQwbZID0PqNGoxIY60fAswhIsJIek8qZMCL8Ikj2uhSDk+W67MsdXli5y3DjTTpbuFC/TJ
FvgpOivYzc/jz08hdbmwRIvzIgx2ub2RSjaaY/GKKtH7KstQF4po9S17BSr1wBaTz0p5EpWWFoL7
WriVLebJ7iBwIJ1GvtJ4fbxw324unIMkEatBbutuVB16lufZ3l1ifYB/SDadUWC43/YtlELbze2n
l8Fq2dWSCjNp6usF8++BrLNnU0+75MwnvYtEVuuvbjjx5IhCNODDkfsKspx/j9dm/LM6PS5jP+sG
SMsuJKU1XHIZhr7zNfIQtYeCPPBs2hCgOPN/n9q4R6M10jJPbmy+2DVVnww+d7xfSi+rXeR3A4yT
zCwDYe+opZENQHeQy+/s0nnp51VmBQd4Z/KzcQmuEM3FiDSHSfZJdWNaFLT+YxlyIDJrJD7c2VT6
Dhn11BX1If2sjbOT6XSrvDaiFFnVmKLjo30H9JS5PiLPYdxgkPuebavrECU+ZwlGM3hf9vA+p9mv
Zsh0pXNOGY2bpbJhW1bjp3a/rkt5BlKRJoDg+QtLM4v2DZeEwlk9pLBeScVWJ1gT1Qcu6gZ1qEoI
EtuAwm5ZzY41il48AQ9nu8RusX/u6RcNOQaAt1WWnLulDTK50rHP0Nw878tJq5qsskeh7s44ubZv
zNxdt8AjZfRypSRw0Kdt1K0VhBhLitb2jScN3quov731ctQo0jWqfisINGRFIcYfBDQtxMlvAIV3
5OFcLIDv96a38TiXM21isLnvStu4POXXH1vB4HNArFIAMp3+cBjR1fZOhMUhL/8Tc7CQv9lTK6hJ
+31yQiVRLke1vpW8gXAzq36D01Yg33WIxHCv0MBHvXG+4EPR7UluAs2DbqMd8HC+le21qmVXi2sy
zJyfudM52C7g26x9SxCCIFZi2VGTeYhGslEdvNFXr+BiTXGp7xph7lpxQCq/wT/9HQ32j7ulEHR3
ktjF6kPVThW8KOc1cVd1MwLCoa8CYj8uPAE9bY7CuI9OSm090oaqsBKKCT9hCAwudyxGc1R0cRPj
K+ONRmY1TmDBRPS2EE/rEVbWoOBgrFdr3yUs/JaBgT0QiYk4OjgG84OCaX3VyPkvCgKhgMnomGb1
9KE/syQp5MGKELKUVHsvJPFFb1W2FH7FN7oHP832jR0kM0cy+lmxL+7JNSHeWXlx4yhMRN2P4yaQ
9ZKRLFLKQ5chjrTdiKF9ara6caSmXqw/XfyQBS2hihHYynTB8H3CgYNnzTJD1GjeQxO8LFFtjx1A
pCU8JwQ5MMJV118W1BmqowXSpLlX6k4MJ4dFfB6RuZKF742wBrZta4jimITEUzV5Be/WM9smOw9A
bsunX/vjYtxqb8ZiFk9+29A7tg9Ol0pHndGHOJC68tPbwvmqEyvMZNqYN2eqUqWzP+UQ3vW/LF/v
efq8ShIKxXBI+ShbXpo35JuXBhb8pQTIRap5X+g9SPRPtPzAf/F12Jj+YnOkqNCnQyVX/gWkw1n0
Thkx5GoJrUoikDRrRjBKmpvXIrsQZAFiEHf895QpyzSIRzNfseot2GwghTgPqcZe294SPQFLTeEu
asdRnegE3y07lBhE1NBRKdOHhRQpA6q96Av196RB81fgkh2FdAxHUeKFkgdnDIZ9r3M+Pu7IRBDy
mTnea0hrS4hrg8Gw6BTCEYKV1rkZ6xXcFXbrz3CgpyxAohs/XTrLb+jlhIN1UBr5MNaiHHj0nNSa
whACCqriJ+yUJG5HuB25x9B/5syRe5ltv9MIQjw2FKr7+m2ERRraqaZOMPpXQyUQXAqXeKRlFqqZ
fXsMzGnpNxQJVysS1CqX2c0OcMmrx9hWbZAH+IT3RE/CZZVES8QnuHDYgizAxt6l2WZw+FtxK/m2
+CaHsapOKx4ktdwa6dKEf1sCSzcX9MEp8FaNn/tIXwpiTqLnLkIOL9oTTrBXfK+Hl6bLDtObTkc9
hbh23y8AKQibVrFbI0AMcJaemWgsdb4nDHEp1NQ4pqmTX1ytZ0XGBGHnWfP7iWuGuTtLv2gdWHk5
fTkOeE4qqeqrxI5voxgZstI7rJIVBi1O/HEyqBJ1kgJ4gbwEGU+V5zEij1CjA0sa1W9nHc0xDmuN
fS7AGyqzTl6+R03gjFHGcQX9VeBmOYM3Xhj6n84eotq2R6Rt2sutUJl2uriaeoZ0puKGl0GkqNwq
A6aVz3GQBILOKtaErqx3TQqTnyE8P23t6zHv5Fmff9SE+9fpXewcJ4V+Jddqu7aZkWYBrwic6c+d
Iw3jWM7tltlLtLrwdmcTigHSopQNe39QQEDstTYB8VdBB0h0SiVeCC+oMBU/sQN6Cj7cgtyljPKu
rJAuJa2StaDO5WpfeRfwSZsh7tDR/yFHgrxDoK32zD5/g7NXuDSTn6vGcsnoja6BQExMGvJlEYQT
hnWBRTBlX1eF6a5982SgMPZS1WG91tp1zE49XXvZw9fFdea2iymncN6P11Xi6K1eKKlgzlVXPiQA
YVX+J6Fu7+jFTqv8k/I//Sm3dqNh9xYzJkIlgNiArnmsiJFA87QSF/wdz9nPKL1G35QeiWIKmUW3
j2/v1iGnV9gxkE7jMaY/2lBSBFw9LwM5dPG933EiVk4z97gVkM+jNRiwe0p5L19eNXv1zpm83JGA
BqWtL4UtuWKMuPNXiQ0MP61dybnO2I9e/zzgsF8JDb83huC/RJq31BI8O885C3pau3CSm2wRWQpD
UxW80sNDAcmqpV3PVzByADEhZ0jyAwq9XuFQ7X0j3XwqBv/GrbsvypOB8bnMUfdKP+zRHeesHePg
kAS8kwmyCVEFJ1eZaYlP0+k2TraVRWCFLLmPVNKwtaiU3KOCF8x1mhtbwZVuPXffMeObuGB2MVyk
poK8lt/AUIk8Ft10+E09Jc20pts1MsssmGSv7KDO+f+0MYHXL6NFATc/0Apxedqgc7lNWq0efRLK
OMbIyH7dRMHwyFo67whN+Z8vhavfxtqdzdH/TDk3xiLHFWQ5ToaQKRf7pWYhs+6kylHfk0y6r7dt
xe1/SqNabyghXFSq6woHBCwTzuLjKIA0MRB+XT6lGJLJ+tBKZw0rVV0j/m7FLLGOUZCVZzyc4qay
1qwdHi6RNiWCfR6vouEe2+JNRHSOyXP0N2XzEG4wnaTNhzUL3SnhAgudVbGzyhlIn6XXUlwyzlts
nWRibYpzA9FPmQhEv3HyjRSmGAM/d5paWmn72V+ME8j6sM4wpjggKz/pLUAAzQRjLNwyELRiczIs
C94gaUEK8wB7YmK2ceNZCSXkexOcUoZavI/i8PPyyW+5tn7hbHKihq6Plb7Udn+S/UzQ9TnqhpWQ
+DiNkH1mHFvq8jjJNVTSiLwAI3hSrdycC82zaCIdm5jIcO7ge3Po/0UDyXgLrodCuCBnPN2UDAe0
ylgbNcKYe/uralxgT9pYdjrJdQdS4Kq0QCNZQjy7NlDTKC+lpIbHM+9mvck1ulCSRz3+gzFKcBwZ
IKOHcEjNwpm/VVepw5xINqhPfYArF1DuDEfOnF4jhU5m6/WDbkdvbUduonkdirvSALq6oyXhnrGk
a0lHnnepIYG6rJO++VRDFe3fXpcN+cKfGbx3gmwNGIDUuPHlMPjWhP0UTegXTodezk0DBxMtSio1
CLyRzvYdXYxWwe0VnkrTBszVY3YHvCtb/uM7Kb4OYoxLnTwx+9BRrnsdjl3fATDykTPPcrhnD/qf
qnvuTBzG3SWwAZeoJYh19PTXhPpJL551ajefmGWfv3ADyJmTbhhQFNt5ElFl5sssDp6SbmpwLuOg
UXYOHQIJFjZ2uUmTvuYN3VvvRxNGXqrerq7sOlSzumwu6pg8ttJmh8hRffBA+aSF5aaLekTMnE2d
Mx7XUEilnVwkmR4cJwOq9NmSHWXQOY13zXb62047X26Q6IP/AkOExwbI4OtqWpT70CwvpGBhUGLl
AfKlDxFPsOGkwoGYRi7ZPQtQraykaOzryRoW/VZHBElptNlP4YSfkr83ycTkSzP166EHnxIUSJfg
8Ds4dbFXdahyp1ysaDaS3yMqhC3feegPQsvzWptqSOqY9BqnPrHqzvr6So8RE/oSN6INohfM4zzg
rZ6G90Gxap2wJxqaSb9fGFotnzHkkDjFgBlL5YKtXI5vBYVRPvhVLUuVQ/83Knlsv9uW/rscrFG9
xFC8x71y8tq9q7HyDHgZKiaGVXcQYCXSOuyKLvGYSgyiDBFNh+0vHib7pus9eL/QiaE7aucRr0my
/rh0T3IGz2Nf2cA4RZrtLTD1hid0JWEwDSXU2fYwstQSWUf9TOwWLi388xJUZRGPW2sxFVYvzTSa
/LjFE30uT5+hfe3sIGPsej2yIyabvHBjGcYK5bPPo9CJkcHotAKMw6htIo7DzZqquLrCBxLoqULJ
FQ7Pq8X6NHLYI9eG+sNumkJjAQ8cNJRc4Jsxf7/NpS3lZv7sTePtjTVG6yFgFPsi3RqwJEL8rvkH
R26C+4IBEQLo8O+gqPpIJW+REyc8ylJ9rv0lb7+ZjrkvkzAljN7W4BFLew1GujKyQb1KPlHrdIN1
6t6EY5XEAzom3MpehQlT9reaNltTP+W5iPM57E/oRnPhQo7fmig3iEHddC4yv0x98f2ciEI/vGTN
O+bNcJtYwjib8qaOJaVBvIQPio2XypQPrlkVS2ksbyFG7tA7RnPBkhxH+VjnD7WyfjSZzE4imh0b
FiCmX3KXoe0QS0+LngLlsqxS/4vJnpYKNa4H55HfG2VYbe+HjVhZ3h8I0jL2LByltel/GX+381+P
CqWI6uywdj9domPB7QtppsY6lORXTFgco0qKs1l4KVQxhqKbTJTxMaAgMOeRJTI/pWLgosAS6AKC
g1IjKp7U4xVBNegYfDx7lCqB0uSNcYe56qGqheDociNmS4MaFyhhQyLqcuClxU7BE2Y+MoBMAWvD
F0lu3mQ6GiAS2fMUZW8fDeUrynXKhC59yFd+h/X82EbDAvXF/k3OFu8YaNdATFyWXab5i8r8DdqH
vY/7Vp8Uflrg/1uEvqNGe4juzweIn/9K0Fn1EjWY1yY/+AEDIhHuEolbyJSy/IvQ6wbhWQAMajB2
abQGaZNa974rb/oEBASnA6/mUO0RB+zP/Ad5SSjff7Nwp+ekUnRXbW9LMFsqtezZ2j8tNqGUYwO9
NzkVU2MKKCMiqB9E0OHbtUvJoPiT4WWlvxDgU4q/Qso5Oyc11uqnQGNLY8gpOyixV/FANySrhoIV
F8i0lawNtjXoMqNi+rVcBbBkz7lHQCqch1eQ0GwRhPpPLhZKI6FCDqzPEglaz8f4LOs5JQHLlnGv
cWL8+hGaSP7V0XJsvTnShIGE3oaVxjGTFDuddS4azeUKPlAXd9wKRDW37u8+rN+n0ltr4W+lNK7W
N/1GH2IOifb3nwAvzIEPCifZzkR/LZcFwy7YmYOCLHlxFhWwtCMBWckcMO9SSjprcxUXE1H61/iV
rfpndw8LiQYQdO2KoHkLlsvNlljW1dUo7a7jKlcDTQ40nH6YIUxhzB6ZfyxxalrBCl4V3hEVkorX
Zto4FvS9oGdVje/xRFzO6kDqwNfK3cuzRvZ8wsuEpV0vl+M618XdsPOroxrGwq4wLf5WadGxUHkn
6AAnEz5leCT9CzUkjXiA7psxCWikMRzOTq1qIO4XB1+k6nbywmRokSbSctNYSVWrp25tmZIbW4cZ
6DWm2u6xFEI7Wco3Hz8c0cn6l71Xm6dWMhLJbJS24DfbA7NFy85pmzQkMqPn7G8p9v9eNDpKSt39
3B7dLJ4wNRrcmDwkuW7x9ibjh1mtlG9c6N1XB9en+YnzedgRZbSkQ82gzXqd+IDiHBrTqlU71bHc
q6gESa0rgXFTwPW7lVa2gar+n8a1ZNAjFfSNc6QqgderElo+OlRt/IOTkmaIe/4hTOIzSZxDeg2P
yNh8o+rBB0xZmriKH3nn3QSWGkSCtLGtqwkeeD0x6rhNW3Iknyo/k28BlrfGt/TDDiuen4EyEbMh
Iyym18UMFRKdhDYkHKf/vVhkXOLL49A30eX6l8JP6dJ+mlu95t0F+5jdDXB78Mikh5e7qvDN+8+t
hzr+bJjNPWHsmGk868DHC0zmV4OsCBbhpxNkykOO83C9TDkrVbhwJDKH8Yc/SR3vZ66OB27GYEsp
qbUXZGYdXwA0qAXPWGI4mO1UNrJvZMKcg0UUIY8K5rUTgSOHLJuk57BAxUMMJV4LISJ1dXbrPlOx
C8iaVryOzkGvXk2kV56yfmTygJ4pGiWxOzVDprCYOVqW/gkJkZFuq1o4/2QwjQb9AluVDlQiY2vr
oW6tCOLA5beY+3wqsxiTlWrYrmwS7C+PV8ejkq9NKu/yQnEFXaKmK9/WbohmRIXzB8OFWQdPuYqJ
u8KnBoOQjVgo782f8kAy9Pmylnw9ipxMCM1n3WiZY0plfrd6Fqys6iQwbqvcvOwKLXM+d5TfwoJ3
syWvrSfBTopKp1iNWxrpG2WA6x+yuGV5ytcpDgXcrQM4sF0+e1zjyAENQrcEbo6ZkAA4H3hNOWnV
nA/z4ZVi57aIadbiEWOlPIQ63I+l5W+gkuUdMxOwF+4ArLCLROLbzpFFxcStYZ1SPxA6nI6Wbsdj
/W2mclsYAVzhc/xdO0Loz6kDRwM468b4/x2kJjZuhFLbSTLikbBipxiCvxsx5kBoSSYU8MlfJ34B
el+IE2iVaX56wBetWwm3rVJmpQ6fnZhOpDmFK3QHex4D/c1fzq2R0Qr8f2T0V/y1LFazyW4aUgY/
8HY37ydZDYXtXbYiR0YyubjHR9XkXKeE88t1t7BSffYQCBwaTAW6+mF0m7sDci22I5a/9Is8tEbQ
aILWjfHSldtj+NyYD6mEW/p+8voUy9xRb5avsmdM/LzLtdI+pKDB78KzzJqbzuPso1sQHs0nUg0M
1HghadIu6Lo4tKauoVSGLemQYPd0xOGqHKbewPdxnTTz2juAOJoWKj2NPZhCA3mA7///iKrYkp43
psmyoYFwju6jToNY8Sdglo3tl5z9AggG3bn5AiEgvL/+ExHVHyOSL+7ahnFFzn7ZeGpb6ot4n2Ew
+QKnfSNtheM7yluPUbYlkp1ydl65rXrhnU/dJYOecECM/or4K+isI/1BDXNXQoW9+lrphEvuGTy1
D049VYLHxjEFkDgsX50gUU1QhkK8s9omjLFNiNqvvZPwB1SPqbP9IhVCj3/gjMftd9XimrYykkx9
WVX404ygsCFDFX1H0HLehdoONs9xAE73Nx3BFcRy5Q4NGjiUTfsB++6B7e47NFmbcA8K844oDu7F
ya84x/xJRv7yfxxQoM4AiPWzwCdEeHWwFoXSM6zhQiNs/TbFqrAV52g2MIZMXj145xs0o0uNo2JF
zOcGp1Zi6a4A9HsdfmF+2nJ+OOdUqnmhAB7p0uMWH+VPg16ILYfhrXzLRrnxoM5GkdqzivuYhMcP
g7tV+JfNn7PzMQtrpoPIbvD6fgfh1xaWzqRheP34OtyGXbciiu/c/JY3ToLbQKADcX2LH1uWoPLy
OEYwMjGsh/JsIJdyLLLYsa4Fu/2AQnycy1no+4wKyTBDfY19E6fjExEA2uk8TykRm9Q1z7nDeWbQ
unLn4M0UU8dm1LEbrdBvlwqAqc7zaEbPiiFCiknLnzPICHeYCJ5cp6j7fEiuGtnGLKeo/lQSzlQG
NlOVfNdLknQf+iC0N9J/Do8l/u3eHGttAxtMNM5vnoncBRDRDkTgn/1B+y9Oi6ixkYSrNSwqvW1j
R3fKa6QtufDWTMxtAe8x7/8a3M02+auRrMyHuYsjQt84d5rNWcvN/BUs6U+jCbIPg1McRtMeTnq3
n6sAXbRFPnzNebu87CB5kJIN294AcRzv7GG+xmp9Amer7Mk1K0VLdkn1e1+6gbJujzJHRhGgbe/k
LLjWioB/AC3nwiAWW9+zfv6yRzpYenzqM4+CZwBgf868RVGHrw+SAQGFN7AjBcgynbeED+3kShNm
PZe9aGuJWnLdvrZoasoNxYM8ZN/VJ6LT2dcCQA+qTJqdUj6tKT/SmkOqtxoAlCCjY8Uia8EyluLa
Xj4Akeaia2v0Ee4dh+Z1yixKJfRPIJKO/0bMSAE1UTAgowePsXePjWHtwPDKAPtNK7oOfZq0Xsiv
D+/iAP8g9lf21uvLCP2GSOvAeyuLoca/aicWZEzAcXiKu+JNVTUElFsv9LESWVli6T2fpEYfQkul
fy4/ldOoy8PjNvEGxF3A8VgG2ZFY9v1P97uwqhlR8Ugh4eYW2h7aXegZDuoj4zDwZ0I6udipMBtO
wmZON6Hk7CfR1WDXyh3SiBg2g6ZI0ghnkmdBRhtMs8vrle3jZEj0ThotxZET8aAKgqfITdg0AT6H
wWcFF2xwLkSXW/6nFjde4mX54O51CGyFKN0uPqA/ClGL5JJpq6/UMSsUC9Zvrwe6TPFUDYAUVmyd
zOivIBH3NrfliEGUqMFTgkXLzbPfhueWKuu1ds0c+VBn7nVagjOlRSTJD3LEwyFJ8O1i4hVEkbuo
N3/Sb1/jooXTUm/uNu4E8UE92q7wIOF4kimsJJcYuDYB2JLOaWFdNlg+DAgOP1Tgc7nu5EPBk26j
MS7MRXsL+97fAxiXIkloZaWYv32TfgFEGM6oM8cqCgvO5kpWPDP+BrVrdRFHBLWzFDtZoIciqoi7
1yUxwZpSQAXt4yfXJBaU8dP7JdI5j6kBda8h1in1lfof+8BAICddyW2AIAfzg6hfidwcZ8uOKV0e
dR41dfOfKIFSa/qS9ktha03LoSlzpb92wW3ThcRASDgSb5+H1nc8LdAQpqFny/SZLugvHh+3O3Q7
9SqW26/3coTrBTAS3f/8XaRqCbydCP4TXB7D5KYodSBAfy5YgjA6/pUQ69llksLgWXhQ2kqAt29f
8NvJ3hiSl9GFBcQBS+5mY/S5Dc6Yh1V7cWZH+5LIk3Gc2E8ProeQ780OhrwPnVHQk/ySUoPXM2rE
F/MoSnArB9nkz1xg7xAPrbz+7k7m1PN3pKPNKAkTGyt7NGjBjb31BLqHKUHSdH3B1mS0RkWEPII/
FVDyIl1Wedyuo1jLHSlnHHfDE2UXfslJwYv1Q16fH66XA9MtjQ7Tk/1CAVjIbLR+mym+4WmM2y60
wP7ON9Tx7/SO6HDtkLe24hkWZofskrUOycWiUWrkEdEHcbFKbeGIhyLO6LIkSQWo1DncOwJlUWrj
fSM8BJ9FEgx8ZdFLaO0NNjcKz0fZZkU9FJQW3nDTvov6FJEkSD8nC8cju5s/LsNypc3FcGA1VIS0
fdpDnRPyKMTeFjvups4z5mvIL7PkPUen1WYz2nGaP9P5YHzbmHOgkc8sgssoQBhGfMXAiIHMKUVd
7Q+EBUIUVmKQu74fKtudlTrDmRhvG59Xc7rW1ZXB3sq6rqQZbV86KZo29NaW1JbifUUPUNMTPCrh
7JQYY7JbL+hFDsfabg+mx0ocG/GQ9zGNFwBY6zIYVi2rlJhCv35/kB80URjtkpGom4zPQt3pOMzG
I3bc2q8pBpit1U9CENgRBTdh4JWLkCxA+8Pvzdd4Ic/gzetw3hMoM0vI47ZcjanYYSkC7qTIrFZ6
1CTp9NKFaMvn5JTNtNomMW+UAGIpZzhsqgoyKZ2cl1AsZssWsAcF9mzJrREJNJnzPXViN3MQUYII
W4QZ0Rl2T639ryL6sN/cYN1aboFAO4RAtE/QdkQOCJtVU/p+cPEdni+Nw5xPfBjIV0OR7R8QlYEI
295SqlOMQBh11r1bM1cF8DrC31oPCdVqrMsPIX4nThs1RuZSO3B2y5E8KF83p0oOH+X98jiK8z/V
m4OVDrn/O7aXuaYLGdz4EkS+m1cVufLkBsbvaDYRgryCiuvM7g7n5vT1mjgv9U8xOqtX5g84pXSl
JjHlGVaMA3lmDyLP2uGQoFOKp58sfts/ko67lsqcd+b9k2tR0XF1APQyP3C6YKD/3U/gk0kh27cs
69tSy5OG1Fwlge36Lo47piC2x0mHhkS+bjxX/UXKLTilxc8sxs5xGfvMFV67fBWANia+4Gfdyx6F
nbPbjzeCI9S7qgzb6UXPhliEJ4rVkIcZGpb33GVNpy1sFwEqV/kMEQLgDpPAoFU1CmJx35MuHXNE
NBt1lX32t7cyEOfDCk5vbidPWXzWmEJXo6T+xEdUSiJ4RENnHt67j7xYDIAOCRtbNTu0drT/oEF5
6WTY0hz/a5YtBUKuC+gQ/e4KMlR5mmXA69PivIYvlT9jyrPDu9okZLnhzS4CnAmk6H8VgBRkYJRf
DloiZQsaxjGTjyR1voi1rcE+ft+7ilKVDYojXYPyh1RN8lCNJD41257aM/evtoQIgdkjeXA9gM3U
Jrvc5aeEs8n0cejcLUmVmhWhSfuJumZdd8i+oZpySguCjl5YxeRoByDoEJjknnwOazDL+YLpeSo6
bgXewAb3SULL6ao0xY19llXtt8OQI2vuPYHbeMxAHTYiWXWvueaLgJN6UtitHKBtVTKNiOAZMlrK
N75Nl1a8RIcb3gA+cSMYbU7Y2qU+AYNG/WB/WrmT9mT+yBHaJagDK1tS3MBES/aSxE/H72o6X5mc
GJv8JX91MAzv8Zg5Z2jvIY581BU/Tu4EEtnGl9yN3gBPh72xb3nd4JR12cdKWXzo18Ih9tkdUiac
tEpC1ukOtiUpahjcAozwe+0xLJnYM02kRJb3Lecniubs+TI4Aj1/WcQ3N0fHigtBxrC5//oNOkmT
bZnHfSpG0dQk+m5VCL18p2f7ZR8UftTb71inI3EoJ+30316XOOewbhY2MyGQsXVjSlMGpIMtT/Hs
u+6/9bVMa/dojoY6K5lKCZ97cTBPiIUghaiR+/7PPk5MOaO3oKJKHhIK94Xsw3pOtm79rVVItd7u
RhTnGTtau7hE/3t8aMx4yFCSq2PwK7YMY6Q12auVA3fozADln40NZBe3W8+IdtSjHD7Y9rw6x63z
zXeKmjOpaHWTAZxbyAYEdhoDWLihrtnY4+R5BY17ysXRneT+XQuq10KZtwrBlQ+XXG+E+sVazxd9
MPnKsVlkm95C1LJDoFZJQZ3axEAtweZpMwp1uMDtRl98i8nIe0ujf3aqV4czpHuJm7UjQX6ZZ5XQ
ozdh4NWjZhtL8kTsQ23Vd9PtOPwNLz/cA4d4RPAPEd+BHW+v8l16WVbLSLDgJ06SDCpnSCrqjr4D
qu9AtPPngvQvQ/ehzsNCjoBz8xI7Mo0TpP0eZgh92PTQ1K9P5jM+4A/61hBILDoR/Pyv6JSfAuHV
eCitNp9KRwrvReVLnOV9ajX5dCSuRfq7qOj/bByD+4cOzz0KpsKbQHRUcJrf52rzDD+gVNNUL+HP
9+gYBjjBkBr8RC17nytXsB2VxMqlfdflYdG5Skl8wmGoufBWosxtd+LK6odTRmcgUDrHJ0XPAecc
/8ZhSQuMGWLQMeYHNutasGYgCI8uC51ao0/q6R16jxDb5WyH5M0gTRAmVSzxl9CYMJIX85ROJjvT
D8X6xpal1b7Tv3ZAxLc0RAB2R0+pw/0b69WOo26rmBz8YM/HcBSpbyOSg441MOy2/H7gJwRU/eVL
jw324htMsnZdJ7tpVSxipPPtU3xATYhWisRv8MXeuiyv+YZoRZv8S7pACYvyAKW2JSWvv1tDhyzn
e2EBYTZseI+afhrr+2HFv2PKT1YEOSb/ZGsb6h+njmOaPleDuGxkPrMRKwcm16dA1Bp/lFRt05Fg
MjlYIBGCtTaAkPe0PvvZgGbUtTo1xLhIj7zRzjldaPZQB27rymNmAMqULVfHOlBYlVmcAjKC6xtr
qbp88V7E3l91uNSAO3DRIDppKW4xAh5P56Olt/o7vJEYK++8a5d+atHX1yF4/vvYpRHL/P6Ye+4M
LjIl0WeKGFGHMWnNraqRg8Cx6gLAiAHusnF94VzrJBYtHo44O/BH99U0G/d1wC8rn3CUHJyCuU1Z
9xuD/eLPzuKNz4rYr0ldvUoL+I5kFfhBk1RmlzjWp5XO/6CTe951OxrEwM7ZGMdf/UOrmfWGh+cO
OeG5xNcjt+RCG6R6iioZEYcSO1QzODMaACHcN+/T4nVL9j4pzTB3sYLNm4AcIpndJ2cboxTmRtQh
vNy49kzSFPNleacr2GNWfQ/LpquavIRPNnXCdKr6qy3AJZAPSeYCWuI+VZAansYrAzKElucDJPoR
83PT/cuio+PzmoGJaCSuA9un/RJk2WaNWycMDL1lVaVNJsWIlJVD1xc8G/prfO2fHNMuSylJE6F5
5B2x+FbfdnkbLIzLNUnmZsbjNaq21Wj9sMpI5o3iLeK1CpEa1f+ggJZzZ35qzT06lvpwak7Zwxtx
kq3RhVgnLL94/ZzFn/igjPWPADSI0/kYLwx4xFkI7MX4W7V5piphXaiv284biXJ+PFXCfFZVGmNG
5o2Dx2lcnsybr/1LlHAx42rLCkGbnpg02soZEYQ5EP0dFxld9UwiX6dbr+Eetk5JtK3M9na91Xb5
nwSTcXJXHTF5osTwREyqHfTQUMe3aNByYu4efGs6oWpOPUrjhhyncn1toLdDUzXFRw4H/pUJQ/gh
OMfvv5TrsvD4WkCWHKtSou2Asr1oI60SuDgH4M/c0ZPAOY1aGot3VyFfR8lZPBRWR0eC77naiYWF
8i11XHyQTezdqN/sD7nj2P4IIfoeV/C0MeNNX0APoEeSu9w/+KRg22Caz4jNIqo6yZeR8RYpN9xa
PjUHISLfRWV+R2dpsDecLmvhMr4okoJ0GAgQQk2njQySK+5UosfHLu0Szxly+UCemeLGYLXkeGC3
96H1JvKYsc0JGZ2/Yi0V7JIqFaoA/KJGWZQ+I8hlQOT9+xcgdM5L313JMxgnL/P5CtTTrLMrXrk9
kUzUNJQfkntzIGU0HLDqMx0QtVv7ZjV0ePav4Z8bOG6RNhOu+jjIj5Xla8VhGweTcq0XYH1A1Im7
7NmNQkLnDhWad2d0lyyNLBKFM3l08nSpdGIJ/QQ++3EbnPK+2QbGUN7VU15hmkhQFXR8qVwQqmnT
xJyDXPbM5qzIvcUTUms8Qj7/+G2HOahO+hSM1VrN3oOtHp3SvNWQj1D0XMx7jqgOpoQgqkgkcemj
1QaAwGNqiyspUZLky281aKTHM34O4jE9uWzIF5P//c5lnuEUeMlwT7+3tUEhTiUP0DYJemziqf/Z
VZx7eNeSBUEDkRtOL5q3FBtyaUyGLPp7QG5sc20PtJaR6dGUTUibIMwUgxVmHCVHOK8FlzRLJQ7P
otT6MV194fe3CFbfAcayj4cZoq6drRjSM9M82Qta337WLF01/sz0HaA7vaqNz9ALedAxa2ef5ujz
iPUE27bopwPNf6tv/AiY6rDfyHjTF64xJH/NUMepF/oeVHD9mPqb+sTLLi6kdzMi8TP4zecSDiEI
+7cGNJ+epe4MA5wyYq9Th1aH4G8D4PP2hyc+3t13aSKTQrZGLOurAlwHRNCjsIOhCjGqajdiC8KO
sIZtFoLi2SsQo3rlIt0yWvYAFsZGVjJL6VQGdnEq7i5FfxHTT3nTdc+o+SG8ljWddwdsM4nOUw0t
R+nTQmTqg8V8lka6UZYmfNkdhLnmCSTBmNKt1j6F9syd0p/VTmkjG8OfvF4y/DL0afixVmvfrQTe
w3Wxs40/Wc+RQiwERN+yWYWrJYsN5f8sQPoViCD3BMil8NBVetNBzdeDqShn72SWFeS9b3Mgwx9x
sIwr+7xoiZRueTKp+R9sHD/ZuQbsOoBiEIjYf0sHuoCRWrYbxrFIAmvre45sT380Zr2Xi8OdBAg7
DqMjB1fgiFwW6Q/F+CfkK3VZ73RfdPwOQOwP2ellyDtboRZTQNmSxc+An+OopH7dfoTubx0nSSbk
GWNAhYKWACSlF4wYj0N7MnW9BCn/JhlZDvSV35hhc0CiP1hBBcU+8rn3zL5XqYdSZq6nm2ivTd0B
+I45Eag+MyGShPas22FJLcktHuiIGl9w0M+/Pcc+zfVOV9eBQlEF9+Lb1FJZ2kWQDdyayYQE8l29
9o/MumEiIMU8x/fNP5Fflk0v1iLm+0ZKtlO+1z0wgepybSPnkfnY2yT3fIUwj3B+MpJONqagzaQR
fTCZsOWaW6sMjsWhPz32YTF6NEp2Nq0nK7tYizfSQrBDjWOsJd42gWrEd3rB3wNvG+GhyR01vbKT
uQIAx/kEi7QXzWokVVgYGPwf775GTFy5sos3xYGhKFLMmVSL9IJq8AJgXJytshb2+cdjhp63nVbW
JQxBjA9S3azKtvHX/g6w+JwybMCFrsaUKAuznsvSZ33DUFkwee8yZJyYruoc5p8fzlwM2ke0cU79
FImjFNC+07ua/u7XFS2pEPifn7eN+U4nooitzHMNqg2vpPrWKpPY+B15TyDwn8fbuRcVqlNwUkNY
tzYIbVBjuS49QgC7COdE4mW7yGy+uL+76Db7T6cloG/TRiQUF5lwrHrm21ex0ulOtpKPWX3Q99YU
tUxL66K6uwaMoZSUnc8DBkIw8ca/3NNCu5bOYT3FGOE9iQEE5tYjtno3h1XUHy7Vv3s/DdImMa5D
pvlp/Ap9e1NP4o5BwI0vmPMHJ49Pf9mTFG+kzmgELWvxnU4rSmZiysrKxR3iKbuH3dx4FZeQ3Q+O
9tsXhLL/HuhqX1SZ3xyfE62DHzP4eoBEP+kyrMIjff1x24u/LdSk9DO3wPoKo38sCZdH+uReEwkO
9MFjmNO+bxha8zOUFVOWvsjrnaO5TxGr9CWeeIirWS/2Yqzf7Vl2CsuQd6bq7jfeZsFTqRmCWCmm
5W9XDAsUtF9xLBA3XZJP6wbnGlq8KiubP/30WPTOJJ8WJHvOeSR8pKXwkfxKk45uCE+0AiE+XFYY
mpepessUXVRqhks2yni9cjuke4BnKmgtzz7gjW+fzGUmvYB7IhkHQG+3gb82o7lbFQmxzsSYg9o2
BAdARlHRxuVdUbVBM4qD27dAYufv1nEv/FCo2rspTG7jiRk4TsTBVJ1kpyIfOUAcg7Ak1T3rtUzY
9wisEg40VwOzSaiQ829O2YX2jHPJNwKV+RJCLFQACUB2v9n1uln9JdF0JkFgpwQrslt52lJsPIbt
hYszKnoQBL18F7hg+qt+RmOhwuZNpjAkCCWDjpLzYeBo1hRnGVDbAXGfZwvOAhvI1oV33Mr6mumV
TbRF6TbbRaZI4dShideCJT9wCTVaCeStmNhxugfqDoX4mGBJ7P/lghFHXJf3F/2UOTwNbQNVI91F
ckDbp0RsUAepSZ5ao6htixFSrrWndn2JBfTdthUuG6GwlgbeYN/KqnVsi6G//wf/nr9paXTuVZ4L
9T5+7k1mnV5sceWlAHHZHjG5hxix11D31293zJPMxGpu2QpUjJOhc+d/wn/u5GZMw8KqBMo4wc6d
84fpzyM4XhtMZh1rEPoq8Ak3jnuMpkJjqviluXn5geVAZajjTqG4l1DBqCZiNhRZ95bq2kgKcYEQ
DTAjFGxAwTXjgZ9eAN9U9kadRrqu0cP4KVKYAoDsZno8nTokyeBCIf7/cQ60Ca+xJuLsyBSL0HUx
kazP2Y7rW7ulZB1vtAdAmGEtffQTgtEe1dLmc9mvWNP6Ds1fuhJVflwketlERik85+nbSUn99EBJ
iRAWmYLnrBVX1EFjlvqxKP+pg/ZGPmAm06DFiI32ZARPYdWNAhfYvG+OJ0oN5eAGoOwJ2glqHgrJ
iIyMRXe7IaLkC0/ndvUqlq/6F+VDYgVRUStjUfOWJICpvpOkiF8eN9ZK+1XpvtviZM9oP54HT3ni
SZhfj6yx+jCGSzYyAMIltdkKSFILfq7guxp4Eme7EdQMTYX9l+Tw8Ft24O/iWoDLRUNBFXYsz+Fv
9G4WTdvtEZRXd83MKk+9+UcwdC51Cu8/IRkosgJ8jDInikPwu5GgSi51hD0PfI/SBBYylA8GsIdp
BKy1h5XVTIe5V3Fhy0YY/atxSd+tMWMESl56Wq0ZTPrOHZ6tVbzR+e4BrkjP7qPDtDmDxJILRHHQ
U0zbWdsQeo87ljfYBy9+Qjs19MgVOD3Nvf5CjOV8nHk72UvKfyCuBs78m1cx+0itEIhEOb3ooEDR
Pu4ce6hr5GmVnTKUh/hyw7uVL4SZVCyXDf+uUCl7u2NXxJG2cwARN6DrIw5t0tNdVJihBV5PcqVI
Kkzj6Y2PK40REUS0ZHUO9nfkK/oH5LhUCJZYflUsFoqt/MVNNA+0PdDoTpsXMlQEDDh/fKPK/bNN
NOFa1CfHqRGdcAaWaKqwBQ85Q0XkKDeJs0tJ4c9Yn7sAVmygyFaHrIVWWZUA9FZv5ZnvFcrdjb5D
yjkhJket0jrJ11Ik3GejFecYlQeFsL3AwZmLc0sbkPvMTTCoxES15gKBmp0Y52sQj+GfD73FrYdz
GryCt07NIikNpwSzLVMvnmfTWwtu44Zz2py84XrOdmhswcTSqQ2vslkvNTLOutxS5LhoyHakiMKG
Kd6Fst7Rpu4OVadeIHHFqN2Xunh2kzZFXQCWAwp5GwGnNJqxtLHdzXDLf5U31JB/EDgc8whdgXCH
VXu2aggGr0eynWzsYMizHODpRty8osGi0hsjwfS2PurqzBmnr88S8c3FP20X2VK9GCL++qw37gsm
ys+5YUzW4jCsX2+8tn6HgYXPXJxZRJz3naz18XxnnyIWXgrbqHYo4Tn4Yw+Z45OhRbp7/9jezBUB
m8Y4RSJOFXSnRMiXbTP43/TQzz9AMZjfa3lAD1QiXvLwRrWpsm4ggVe33p/VAH2bKG/VjeJnM2dK
QHtuwuNDgCu/Rq885O2w5aAOow4hf0fCVSLKHi4B5HiMwkOJMVi22pMa00N6KqusowxcJh/ykGZl
b0Z+SX5kFLcDYJbv2ECaWzr/CbWRCfNColhSW4DC3oXocQMzWsoKqHAfNiQh7CWkzZBsP5mYKM9j
aQ4dm6w4mKM90R0oqs+ps9SLWsUK0N3hrKnNDgHjcf08bSuJq9HJZBMlw2VYy1k2FVF3utsFnRL7
xSzPP0e3DzI/WMaKzsq3uzBAD+jH1h88REY+04koJg21AJmYPBNmzF5VkndrFLUYsvX81jkL4BRB
4xYocQPPXDuw7My2ts3HvU7OUu9WXNBfgAwkTt2O1Ss1QIbQiFyMzWbditslq8byyF2lasUCEIG1
jKeRYtNSHnRGuahWl0kK62asTwgK+vmYiav7kgRpH3GZS2oTX9F6oo0X+LFZ0RWyYCYhcrXX5XhT
CNfhENA9gZvDWr70qV7SEfUN85W1vPh9EjjDGAqx+ZONenchHka2P2g2Fxsid6GcFEmRl1D+Kp/d
+KFxP+mP65ephTL/lHTCzp1R65flS767R2qFUlSY3NZqF07G2SX/XQJ30EXIU9TCJTvYz8BcYwon
8yXfMv1yGVrIHXk0QBbJ5v6+0iZECjWiYtQG5LQ51NGWJhUMf2JUGFfOJH+O7rYLpq78io1WI406
H3d9gNghfqXh103FHlwPnQ9JBQixEtM78+3tpUfkkakaau3E/WMLT74qhvJnupHnje3PNwj6zqw0
MxgeoQyZsoLHArsZuc83yrBr+JC33JacXC9wLErTYzjGc1blT3FFoD/JBiCA4tctimKhMlREYqF+
xODFFHY/Gz4gLcJX+QtAcTORxEnNkDrYJQGiXb4CnSPujWKRrLaBuu7xik+W48mJ7LKy5DPNA6Nb
cFp14SNCp8tnN9gyvrmPus8/DCtLjy582oMQSOVeY6kD3vy7XcQircFa5myEnHPY2at25b3WnMpy
1dEc7nYtNzDEt40u9musrqbacxJ1QWMbVYrnYkmAg7IqhCYRnZIr8SeHfQzkhJkGXLk+Xhk69yaz
1ZmRBPculLeAQWFw2sm9ev957oOPNTWDxjm5qT5FkTFlVlFIO6+g13wV782OMDKFAuewv0M3K3Ww
lO7yUgZZLzmZzTyAFxWrd+q/PPSXn62y1q2vw+iK6w8SlDWQuFBBtpsYxdiIrCEPjTB9aO2t3KsK
XiO93igr4yGRJwWeWTcolB/n+kHCYmy7iYqbBuZjEWwdRFmNEcLOmWISfgA/47zvbZf1fY25qRQm
yPp8vOKg6SIihBwXxDFIuGE2tYVJLnPcsInLUJegF0QZoOelpGHsNmaquOWQdibfMsDOV97H480o
frONrHIwn7Nzx0nlrRaNDtxW4OAkvv9hlG9Tsnz53M+3aiWOL2Hr/70DePD7zZuYAxz/kb3imscE
2iN/cbCALRNqfiXA23WF49+8cz0cyO3ZzroOGT7IMOLVuUPMvizh0q+Jt03nalrMP47Ujhw8tt1y
PkhsJeDi4o7h5H4M413e6uXMhyyWEY/O1NZGirEtaZRDbeT0FFjRAPdoAGAolKFfii4g/F9Kec7C
Uk+hBRVHonh1z70R9WAhOI+QQoZ+H7xSKExM7EWFAqYde8JlSkPP8s4GGbDO/rgdXXwgJjnn3Rq8
IdIAP9PBRs5eauBEnQFhFPabp4ABLv+CJGjWWp4VpLu5++V6LxKc5gpFQIoOnDfeiGtOKmN5EUH8
ChBnlA3KF3sSz94sWbLuhmUkaOCB7BEpHb7WBLdT9Z83LAqFoLPk6Tr32CSYVrVqU6yW3fZiTUHD
DPUA4MqWbh6B8JJc1JS/qyc1YDBSgFlRQUdw6HRliUI0DdR68ryachdOlN09gU7IBsQoA8qDF+kF
X0YYKTr8OpUqZVSa5diQsuh4YuQJI57Acw67adtXNjQJYaC8d2Kn0J6xFRBH2OhX6bIVvCHh9YZl
9aotquAbkIV7BCbdxx7KmYilg3n/o9q80CL+A5feYq25OD62H9BhugkwKL53pd2eTsqGbuky58W3
PJukySPg8PmN5h7H/SEoDKQe2dqFBy6B8nct3k5hCkKS8Pe8R1Fl19slJUxMe6UH6wjxXH57gaUr
eHUQZ/cLTw9NukRdvUGgQA9GJacwl4pCTfqgMvAM9lxhl0Sisc+T5PtudVxJa4CtpXU65telu+yf
y8r3ZBIPNiiyxtZ+YDugANT6aJCdsw+YhBzwgyLLlW7mc8cjZCxTSHbP8zbkB7cT+vCfy2/oYNKC
HuCO55K6U1vWZgbjZ99DGgmnyaY5yx/LbCLy4Kdh1XEX+H8WFJ5AnvQHeuB00MHXqsbDlTBTxYh9
l8d9HoTJSEBPGvCgMRaw0gdubgghbKnbgqabPp0UztO5d3nkKAsimbP386csjfqiqb8kSkc23kLJ
B5r7SaBHWCjgud/ph+EEYuKNd9HLhYswzBRXMwCCisdOcRxGV568XTuScv6Njy4Y505dCka4bvJ8
5/Ler+UP3+DEy8OEASbbkirfjCptwK9bW2VFT0qwKyzTRKwMophe7gaEnt4ZPixP/gxtcayw+yhk
/9QbJ2xuX68TCDsJcAFhH0HIMh8s8kyIl+YvjbjdaISxKWDAAVvCER7FDtIyrx0jwLIwj2CGX9vk
STdRCA3qHZbYmLEcwNEIPIPYQQ+jBP8A7XRpR3iNQ1xTKDYq9o4TaSxGOmU0HvpfYlnXt5L+1StT
APjBjSgDRh+f6/rpT/7c0aijbCOv8ecDUHkvTj/ii8ZSzM2kK5rpc+tam8xGwpybu9Kw0mpGkClt
Myd0jccEhkm73iz8vytuqKdfYtpskw2shCLJ7z4N831Rn8MEOhLAGzV5k3bUqB2CID0D5I1q9945
otaBBN+TR8Ej5gYMCjiuYIj6XjjmNFfWSUI5WOxkonCVQzccyTEHncuGHKb/FqigTPWA1UrGZaA9
Hn1PFNFFfllRTnfg088FLApGB9wARQyK2CHG+tQYEuq2KiIE4U4xaHcixdlulGm5L96qO0NdJmqW
b6RNGSrQiRNNNoMqMbUoNbhs0oxa3dxNr3vZdsiUwBprgGAD823qJcbDD88LHHV8oUkJQxH08eQo
MVqfL/X5ZdiQXk56LNU/4AANlYkmHfvY4skklLcUp+iYMfitfCwTid0RDQchTecMLBIKkYAOc9jQ
77RrOlrEHhyTlaJIIjEZHhVK+5pdMxqK2VEkywTupSf/aB0X7OEqP2Q5LoemNrT0/rK64ixgQoPR
Wqt7kaHUeu+gXSCMdIOwapjuw0gcNNt8KIyC6QkPEwaG3fOQySM+/80YcCyglCZqG6as7YAHmcEq
pOZBhK1oaoZSbqDf/J2+itW4OcNvDPNAQGxYeKQuHL+VRiT8WTW5CjFODtEBx1havP5OjWF31QIY
mdy9AoeMeJVWmo9ZwIgaTZ5BDmbbzQBBSQXawyglGhNjvB+Y2FpVSe7x7230GMCeN+OjLvD78LwY
U8WCl/5kStBsbYs3euAmN1hRCHbCNAJ6gwWFUnSL5Y/5tk205IJFjRhmv0Ig3AqNbpdRaB1XkUW1
bdDTYOiZKFKgOW4Y7NQkhz+EWQs+hUCAl6szXdl0Zr41biOcLNcXBwa/UovtYlimTuPK2HMJSMbb
Ck58uZrDIqsIM3QNot7MHrkteAGtYpYyLSdb6/iQbH8rhauOWip6MToaewrEbEbz9eUap9WdilL6
8/egOMZqiQJyl7RNBLzl/McnLqc3VgEJ18ATBuixaUCjMMjORqg6sigDMu9UjQ/u9U13haO+5Kjp
QX7kCZNAvnP5AgnAYEiSilnC2X2lVa1F6GtkisgeF7+J3r9cTBhYjFdBFmPxn5Jom0Cm+09Gj+fh
qr3sDwJYme7HsF8PTpqWzlS0I5qiXNfHIUsKNxbh/kimfu1kHsMU79cdCKYli6hwbIu6tEB6c/Hg
zqCK6oMVl1YwSBfU7ZXtRvz+leO5J/x35uhn4SFjbemUkCLFQKZcXqqwehyf7exIf4FfR8J39lwT
coZpIA4cD2PVP3BUPRHcyOB4dh9xb17JLrNb+4HkP0CgWlrmSx6em4QUhiXEkWDzzvHHfKD9k6qu
AZRHjDGjah1X0NTNx8Fw+1ryTyhM6egTb+BSI+tY2lMG/FHqIWPhUFd1Pu54FWO9fZOI/50+kY+U
pLXrmYVAR6b7YlrjqVpYjCskbS27bZCB6p/53X9sEv77O4y0NQCfmIL7yKcbkD7tELodYNDjunEH
L7rYMTio7ik/gw824esg3tZFkUGQ6LQdNK+er4AWNmy4KbQ97cLhvVblQyXFBoUzX5oJOImoNGrZ
nMGOhOJ/CTGZe5iHIxVOmgo3+vvZ2R7vWikaDUoihYkPd7Ui16sBA0/WMgRpkxXE4XHGbMGvcAtH
CtEBPt5c+NVhyGqrbt9CMgxSjOxfPbjWLhQENM7wyaYPFvDEo5pUcuYV6bcuIdoz5KLS2hU2KA15
BHPXYpnggFF6ti3am4CxBryRgFwY1bmA3vHUrOdCauJ+p7nYOJA3MQt7vKiTCHgdYbMMkKClFj1+
9NPkn0rQZbCDvGQuZIq9CpwcUseRPlJIqfgR3pEhdnuYjl9G14kA0jxxPU6b41AVAX5naNF4+znn
ATyWt1q8j4elviVAfxWi0SxOmeVysLebaoG6dpvCfXHeDHlo5Au55Np6XKsuELJ9R7HYcA+c/PLu
Gu7+d/eCVszCi/xJW9DHHS3PNORjUQm2fagu7GlVJz/hHve6A1+3kgl9Kxu/OWpNGUOZeU/FDlwZ
byR7IhNnFzM+Ui1GoKOS5wFGY8+RW0aM+IXjn9KeKMRcfZpiT4VP+sMdyIhglze+svU4dyzeNiqc
kkifkYGM0zljVkfGMIQshkldRbOcuSlRKjkK7YCOe6t6VKgslPrAUQ4hyElpepmCBLHG1WB8TdDR
wP3q0c7Co8iA/fiHv6zDiTtUKdCVvzh3x4TTNj1QElHfPgGT1hMR4+CmvkpX1b3PuaX6jIAVOK5Q
kcowiA7YrwPoiPXOUfifesE7p4+d0VydPcRoPBKPmnVr4aBGe3tHwyQjU5TLCzAzvgjJku2/93jt
cjgsTqNHvVbnioXnh7zsAVtwzHfyN0K145ci2NOtYsnwBenvsDmKSA7iz2MeJ7TVjzieaxXD9/cp
5gcHzBIlqmXP/fp2g9b/LRJEBnsbHN2prMlmaghdK0NZDubzd7De95vFDjYUj5Wx5xfMxfokrN/F
7yedp16UrDq5BSszQjZgxUCHM6BQxPwukO3OD/EMbABLzhWQIvdA5muRkLvpNizs88qUNzLCsJgZ
af8ekJwaA9fReertKkF1B+WiiMwIvWMxqOZylHrCTc452gge5dfjDmEqZXSPltEbbdU6Va7nYLhA
IbAd6f1kAuzvQZkQXhqElbOsLc35eQZbDJCgx0lxQC9EeU/lomCVqvnh7ticdnLXsTI4GbAWfqNg
XO+9YarjEI+eIsM5uIGg4YQTRt/Zn2bl2rbwXNkd5/M3zJcEN1iwv7lhnKsxdgkjsIgBXv+x1Nfu
9+gDfbVvUgXzV6PCMrgrwXAzK0CFBFU1cAQ5WdobS0t/pyIs3duxOLAcvzObDG9LeBs/GKZFhLGf
ei4IBCFyR+NmL7I87OAiRFdcKQvzKxEaDb3M2k7a7yLB3uazPzpOyT5z8OgCeNzHjYRlhOtq6GSW
/qCDkx776vk6kwSrCKMCFeu+hDKLUXOq1zdhqEg+tZXcLYKM+aJ0Ocjx7NsPGvdIcVYvuDm5P8/q
cnpc7VwFTjlqxCLnAMZtlfB+ozUjnKeFXfRin910Ca79902U874J/hv7cfoBDB7XhrH9w3tmzoQ6
LyE51LQGPsyPS9wzIHJk/cdSL63gxkvvP/tlnN1rUtCuQyci9cWoLcuMjQTl78QovNUA6OVGLCdd
gY2rPkH61hQXTV7qM1IMO3fX14QLG83LYr5Gnlz0qRbM/6HRu1BUMs5BiYSuY4QzQAg5P3aip7MH
l8tFJ6x563xW/lgcdkacchfd0maAM6Z/IaGIlgF7oHyOBC7TlytWMGPzUE+YJzgxxF3kWnkvRNpx
3y+rGqQA368LCUhWdf8D5XqXjC4mEyFiu618Lhy6NuC3TG62z251TELCKlA5+mOq2nsXwkcH478k
WfZU9a+O6ptxvmcA33h4mtQTyHp2bWUmU5Bu2vLWZPLtoDYcTDIS2RscNRjCxFmOYb37PU/fozMz
D8rNQsDIozjstBNbHWcUjuIJVuTgHsAEJMGci2kdXYZQb5zJa0Ee5OJABdqk8nysBUs3B4wrRIk/
iD1wUN0xAdWuJeSZBmKiqTIlmZtm3SVKhisVJqf08VJAF0d298zAZx6eqXKey5jB1Q64oH+Cj5pC
jPiN2Qpu0rZDa6CtcDGjgVDBPEuidknOb9FHPNYJqREP2RcrIV31Q9mPG27BQ/n//XcvA0NDrc+3
enO+7rI8uMz/a+NnF3D7CAzPxg3TNvbx5JbQQSzjtoA1Jw1e/WOI5Vwh059Q8a4BC1oe3cfDRGze
aZcE4kT+0imU8TBi/3D94k2JBXWJQRAO1ujC2LZlxt2WJmhZbockEo+lSCyEevLvk58wV3Fh8STv
33l5NdrOtadqvdZbilsXBEHnwJoJ+QFYqclM2RrPf2VXbo+HPrf1AcfWvLu3Z3QX1E/auMFKir3Q
GVugVGHIZHm23TR5KmrvnoEfRykcgwjlyAFgLxkWWihEvZg0LlkgPCw3UCxhNhZWIiS5thDmpwkm
euSIPRLbqPNMj1YNYx6nY+1hErg+kOuBxl3V+AVw4kcq+M0lnTEVRV2nTqobFXSMVfkwty+F/zs6
hlrv+Mvuu3rfS2vd/cMCp4WEztVM/9ZrlPnNfavJpM7zNMdtimU+cjQAiC3ms72rH0i8IShxN5Rf
DYKEE75FgV+b6V1XZWPbtwV6MHhDUHAQyxZkdTciPSlv9J/xsmP2U+8rddpwLmYjW2Bt6S1A5f4w
hoCkNw6UYw5UxAR0zs4g/N3rDDnfgTgf1Ez590daAe8AMgN0eFiqUeSZhPcROuZ7HLFHb11oKhU8
Lb9Ty+jsGOpupqpaePXRcRIAPo1OXqTl3YZ49vBMUqrCU8DlzZrRofs7yDK+YytKGPRHWAfcz1gk
ZpMUmTdBGV/jK1jMedKvoksIVmf9YQ5Ln3kaIS1VVttDFk4FDhlY9p1VI3o0Jr93NdTwcn7J2w4L
kUVd6YYL8eOZZeyLaJSVNOomyzqg9XsDcFj5/bNFg6sIr8fzxJrM3hZCPBJ88bK13G61avnaTpzr
+jSYSaLYk4cC1Q4I6RYCrX23SkXCEhup4uCLGx5EgDtwrQZ3SkPyEDk72y09QXo4WQXG/SsAHEZG
mGoqIeiZNF4wHXGjNA8kqTIRw5aFoqNvn/jvG5h5isseXGQ44iEhO+byf/yWW+IWFZi//1ZabjzK
z/lwiT0jJ7jz7tcsvX9z8xTvcTvtEcSRD70rfNaeC+wtC7CSEB5wk57aNTiRdxeKtDRUDW3GC8bj
9B/HhP0TPzjrwydopNm6dvPuiFzLN3r3QekSQasaG1XtiIbd3sliHgKIKLM4m86jzFXdGRJhQU4D
e/77PhkInMuk4CKK/Lne9FhgW35/bXNJzvqT8BEBb7xNAEr+rrUksncqyChwPBvC0RfZjEqF6gzN
ATZa3gGMAoE7Hc48RlMSq655cDYR8nTNQNhQD87DI2n3qOJl7WbtNHM22g5jrdfHnxULgtiA2xeh
bJLfuDH6oSEEonSnQ+VLxv+lB40fE4pY+CVKv/qYaiOC+d94ICgIJ5Ny824f7hFguLpMF3Hf/Tkl
vtMuqwoGCagt3XL+RKIIMP3q+T17NqRbOsIpF//Y/DKAtTJqvwHVFKm7WfKsyD7j6fH0V+WEVT6R
tFGZfYpZpAwiMN6Kzbhb9oumzI00fqGvY6LZF5UCqsyRSNFgl351xpCBOxXz/3p75GTbtTdOGaQM
uelrwKEBkysqEb7TrDHV4hxRpoYmKyjNjj+0zDNwU2NMhXiiqTUqbghCqgPSVUFZqLx9yy5vYJjm
Q6bi5qtTHoSrLLhi4IDHFyPw7Mv3OyVsPlcaaY1JLadZLwSFlxwq6gkl8+LIOZcJcIsDznnkiSs3
7Xri/v59AYgfcp5vHaqUdplmTza+wp9SY522evmHL+yyzLkcqa1fCKXyQkRhD84yfT6Pa5KL/bFL
nPZdeqNZ2GDbEqQN8PXok0rRaSvZagWXyP1PXVUt3O0NW/MEqRhppiOdr5TqYoAREMfVvHksVNh8
+nFNfR3dyIEeKmhgdS8TFk8+z+2/TonU8DYTEe5Bc7uwQbPm6wk1Aej7hHIHmymnBMsoYZVBnN8f
pMa50Ng45tIM0x5pchF6yRhmIVjNxiSgUTK+3UrWOp/yoKoz4iWaCcp9BQu4zWx+QFQ1S/QNS39c
EcSaJH44gZg2h+UoeZj7ks6PZIKa1iF7/GFA7RvtfsOYM07KrJQE41X6/lo5uSORs90S1WekMo9y
hDQ92iT9y00x08d5iZ3oU5uOaoEOjq4D4m6isOIoXk6ok+Ua/wh9jVW91mVFg54DVeVGIqQaT9Dv
nYOCkCH0L5v+5V3lDZGExr6K3BnwUCa1nqNNb82syYqad8lgXtalccxvGtVDj5O0vO6+wG9KmFqv
tqU+BTzm45yajok5Mb08z1CZ3HBrwTZuV2R1pybHEl0raS8elBOSmYm/sWPF05Arsqdn3pO9pohl
po5NMntRhPdsNEJ9cyk/pFc46l4l5jnhrYI3VzT2iyicFy+IMh6DoynaQct8joI8X8d+72mcs1NR
V59D06U+PEAR2yd63tMJt+OGAjuBCmieMphNA38dME4Te932YWaVoSPzNP9bky0dP5N6fpUEvlm1
xXznBZzc+4zKb/u3x9zR2dJMrmPqT/j0/zTVB8DNl/PVzUK9mGp+2gUjHA5Q4dXtiAu5JrwOW+yn
VkOTXKbIXjiFWeEQ6y/4mNJ/gSWJKGwOjsv7TAIiNJ8nodh91zFWzMagV4v++1625Wv2flIkMPFc
3jpXJULig3E0i5pffVouXkm2OLpSos16frd/NAFOIRMWzh62w483F1l7bWaBC3nIWh8llkufKfvU
jWM3652Eri3LhE1gNxlVP6Yebt4RoqKyZYYrJ3A+SGCqFgo+/BknD2mq4/jBlX2eQIUIpFQ7ce0S
uWk6EG0elKJXI/dolwVxxLE6McZ0SCXkPCmZoQ616ZInZw1sz0EgVi3DKWt0GclwSxPfwpPyPaPx
aXoBk5GhMV9v9s/zOCkWZzt9vxljd3AUs/WogbkO8ySm8eC1OL8o3ZcmM0FlUXYPxQjKk7varK1K
JKmMMcMiT1RJuq3BIS3RHNynHsn0C700jfuWZS1MJUAX6GioP+Huy+66wVnEi5lI8Y7Jh9V0qY/P
YQ0GukRhtUKSsOU3jVb/HH2P/QP2K4NQH81jk4co13so0JOJYuIvV0jXVqk1nxrl4XHpD7uOqJhq
zgvxpMRgtAdY956eq7CbRYbgjXyBAJ+xCVjWwR+VcSXkoxhVTXLefktN5jC2L0W2HyA07rp3Oo+c
lBM4Gl/JQUcbPI93G8tpQDHkeBCPGcxUAjmSFP95Xq1tnhzByv7tmVqtHsUKP0gAJo5t+opE1ZH4
1hfnaYZ4VElax79j1DZ8EyqsYPLp56nEctlqRo4w8201cpfuOTgKY/Qun0U78xL7Oka6bS4A1E2U
8IcyjZkAiNMU/QGbOTvzRjVqJDHuI/5RDC3hKfxM/bm0ID6OMu8KdxqyUyOP5uN4CTpEw2xmOXEh
G5KwsjSGBvcaDUPt8kzU0Pvutc2WZi21G/JQ6x1nyyqi92L655+MO0k0LxddlYo4r0M4yabQhOnl
9WjVw04ubKVMnWewAE8+FlNDo/0QKRTzBTCfBf1fSImU+QxUNm1jnSPX7iz0L+Lo7K8kzsx3t0zn
AiTlT6pY0L4PdPyewlTtOk1GuvY6d5IKxbq1ZMYhbgmpX74Zdek9+NsQZwIxKqUM22y62tImgGkP
jiCMHWMMczgxMV/QbtR9r/SmobLmFGLRFbrv9AxE7H3pM/9uBRppiGJG76zccqIzFESjrDxU24S3
q1s+CmUrjJ+UWlV8P+FA/8pHMuRb4RtSnb32ptr3iHNa8iDJjzkd3Kv2A4mFf4RVmBNCOr6/Ql5E
WvXhsx7seyU1/yzVBnamBVfjP3f3N48GLTnw4wN6kgerSaLL6GpUn7lLJQAreqzQCedhjWZIqy7M
GbWW8oEsEzGfJ89INP0Zs8mTqkv92K6I3SQxgjyS48r92bV4X/6vzkfeWvTCccDvNjg2hlOGt1tc
3poL+IeJY3GAjcWGOWHTOEVgyd8ppNHq+ReoLe+XhrGvONZFSqII7uMq3aFkfqQX/VHNIAoQ/oVH
l75fXuDYI1D65b7l3+1Hf8NdW5Q68OAApGNWPmBfRr/T36Jacyj8Ie2kzCCzmmtpJU/qWqYj102Z
F5uLC1EMN+yMmW4kMbwAVljizQbvO2LBZvSYa2ePAnuT8rrY/JQpgHvS2p7P/0mQSe12tZ/xvNdT
zmZ90lrnkw0eh+32SgqHKEy8sIcaGIvNd81HGVP0e+NrDpun0cQ9L4jDWD9FdOVdUfwNQ25r0s2d
AZVKyNLhnnWtBkpim2aFgY/OV9eha2mOcGtRnMYoO8R2/4QAdC9V8IrTvztQdlTqtZHhq61EtFT3
w9IJDvbdymHPEtIV6wNnK3ps95XuxlrOH1+t/QPI4KziJS2vQRT3RgLsgbeWf+n+qwHZFc45YJOk
lIVkCgybw/qb8NWf32F2IhjS0LsLuhV8PlEBpMY+doMXWob31xvuoix9Vs+K4GBQPh6xYWQ4BkaV
+pr+A8Jx+QJTn3Btal1R9O0nPJEQDzT3Q27mSO/srKBNriyezOEWmjs4fOUsn+RRnl0/WF907brM
lXfRLrNCMezjhxDXNPKvcgyz1weMwXwo3z6Zhszq4z5Pl0vGxIuIAVclSQHNyEOgFwCXgyBqlcrj
lbHdZ05KGZqtCDMOng5k1Q6nM60UptDvTnPG/ro4Q/LV+DZRPnoW2S6fSgl5Y15gKT2m3z2vVY8V
skOPHN4PG/5laOoNUIj5ePWoiP7bJMZJRIuP3gqwMGVpMgPWRvbuM4LQ8itAXIH1BPmt5gKoztvH
V7c12kLhOVJshOrDShNKisttSqN/JBeQyB4JivKZ23kqUvBXlI3uvaSfS6Vgo+kgUjO095YgJs0t
REEKcK4jbP34Osd1AaaW0kEgnyvYZFcRDRY4IvZvJuq+lE5mj6GSUDUovDVgrTQXnd70DHmtsWY+
3Wi1PthVA0/3xuH5pkPlB8qt3p9lORp+PWa7bKxXmhCvZAjRRYtKX5xJUS9Ww6biQmopg8vVcMYD
Vzp50hvSAc1xBn2aroQDz6Ue8cakqLFByrX0ozyJGbv+OQ6tzrGiAKj9vczn1dyowGLd6AA/oeLW
6zwpwXAjy4Hwq6H70QH4cjZ8C6pXU1OZf16UFQRMLgP2292Q27vI0mw29/syNmvEci4tmkWX6MiG
qemA6fJEWGHyPNblDQ+j8fmYaKxuPqy3lDAJkDeU/M+9edL7+HExoJ4x1CVO/dcvqfHi2xwQi/hJ
yFCwd5qBMfaRQBM0CYbN5VzfFEkOl68E8IP4c8svouS2TEQae1snvYlpRKhX/HPGNFycKiP8J++U
FSyZ6Ngc+Bg4bQMRQBSOs26sV0x93LNetpmR4oAMbeuE52ex4ufJz4LHt4vJaOigDZC2sNcHwdmm
a17RBbqZMxyNOT9a+FYQT2xHAQ+SD7y0etCgwX0Ko7UNbTdDvaAc78WVCdC/IO6LC4c/wveqOKbz
7MVpbXjtT52dgDy3bIRmNmp4HF+NHomeamsKbApEZnJRmyJXCBSDXuUWf/dfwsgA5YLQyLT/JTXg
ShjBBp9ISgAHqqcjODPqA1wsYXtXWDaq2fzTl21GUgDUIJ2vspFZMY8pvjIR+V0rsIl4yrEuYMTz
vcN5Z2HjRQBjdizDWX5GzXziFRIvxGr9bKcQD+P042O0fPD0a8QhchAybKyQMQn8hBjutyQoQn14
xZm0KcJNd47HGkXQ3g5KS0fcCzp9NuBLkT4Rh2ngAv7Y5NYKm3tHgx2GFcVF8oCB1d/8q/b3WfQy
zlIqUh1E4tXgoD7mu09YAiltQBJBznyaictrRuIqhXHiiidWjNI6dbuop6+xscHvC8nnmVB4WQjc
6dhvSP0F16uLw4wrM+e8Of9TcZHuFkNHzk4OetZEuO+qoexEFk6ajP9E/zbTa2EYqkHHKsrt3trh
kLqy9VjLf0S8Iz1+rxKlP9IkGvsyx41oHg/8Q3UFk+7vP74+6VlXihKPjTlNXp1Klb4nK3aNGUyk
caMots9ei04r9YABHPbqPCSKGCbjG6WQkDRsMiXpglkCVLEsi3nN9hktGoNuSJAkgHJUzNKNSOvj
MymJebKt3ntEOubjiFMkJM+QEEEeYRLcI8CyyJ0SBoajjySsh04+s+7CYeepeJFs2Wn83Wm6XIaW
mYflYqSRvNym3Yw+EHeB9IFFFMxnw0e2Hx64oX4P6hJcrHo72DIZJFqJvKTgMFUZtqJDChzxGDhS
uiMIhZUiNwntPB+Cx6tKJ/lFe9ZVgJdqZCS2hD3NZgbHwe1bVuds5qSLGD3Wclt1LtPujyh2L/uJ
r+be1lDhfiQhTkIZvC3UjHMH95QbL5jAhpNW8yEdLEs6g17rxaAiVSiHXph11UGXLwjK7xGoscc0
rzhzVyGo7SH+ZfQTNG00xjgmMCxAeSHeWmULTVXRzIcfSNt9Egxc9TmnFE0g1swfh5w5AVk9g1gl
vyEuWzh7w2tYD1HhFPrq4mshM+VdB+bpsAGdOiG0FT2uWxOXK+8KjvT+EvVkYydKjOXQqBk5gNra
azLXuM3UczMDMOcG0ZuD9aY605h7K7nSFH4Jwmz122fDt33R9bqZx9RVHSE81jiFN6k77hjFlKRF
AbBw0ZyFRR29wBvgmI8nUXCynJhYS4Kc8Eh8pVD02EfFKrjhJrHLAO4uBy/n3zJx62u/yT3TmZsf
XepygDmllQXfddiFNLY9ed33IUh4MxEtDiwu+lA0B6LcpIynsX61xQ8AY+SZtrih+ZSqLoVOa3OP
ya9QcqjbedRil/38Q6lSpE54d93a9etnaLluvO4AsDv+A02bbQ2bB56bZh9hZds8AhiVa4vuzNSw
7UZcbWoj0orzQAKmbSetUnuIr2MBgiMwOu2yzN075SgX0ZRpPKdy62woauM6iRnBmCfSnHs2ZOgs
BiGex8rKc7jTDuc21K4BwLJkCWdLCaNOL37calkVy6EDaGnDZgb3ml+r9XKo9ply6nCS7/YgaJBx
L3cEK0Dd73UmzpwD0mk/7Idc9yfwLksW0fgTgu4ofsrZkY3lbfuARmK2MsygwaHgbQ1v9+kAWnxt
5BIwz4vZvCs/IDzbsTv0SauxMJYA7pd1d8RmSSiA7jR5OprE5T+ozwzN07/SjEcZQV5xMldJi3yD
RE0Ie30/XtXDwKDdCDMEX3LW9E0NXOJ8JsBj9xCXhs2T92gKv3FY/PRSNmbORaIS90E5vshTj8fs
S5en/Mf+Nrg9c+sj3BCEUsE5Nl26Vr9mtMzED7IWueF5rQTQWjSJpopP68eXCOj3zdC9UDl/QyyQ
Cpw2SCpwiZTbS1ki2iz4Ev27NSNDNCNtZyGB3rZs3wIo11hyMg4WDWblavkpha1ytLQpTQEuMtCD
SCzEQns0fdaAXgolDWKE5G+8vVaSWd4D4pFFHIGCaGRBQP6Bji8uIWn3OviBpIJSb7pnRRMS3dnb
MTyE3ZVZDBgYwmi7azRePjPajvD2ZlbmINXiv8lAhFSbuU3w7sBbrjzkjtwWcF0+6vy6rePO/gLT
Zzk/ZiOU7gMdjsCaUNEaFSwiT6Iw7IJ/RQHF1nB2h9DBn36ssSes6VtRu895GvIACM+H+JmDSali
OsuWVvikhmC2XllF9rfT/fuSDnNwq0LJYSkgO3eq5Q1cpI9skPcKoeWqvluUxfIxN+7iX+ztpwRN
g2E1B9ks9bArVW8Tetdzr6rAkM6F0wsNlX8bpoEmXlYpwGZ1tFbxc0Afr1o4x4q26s3HSryWehyU
9I2Tkubi/rfOPff3nOLBJebTQJe84PWynAMBTevFIXT0iS9ifTd/gwnqBT8d9XivCoM2wpn+XH/e
P8014TBx6qqjTtwcYVvFNnxcZOqZQdiILuX+QAv15FoK4laihcuO7Ecv4bYRbdFDX1p+3/yHAnQ9
G1CCVKYrZyAS1eIg8ZhN9EsncWnoe2TsYFSUuWu2Pry1ohOY7BEJvqTb/YBvIhqzR5/QrkrrkFYe
NKt/HhsDk1IXoLltUegzTKA+/x+QP1rlrjxiHwMB7I/O5esGkCQ6xaFmPAmtoO0o7SVyqlTG7F3z
reag8FUQV8R1tecTh82lBuWyjMXE6nPn5wb3hogYHGvQ8Bk7ZvE/Vi5QSWwmvUM7hRjF0Zq2jDuv
pea0tOuaZdELtrAmMtRVAMLKYjIy9Qs3K6hNUcDZqfvMCU4DDeJvZPeqrMgjcTNCRw9y5+XQaYSJ
lx56AKShQTY3IKY0qrpODu6jwQAZTWM75ybxa3UQ3ECWLOUC+HmFsgCQr4xId0WOxj+qmYnfFVl6
Fwtz58sU+DE6qtJl08XVnOSYEPWO4Z9WL5jZUoGjCRi5fOy2o+4fc+5w80uFpcj/9ArfvPbyDK1o
EOX+3jF3wp2XhldF6D59IpMgtzc/4kepGmoVLHuwzMCt6MgqpF3C/qLJxWhcektPW0D4P0NVYdnf
bXEZmaA+W2q32f9zP/e7tIdR0eUE6vSIYhNDbwUouUv6h0akXI+b1AAGwzQh9lHEgFA+a0z3Mhye
2Gx4QMbE/tWI7nRRUX4/icdXgermKxzh03Qgjg04WVzefDlI6PnIPSZuOtn+VL6Bv/mI4C8PtrMU
dYZOhRsG6frlfVkClRL2wzrfJeGvL4vkN5n6ZILJmXkwGl3VvpTHEstJAQg9Q6tSVmswqPrylUaD
TjBmDrDOPSuTDHApPEX+A+jgjZ8vN18lLDUEf24WBELQSHoKQvZFoQguEjzrNPnTzvU2T7Y2+W+s
fdwAYyYcGW880xNKcxEmpnmb7k/Ygt83KFIF00Li87nvrwYvrg9oRAHCM4dpna5cCwP9j/SgygPk
qwgQjlRgfX3nLGoVqww23au6EZnTgo48tus7QSP7qyyH6P0g/DQWk69LAA1AAwxD7BVF3M2JDEXw
PKzGlc7gv2VBDbUHulmdRIl6/U1XiBp0KE2cpb9liNzH1NuHeYVUub49YFC+iYHxSVIPY5OdOPDX
3K+sPVnLveGhUF6r/PiZlucDMpiIgJBQpqd0ddAq8sV6F70sEybWGPM0Q6cshZmrOAiVfXfDL6wO
ZinIIlNO2WTGKlkrFRwZQSONnt1gZjWLX4MM/jZ6k49ch3pw2XZ37Ty+i9hj5ryzfH3eZ5K/8Hlf
G8RsYuuV1IbQk8GpQ/CdHedaEUN+GfFWxMQ4JVNePyiM6yxnQgpFsvMNq68uFYkSbJe45rwsJepe
C0H0udlt+5fiDFxrSSvyJUXJTu5IToQuSlxOa1tnYHT68YKVJkezLoTjXEwV9QX0Ia8fzT+VBtO7
jXBXdWeElpjg9NiwAPznPytase4LW3+U2pdQX0hSmNgticlupOFc97DyvMvYvOV02Upn9Z+wNMjX
nSK8v7SfYSyETKuubQPm0tM+NjPaPyxwt0U0tt76qNKn1Vi9bLMbdOkdOUQ66V/ClhJbjN1t87Dw
ak292/22bkJ6sY6TmjQ9+1atUvJIqptrGjiGnwQ/NjYAizs4mEhcChS/RoIwT7jaYTZPQFVTEmls
rv3aWYOgAY+2Bx+CJn1P790bkqlieJ28Vy2Zc15giqGD67mnd0aB/twFmDwXuJXle83dMxkwtNnL
kPfhPRlrfU9JjCyhNFenmA3Qx8zz1WgS+yZlttLQrAETaGD626ZPfGuaoUFQR2uoUYygpPGxeLaQ
bWdck6RzVYYpemm63NYmP8J7xJnQgrVCa5POj1iPjviAzBEnZDGwy7UVFJYottfzRGN+EmkWkMgR
MtUse49R4QeCcdJgFdAu1vs+pyuAMvlFVAy9Et6KfEd4KiicOzOrFQbnR6Y5OmQZm16nI0Wou+X8
5yFgNHdz8g5sEs5QUPJwpyMyVXiWUdiVARQb/+bHvE9nzNe5J+xbmyHBXR25jMzK7nXZa0s0W4W+
WS+sOwCi/d7LEIMndYWij2b8OvpHotTDEsFF7bOg2RY2cRh5vV04zx182/WDI8iGQvO2HHm5zJFb
RuX1zJXGPVpiJTPKSTnHg2ZUGv5Dw8svTU94rewquvENeOjunaH6U81I5hzVpUEKp5dGHmWyuo16
p/84gYM/NOsEaWZrOrEvesIuR7JwgR+OJEtErFEvS+xmTE75B51vmNcVB5FKIcOxCPRTwki27519
AyGY6MW7p7HODG2bZTx/Bhbmo4LRIOCqeIQlIl9weNh1YJtKcP12A7ALXpKcwNqQU0I7KaWcB8rt
nTr5QDtMdsqzKoNHS6gH65u2dvcWqPaC3ANeq8vmMJr55suRutXXpQaKFLpsdb+6dxwI+OInT2Eu
zV7jHBYcD/RBjmQ6By8CkSTdaOvZV9uU9MCcZN/O4/RPpUk4Vk3dHazFpZ/DA+yVvvKWRkzfsp/t
H85G0wCSipsAcQJGcwOV19BhWhS3uHux1l6hGw9DKFVEOhBPsCDdMjGxeHQbyzdCcqa/orMNRaCK
nUgc5O8Q6gx1NRObCY7kbDM2eC7rNpcAycZRsN+7M3C5uMbP4Zrr+qxakmBONpMN/SvGYuXFvNt1
rb/w6faZEznIjai8aXi/+bZ7tF2sy2c0W0Qob9eYmV9nblsvqyKIhm+y4RDcl/Sl5/HP1FgiOu/D
Yj3n75T2N9OiCVYcj/uHaL57ovmvIhFtZP70VzGoM8B2EQUQcxxseA8Yf3yhZCFxlSqfPIUYfeth
U77cBMd7Sv1siqI125vczP3zHMFZRl/dTZ77Kdc859Mqd0KwItlMfuO+Tgagu8wLo7ktH5ymvD1R
tI6Be/ZOT+CgTOEELR7kB4vkN2WcCWMwLN3TjFSVvIWHlizRKdrMVWI2SoFmpRXpyZSMqgl/DGsQ
yNx1Pp+LwLo/nv/0nS7giPvwpKCxvglm7tm7YSeI3q1/TcZnEORxIEdKm6VkQjsWwDciqyLlhBZZ
nn6fGci/zMQdsOY8l32vn6m0/iH8D8E1JBhyKT339q6q/js1PJ1HSkVMBGxyi+1Q58bwjY9NaEh4
Je4RpX/edo7DiluScV0SZwHmeXeDIsFhMwLLaO97v1IiivTFQ1BPSXSuW+l6dBPAn/Xg7R54Mitg
H49wsbaIk0aEXIbcQK35ndSWyxcmt8h28T+KufZ1NQwGUfngt+y6SojUdd18Y5kWnL2/j+mia0DO
3QQWDq2/N7oBSxtqxVk/Nq9hX41QvnPt8nbUI5hHxjiymPi58c+pjN/93iamCD12uhUGMkhn/RTF
vTeOYDE8eGWRYyDfsGFOqpFg5r1O/KQiLiv8lB49tyXWUdVbH3WG8/eQtLF5WvVu0QmbqEJUQGkj
0UrvOk90A9gJI36OH2iRD6+3ilRfZYpMhJBzzgIDpTlpw/xiPFTinsNUSu7Mk35NO27DFc1c/eXB
Mkog4iDir90I44p4KekDLMkOpPq67lilEV9crWwSNhmKixf+VDSdsnYHZ7HyI90OQLlqtcY6wTG3
hT267Luktbt31bMdoNSwFlLAdgQ8O5NFmznvY0uv6lD8qVL8r4hngxmRbei0nyEnZ8ibYd2KVXkp
jnACRsJKHDaYb7f495fY7XcDlRBu4iCk8DfZyfDr+DZrK6C3LJV+Nn8LPoX+DNP30Bhw7u226M0A
llmYUTnrDqjvSxhvKjiBkY8FhCQFnQKPPOyJXeHR1ZYFh3J1pu2DBP47tEY34ZnzWZhV98V6/O3u
9C3BNFS++Hyk+fkwg6RCPFEYmRo4ebdJSVI5yONNAy8ASDQ+7q5HMsD2EJfGEIolRdhMDQpU8Bbc
vx7VUrHdpntE1nnYen+Q2ZvUlU4de81KKvCyON0Ifcj2T+f4dbEkBSmipUK+uYOIxM2UhaMXI/7b
Ppeui55RKW7fl0ODutNiPI2ealHhczDaArCcVzgL8qg3tIygdIkpO2V3uhH3krenPqaoFd0bhjfq
QNiSLNMs+ix2JZ7TXmXZdhs8aHo/WxL+y87xeFv7mvwUsGJRk4gWannFyuE8PSP+ewtb/5mY9jPc
nKbJA2Dh0OLoe/Lt/H1BjbI4UoYEG82I4X/tDG2X5JuTkLWJquGquueqqFZCs+FmrEITD8GL6HE/
ncnJNvQ2/bLRUeg4rz8ci5I2+CPFNaTI+AzZGkoeeoYPEY9o6Oel5bHhz8mQrdeE+lDPPcWVWB81
Wf+8rQLSVQmDsES8ydk0lawCc/c2q0Aj7pmK6DvgCiNjPSMBSmolLGO/sqc0/F++NDKeG0BgyBSl
HCuN4MMHISogZMO3bbYHeIu4B0JYt0MnWObnSVHNji2HsjpzItDhfmCU/1gUmPdQyJnsa0tF4X9N
rKmxSF0osZSwKMYlVhin6bFX9LsEUSQFNlcCRpYmCDvyHq0F34vus+4+0EC0fM3FavB+aCCOOjxP
7j0E7rx5BVCnXZG3ohC0S/iDieS8dfHoCwzVpb5yR4drvCVuGZACRDCmaZZ/+MUp4W5EsCx1Lkd1
UbGAlI2WDFQjUFcHmIwhH81HQQxBreoovKVMnaN8FZfp7pazsKVOA2vK7zeIaNDHDUGUfRhwD8tx
HvHDhx+jbIz1PRjxX1uqGhlZrVRUzTxp6tChaUz8S4zFTZegN3ASJgou4brgUZnigQye9Jv3EbfI
evyzKO5FI/nQqCbeIg8R4lBJdniN8kYD3d2X88SmTDie0+2d9HUUfToZ5D60PNov0+qpn+M9d11G
vwy4OZet+3Ef57byu0oFXE/YnhIL/azZBxuoSYk5dCiwOPIafhPdF8XF7nBYSGEdWHZ0uoKsNUOa
bj7frFAErYZnCmCRKP5Q3PW1y47TTodXMzeOER1u/GaN2UPGRB2BKMVHxEaHJlJKZvt7YHUujIFH
mlNduDf5tHq2Q7zBnvqS1zvr1qiKgeKjkqAmDh7TaZMpHkei1ZtZcHG8dQZY90Jv6sdffUBAK7AK
2y9YNzArG9Os4ERj/eN1Yk/cUnHmzhCWGk/KGIGtlhxcPlzRvHim5q/dSnHGM9txomLkagGs2tnR
jxCqhonKyNZY8LA24lHecFONAbd3L9fLHosNgYyTX3FiLznkNYRZqT5IkjLQgRSC5BBAi89qJEHU
mmx5fh3Y4/OuFhPGCIaZDp6ycWo3w46Kms9dl7l995KQLodPd0SpHDzLPxzRd44xR6obKiBRco6l
7gVaZbptWeL1PQxH8WCytPJnggFYMEi+6fzelqGkXnfaaI0czFyYnKSkJg1De55nk7oxx9hW8kb3
A9CDnF3QhBWfEHR/jSYfvff0kqsO0XOEFSIkhPtvL8uQXFBiWatmkLDyM5clLn3SrlAJCg++9u2p
zgfHrUK0H875oiKPdlzBtC/fhLfN+Tcpx/XiX0jysADH9l3Y2WcbrcaBAVkmReSYMP0wG5ww3Hh+
ogw0ml+TaJC1XDd2DLLtNbef/F9BnccrjNtQEsVNOI+NRHeBVuY/2cC3f8mguKbHWLCvopixHVE9
pT1CRWxHldlMaRmQW1iFnkUEotLS4uSbN8/RzIsRSooqZMpFitQnuAwxNcmzBRwg6a5wPcxTwzX5
Qqg3D9/FVp9KmQR4KdI37fzg0zX7Bn2v2qbM4X8+PGRk5Xi53TW2Hf51XZj3p66DEqIj4XY4M8fJ
fcASVGrPy+JYbCcRQNz/WqTvDA9fyIiWp9kf9bjp9E7znyLw2cRC2ZFt7AGE5FIIdtrIU3CzR0Mz
oHZ70vbJn7NHYjWozZwKH/vXYMumMUwt6vH/lJIP3EuFMS4r00HvMPVTdSlkx+m73EXwwZALqLXp
KHHU2zI3bpHp0On6D4pZinfxVuBVKzHnb+nRA9Iz66sMp/OHZqUf5dX/91hpB3LwAx79meH1AypI
9R561kw2bLZeS1JRZpTOFLb7IEh9inTXIML9Zd8Sor02PQ12wYINyeBPmTCLn903Pg63rkc9W7kU
P9O9TIssRfWpDUmYsu+N18Tlc19VMmPDervAFcBZ/x4ZQYq67tON7qoKIRrtOdpmyX9sGJ1FZUQ0
ols4PXvmfILQhLLydrcj5qtFeUs2MUaK+0CwgjpSoQitAei7C+O2Wu7wVeAEwXZxQ1ZvcqemfacO
OoXVvEBB/RSlZH2idPfpwhc10sxsz9LzrOIwytWkWsiBJ9El1JoUNnrGH91/ro0i4VszLMwA4ub8
IiavVzBB6hqiqol6pE/h0r6/0NAFWQRMsJPLh9Kplm3yYLPkuOGQc0JEQIMXFsfdfqSo395RcUZl
hsiYOBZSySgTkCOI3ud+1oPY1cLie/iu5alVCK7fbDXWAIynMrd+MHFWdrGIH9TfDUBHb70HJQgq
X+9pVLFCBl5GjmcfpRvYKnsPti1IDoZknSsYEJBmTkm7ElpzUIZuhHsTNiSP7n23U+S6PTpLQ/RE
w000WnyXrt3n3GuaI6iyKDQvfJ5cvgdSoWLAbsdX1XEGoemQ8M6Z/uiZsYNhTFJtD1wrNx4ThfXd
IfFECwVG4RyEBelAW33ZG7Wxw9s082LsCPIVdz+Ri4E+gwVN5EsYO6lyOlED5iId8NrBejVu3A9H
eqzndXKvTidCqaQIEck8GQ5rlGOmzF6PtKN4Gjmbw/Si4lK5fnKZ1UhOt8cNXwBq/amUWYrgJ6Ih
DoQOiSDYc5HoUW/Zy3/Vj0+0+McIuELCyqVi7HS2HmbC81wEyMD64wGmVoIrC5zJrq3X2C6bYWdy
PShZx6j86M4zxNdx5afpXa2kUrCtdNQe354liixOxK/gWlUGmi4GeLMXONtnEqjpOE2MS+iEra/h
S8kN3ZNUnbbZmYBVbt2GymLTW1DrGl+uQUlxglpHxfB+dNpTWzlD10kWhiGA4TDcmXOnfHBd1nd3
6EO/n1y0c+M4rvNi0fVB5cHtdKh0YIv1FKFRdZoYue5vu6tbc26e7WP8gSSXsWbxGVfHpWNTQy7T
ER9KDlJTNylVZwttq93YY6noPFuZKuG1N85NN1S4JflOdUYlPG6wTJrdj9qQjPewY2IUVT/fP3kH
GSi+BJ1y+IfLqJkGMfqrpTcoAL3kw3rJZrpcd1+5saWT6dgX0fH63z1wLv8rEdoEhx6JY+vaoMc/
HIZLcY7yosU1oQuFnt0f/6HhjEWgAXwztcS8IGKNbA8ou56kbubLWJZiRMGhiXbUk7p/loUejdsT
DauROvhuUN+orFi6PnztgxpAUu4ej7cVtgzdsIcDsXPYQYnRlQgqYLEmwIzgSa+27YLXBCrnFhxj
hkAvyf+JEp2A54305SxoxSljMZrnhl1WcrdAxCj/XT985UzeA/COkoEfexqSR+EEHFbyZd+IUTJr
DaqIujbzSZFoN4YNBFrjJp0YZFKLK/2zfaE1UcRfH4HudUHLcrrLjwNomKDkhMYOWxNvgPASA+N0
sOInAkAMF7QEYtjB2O9cvNphuXrTMdpVnYraCxlWBqA2eybNO+qZBD4zitwAf3T/mZ5YxpU+oQ/3
f7UUnq4IYnfJSGVdp1GpOt5PQ5MHG+Ap5HTV1unC6gMB3r6TZU0fbTzeWgO/tHQv0RjlAeY7bIlr
ojss9n3SeyDdkRM55qfN6ixG2RAC//f2UqTplbNjPt3bGm0fAd0l9xgut6hIz3THa6rlyHBPjzoU
tjWslz5snLyUXYvCRCTAnJoyRIT/l6fgLtq3Qo5dmna5FU3t8N1E/+2INm5pvxkYbOiwYlRx0Zs8
jjhH2C7GpiowFgdbY8cP+iWDcW8i2DU2XmTVmwt74n0DbzKLUC6zrdjwvSBl3QmM9tanClZh1rKy
jO9wCegFOyI2BA8pBQdaF9lLzSKt8cC4WuJLkaYhhgeRS4QDmMWXzhfnjdchuN2RlJBomhpRtpWp
q31DIlkBpyJ2vjzwjvQBibdeGcXEjsugQDzy36hfHUlK4eB2Efl05jeQDLOIf1lFwAbkaPsIDASK
LMdrgdBKDEZgai/uiTN2PkRmcMUkAEIwVxRbcv8vCUErLcEdWjv9iBH8scxDBfVAmA9kUwpVAA30
0jxbt3Kle2lOUu1hzz2DxKE/Uig6oPHVqmKkM8Rdppzkl5kcadZ5Jb2Bltlcd1w1zNkZyJbs8sBk
kyJkduMHyYo96UANjLQ17defNbt2XZFh7bLpPhdNpl1bjg4CDYHwm2ZMqPKWP5PXZEblMaMs4U3H
MYo5SiXrqgKBf7iCtaSongHTWI6hKdN5ocZxzXBJAxO+EgiN7hzCu/amBVkHLwDc63pVV6puff4C
Dmxx29aP+5RcmDDZtUC/duD+7LngzzZOVBgQrtiNysrDjYOdfNnyctJKpk4i/fiUU8ggpjIrGDta
syY/8Z1sqWQm83Z5hHs9dX6sS4//thQiTMWyMSVWA8RDz3vGIdOQMftUtjjACetj/bjNAW3Eovnm
WeORTo4GVw6qEEhM6wICfOC42nbu66BHBZCbZf8sol4Dg/9FEMrdfEaOcWS6j5DIsUiVs9b0tX3g
mPn9G1tr+8fxFrIAw4hbtsowprVxFV8CSC/ALCdNKoHdjdpvyY7i0rBwztG7d11AzNZkgbNCMRzR
iBP1SIKs56ZG7NetnKr2yNujG0e8Cp4tqkHzxdXJp61KDhWQKsJVYz8mFc9jSHyZto3uTTrM0MiT
i7g6RMSwxAiw2IaCndK6khSuGxJI3vDsuccmYBbBOgVPnQaG9l9QuiPGQis6AP7V+F/3dykbKNn4
hIUNEJYwHK8QBLXG0Hly3m8JW0gaEY9T7h9onNDpZ9INik37s1jUKiVJKMK2cv/5tetir9NnvGeH
vu2ErNHR2K43jfPunUdyezP1LKpgra96apAPl4P/9PpUUx/G1UIw8F/3tOr65wbVR7fbmgGuZpb2
Qz4n40BzXbXuOfbTAcyuDvxQdbrpO6M0UdcrJGGEUijjClZ/Pp9vnc213hAkr/p7TXkN1DJPku0o
LtBmuCfijx++bPlC/4nRg+nPwY/MTRCOPpq92NASc5l4xSG3QYfK0akdCVzN0Uymp5x/cjouIPet
LSDzBlYgUTC6yM3TB1nQm9jUAsP9vy8xXskxtQBBPh5LEoxzpbBvqcFOESQOgCp6PI9j7C+J14q5
JEYaiIsySfeQl9lqGnEk8JwSHyRpbeZN0lHFGkzSiiH46H1Q01XQJ0ZhvcRTgJLbsaBXHdG1xVyV
Nj5P1FIif01ZKU4CvmvdjzSxcqLwwPzymiwsfqQbx5Avd5AsHi3fde4PFqXQjYNlP3JOLAGT5VQA
xjjbXju2Up5qpaCXzgLGMOzcJvX+Z8AIzRLfP1oxtauKHKoKXk485CZSlS25JkeIBxSzWKp5pY16
YSO3CgxLSUYqasZv+ybat42U809955kd2oNS5+OGu4q077QbAQ7GwYMOzcAnACSlBKN/PyhlXqr4
AXlXuFIs4RGtchuLQMom1QiwIQHNKwHKj3sfE8zcivoa39sKXBE46QQ04yXBwHZlGNzSj/EeYOX/
4ctP71scFqs/Hv3sghTLQrhzQ7TIxTzzwTmPYAVlbPqxJUmMaJOgPhUvBsn7FRIJGjNHAC6Qo4iY
O0A4TKAXRK4RDeL/gC0ppqK9HPf2KOSlQ8ojhx+Y4UvCuOgG3IuMuQW7HlU/TuqDrpXozvDDzrWo
dgX4c1M/Vk4Pdd8yD1w80xz1uk+18URTZpEPkC5TyINAwgVdL+5MOaB3CRJgA+wg/13K+qf97YwB
s6/rUi6QAL8z4dG3hzAXRrF577/yCqfes4+jwzB5QTyjSvgXfgsIn5oixLYWTNE8R0YUn0u7bW6O
50ElkVAggPLX1wj0Dt2ATkrno0sQrhIUnQsw8x/xkSHshBmniMoMhcT/qGfphJNZLPOnI8M1cjQz
zLi4AZK6YFxMc8LHr8DUEUvjgcP0g11UbfvaRb+Xuh26O2C2h68MjymVS/OSfQMO8Ld1m0LjTqE5
BPz49B2Rp7GENEiF7qMY++5yMu/LbfqjBqRyBwWvo/X//dGslp2G/mKN8g4SeOrDGZkZxQTiThbA
YCKfrcwgiYodyxZSeRSCwQ5vSSc7EpbNUhacEdKOYlUCiL1Bvb8JL6L7UrhhteuWfti/M9AlRXqa
jwxyC9iOL2YZd5upEw9Ujxaj4V3B3aY9XM0HOzxbauXdaRa8RdS/qa9w2VaPeskMYAkneslNVjSG
SY3kbO5jrqOIFKuu+EBDOoeKzITFxXwJ14ZN0GneAcveW+zei14G46MH58Uy1roW7zCaUBrIcghx
G/vikCv/JhPU4f8SChENYvcq3C708jRYX/MWXYJxFxjbucFkP5YINEyEWKI+Lw0pn6eSnkIzM49h
qy8IgmP8RIo72CHfn9P86ST2kdItWqVnWnduSW1A8SnpkGWRRZ8Ci2BV1515Kq5/2ro5zQqeUVf1
dD1Ul4W/CHyAV/sNwprkDsrvHZ4j6dxevMokmxzGqN+vdIjaW9KudsJM1TDBxLNYdxUlGNdUczpt
CHiNP1zb8V61B9FXPOiSExy+VNAZHzIxCSpZ+xu9AQfxsW3Up5u7PFlzBOdvEwip7+922OL2yL22
HEzlCbzuCVLmNyMqdjW6yGAffEezfy0edQbFOYUNINWUFjok59TspxNghLoh2LSQ4TfssGZgL+VY
R+Oqz+3PFaQOJqcTmv8Ax1lDf4FkfjkUKSox9wr86hy9u5el8MtKRf6Smg4BvZYwzIjCxbVvf4lp
+6atJzLXkQ2XWM5TvS1Ok1X3WuVUAYCmLEOv+AIetjIoDQeb79bD0FdLl9LWv788twDFxYV5s144
tDcYHInwZK0JcXZOPnyFvK5nOdMOchgpeXwL9wsRlNwgonLwePgUUuAoEBQhx4auRRlcxNstQHV4
Ufkl52qUfQylbZvmu4zN5WUxtO0I8e0huRPd1X+idY4jqpVc0uhQMkT4lIA1ONde1RJMBE4HGQsO
sYKa3huyBa0jzvAY4IJZFbkJcCQQyo99ZFA9QFW2K8K/Z/WcPAiYAb/BJYm9rrDSOrNhhMrI1BID
2jwf08OpctrjyAte8d6SgO9wC7o/HhpCyNUE1IjvsX1LjmLBUoDQmG6EhlQxifBNO6DhSkyayo08
6HbsVu/zO5WRfIBrViZYicgNVDAglEFSS71flavYDunkt5wV576+BMDkTF0OIxua/32PjcnVYujA
jgYZ1nIC1JAK1BAqYSo+JD73jzf0zDKt/epyHykypnsH6syjp0S+yEBpIAJHOi5NApfGAtr6niZa
wQ6hIQP2jllx7OpEWtcFLSdnKCgFVGh4/TOYrtnrEAcAnanV3GHUsnwZi5SPTLMSpBgITIL4QOID
qmG4MfjmeqsgWAIls+LiooQAD2lubiIL/TB3y7h1oFVrZOwUX173LGz6IbMJsFFQCUmlebB6/Osg
bnaYGcSgCcwGXCsrXTCDqoEILl7CUTzqV9/FCDTyx6uvQIyWlEzzS0kRqYpdsezGFblQT3HuB/Wy
YZ9YUsQOz1A0wLtmC/cGPEzee54GnxR4Njs6RO/TJG+bfeV3vc5zRCrqDL+YfErCNIZkDq5voNc7
k3YyL2PEsJuiTpK2rRKzIkkfZwbnP95mCqEUKzAicqP29zOdlegQ94ogkXzLex1FLJGCYJLs02QG
efwzSHVc3qc47KVzQctwRWOpLBOZBI8WM8FCPk977uYHliJU3Ll9B+56JlS1JJpGkD8b1jwRwxdW
BlG85wvNMX07NHUzxqXvRKkuDTx4+dk3u4GFKTf71rQLdGa7DC5kqEwzvzg6iCBy1XsuYDcI3o0J
sSsmCUVyOl0oKKuqWXf1KDegTh4xPeUAbvetm4PLYqV34X1E4EG3FRB1iM20PSa/G7Jd3T/YLLyd
MCmDR+BqJnMSpyUdnCB8+udDzCyDRVSeRswAMpIBgM/b8BkIHczNzx1mx/NzaNWmTVNxkMllXuWI
g/xSksS5HlzGMxpDtu2tbJj0hI3ctmAStsGxv7XMpOqwhxlj6xQSkuUqrzBOeAWe3S5yojZYoEVn
4W8STnGgtf4oLwq1bYmB+WVpKdn23wI53s+Rgg4qCuXkRe5CKWg4sfy9He6hqSFiaiCZwhHNc3fu
bPwyIZJx0vBURwMvKyoH0obX33dZCR0ZdxeIi0er4p2g4g5tzyA1evnEW14Z0YYZxrbk9Tmj+Rh0
RGMTiTmS0g4jPmMDfTxGAAQeefM2ZNEivrElvkcNZ9lVpVlhx63pn5YLkPwcfVd+TjrlhjpeQlg9
J5vgbBZ37ZPD3BhzYcCu4SR7brbOKYRbFvSOQbw/phgf91zUXjE+PHYyEL+hAyCiZ2ei14emA1p7
8RxlNdonmdCOdHdjc2sUfZ7ltQAHmAeNoRmXTENFgqK98df7UR2br3t+m0gIKbKrXKuuBdpNvCvI
sr+CC1gRRcFr8BZUG7I0AeL+Alh2a1CKEpeguJ42/OH2E5NM/8wlnKZH3oqXZgs45cbfZj5w2cIn
FSbk3noQ+1tZLvcT0/yE/wQbkbFq50qIbzXqdvqmbcyOewlxv5e5gGEUoagtadOAf525yc0TBaFt
nyIJouzBnGOLhVL2gCfk7AycagPAYUBnkJk3TggxhJJjPTkaUIpFfHJkQ8WySANnTG9NtMDcjiKy
Xq5xprJ89uYf+h+FVW2VY3U1krwY/2kkgjZ+MvX1KxFIJQoi6BHYJrueXcasnnrQXDkDMXNYQs5O
0QUv9t1gP9zs3TptUsSNduPhH5hbgVbYzndVSACLn0I7f2oaqG9VksUshlEg1Ojt/y42IG4vNuXv
tln0sNns0/b/meUBfMkAAUZp6x3jeLfg5YaVZJQPWnPmMxlIaeIRTOAFdkOm5GLjhEESv2ZekgSt
Z+pxs9F/QTTggY7LPzR4gK3JR5ahXgl9c7jjj/221lo0HX4KCDRKbw78pvYhk3JEpeBFfPsvNiNU
yIJdOZuZFhG8Tk3DQ3za4Y24O6/CgrmasiWI3nX8HEPCOusKojSP9RxnE4ZP1MvW9joki+pnaNd/
KzKMi1y0v0l+hmeWKNqMpk9gf6q2N5o63OFcoogsIZGD2CcZoygx/AR0p46lveqTrQf7fCMFLFca
RJyhajvpUZxB9T7mL9AgB+uoSG8MUNXs/wBAHgYSf4afNhnCm/DuOiGm0weFg/BxM4FYWlWtw/lH
q7nMGtoYIZ//OaxJZ/CJQKCNR3AR9nL68sjzHW5LFQLYZ6tvSA3tS/zYusl+dujfyEPXjzOLkZyC
Pn+k3x/mE24CXSnNxNlVPaiDpMwgBGONM5885KhZbxo2tR9vYMg3okZ/kWTBZJXpN/1pgiLRPJiy
PizNFInN4/0A06eHds93P6gjw3K7cU6uc7X8K8ZlwqYQ8p6f3gT+ibhYaJPt+9plJ3d4dY2IGIsI
sjGeNh/yYOBfQF5Eyqaq7spJhpmM//2qBSP0Lyhok3gImIvua75rxmc5wrT/VsvqOpZPJ21nEhJL
AzSJSc2RVBdvljEt3JQNMBoOAmKHxMi0N1nKlDpOshoetlJftNdHgyBJLt2Wlw8hfC+zgDPxLdCg
6puXMetRMjfN7EoDzp+7TcFmN0DAXfJtrN1kiySzfYvIsH2YLlU3pQMG85pud00Z+dcMDNJEDTr3
8EIDO1iGfHU1qb4oXXzahSllWZM+2w5XKjevDQMlX0j4bkDG6iJ2gebfpHxlunoOHUgchk+MwIOx
AW4VOZcgPyUKppowYOhYku02wcgWfnQInjec3j0yRNmppMOzQLpeW2mfgGvPKmjjcQKqq/VF35yI
ll7U1zuaNqdlDZ13y3Fs+FLNP3b67M/DSB1Qncl6QaQ+xQIwldVpwgofxzxrxCvCQv4yqXIBkTWv
s8wV8hWBIYA1VM929bZkUQKrM+mroMPQGLpatQZbXcJeSjzGp+f+/ey9oTcED8DMWYeL6YOWd24R
hZzI2RhuWVkXf3Fwp5MYdTf9OX4VlGTSey9YslsGj41TfWp8D/I3TDMrvr9X5sLzva0S2TWq7q8t
Ls+r0hSiSLBNUAtaHMlPKbtucqjfCdRr23Z5xSKjnZiZVGfNyN5ih3bezaTSmqSNJ6izekF4+ThM
qsOrjK+oEszDB0ew8SReAByIgTF55osblTPyGkUOk6d6DirpY7vvoYhft42Aeb6C/dkapIHEi/uR
6wl3/3IBHm42q7lyFzw9V/kBybNSRRCPZxfsN2BNWeGfRWxoqPzOUllQJ1jjITcu4pZ9KmXARq2d
+SMHq+7BoH5tqPg25fCuj5eIz/zOfPDSaZ80Lpky4rYzEg7+L5glLpdEv6tOw7dyzTASG3d2XFNE
sZOlpi7rVT4rG4aYRPEZlW/iIDC3qbZYekdvkgmwI3hqgQRjkY/D1VWSc5spwRfMC1Hz5Yt4lPTY
Yi6+U4wwqYmg4t2DMU1hf5ZlCAfgjmIZ/KkXjZ39Mfzt00kRMUDmD6As5sjsYtcUU4DbjvDAaRIr
hbwLI+EWd4Sce1JSHTEJG/CTrPj0wrgWHdD5HC9VoLMFI2FXCUdxLi47yZpNYHTZarx+MMG57Joz
LTgBfn/EYY5IEpmdaG5a+Ky2f1Pa9lGnWhcUAvpLSjxJDSSvclbnm4CKlkXAQ+wvjAog71e+p7FY
115Fpkic6kCLDxhcbaXea//hm3BZqL3/hbN8VPEQIHIAWOFyoh/NznihV5aE4RGWF/Z9cAiBsaKE
nzViTHgv+bOP5PjizUmrhkvkZhQf/KAnXwA53voNt0cMp73+N7UDVrAm2gX9vtx8JRqRgOO43Bd7
i3aBpHBwRPdV5WF2H8Cm5plnhzQERmYf7fZOTASWscwpHbP2Y+tE5wwh6KhgATxY5XTL/NZI414L
DhGZc36ETCZyHffcHHNSPuJk+b9i8m1G+n8r/1K+xubzKySdAUWd603NAvs8C/cklERJrPewA7Ml
MYwU60uAR0sqeiEIDJ5aSCzXjjgx+S7mFrl4cyd0wxqMhjtf+wRJ3V/3YUrQotFBt8aVkLfurZam
u442qaIlNPfj+aQUEJEDRlLDn+B/KQy5f0W+Kd+ZScJCCZgS/6nLFFJ/StjoAqkXFt1oUfS6EPTB
W/jNiMWveA3O3iN0PovSSiaxV7x1xCwvZC+ov7tGLnVwbRQGV+1Y2+pX0GXgY/cJGOwpga0vXKS8
ioahvj+bBlfEWk+ZPSsdSPqrZ8xSk4l8CnePVlalFKhX8lQI1m98btAHPKuhKC4CodmAJt4REU2U
SvyG19jIrp2GZ6qbC2Z8dpUprEN0mcYcG5fz7XXPSBcEbFN60lOrHr6AsNTM60s0prf0VGaKdmOR
sUbV4+Km4LrCqMen3cK2AYZ9kA1hyMDjs1lXanTDpHl290T1SCMR4S6UO5OmMDL4GBMoUDf7Xil7
Q43QDF8VmEjpHXmrRxYeKFlcCSvzfJmZPDohd9Q9pPCCPy4V4sJnWkRsEXe4jwF7rRSVD/yTzli+
M6X8hR/IabkmIjp4pX5NgQQ0K0e34LuT6amqqHVgDWXT1y619YGwvxDh/i0RVGd5tBXdSIUnrUDY
LjZ7X7D70T9hxLJg9k7VvfA/r8uqAq5lBMGIIBoc7isGoJ4mnydABDoZbjzrKoum/qqTtUFNaw9y
BJ3BxyCrVPCXt/zLbg6rZefNnb4rqubOr/ZAgsizmJo5M7IQh6PzPZB7sT8bgQ9SyONOohYBLPFD
cLgsLhdeSoG6cCP0TGgnMAtEgtHSpjP4m/FcgE8mtu+FMuny3C07UGduVhrc6zCz4mFEM2+jCMQx
O0nNtFzil3OVdMsnpMF/8YrRojybul9jEw6dr1A/nfow8eEGhKaCMMT8rsT0I0dksJ8TQNaem3Wq
HePXCXW5X2mhgNhS3y3EADxw8FKSHy23gNIwOzcTvxdTfrOiFN3yOyceXjySM0yZ7m1JbSu4c82z
CBAftMSPgzZ4wUuOORor2pmJKZnd3z6wTgGHJg3u6QQxsYsxmI89RkU3FHxWW2+RKateVq8HkeEe
0ne6WIKJuVp6wGOpH4PsMT/L6v5FYKrAKWmLaADC6aMZ15QJi9invJj/bNSL3qwEnI9DaZ5mPuYH
wYgukrXldfXVdJYgs4aQ0zsw4FqaVEgaupS2kyLOlYQeR1XhVPH/d7ZjRelxvIwbyvJ9cybDn8UX
8ip7bXiFRhZx9GrldzFPfxEbai+1dSHL1rj5FJJccNCUd1KPRpKfmwu1KCowngKiaRiV57JshWYr
TBxJjyBTfoymzs0EK4ZfRWNHzc4Kye6XuxigeCo8950MbtMTmESUs+P8vhjoMpr78Y2a9rHiwx+G
nNcwbk9G4WXGNTgFPK5VPh2Sbjb2koFPcvU/LgaOUUYmewCkuUnmAEvlN9btDXk2p9jf7f2Ub4CW
dQ8pqI6KoHJOaX+4ixwN4Blj4G0iGUw2dIxVYlK64PA7t64K+ZKq27NRUDeijNRTlmNRq9dz585X
CSAjJca01t/meHfu7Uw/n1BYLzHaeqJOvE3AmtqPrYTugdfsPH6l3HtaUi/IoLgDYPFCIU9x4QEs
EbkNphhE3a+PnEE3+1gHrYBz9h70GA+eBfrFOFuvuoKxmcC1a6bmU8HieQya79I0XLQXXAVMzpKo
zAws8JaLkV3e4dAvgokizgoHuarZu29mBaLEMwOgchAIeiPQeq/e8JOqV0K++BP1FjIntyR3FYJE
9YhXqFhUQ/7Zh71JPpSh0oXvIbnFzJb/UFnp4IJXoE/u7d3+ziqMtEpm7q6XJdrDE8vrPDiOhetB
spT9jy3r3ya5k+bu5t7XEapmmDxAh15RK0q9lAvFgURcqLRXtUQpeoSWb1U6WmtzEH6kOAkdzgp/
O+8yOnlzR4H69LDOMtKm5mtk4sqNuzBWS8S+NIXxNK9E16oCba1sf/mc0bw2LMlDFz+8MZIVLl/d
6P2Yb0HWl84v61CjIPS1vwQFkxDs5UGrpBwMcwfOrOED9y6BaRYA40ERbnxcAZY+bahuOKLMFgxm
djgAl+XtXIbT7FfBNsTKiMcb87LE2DDl043JjfFMAk2/dSpe4hr9hIMmsa132ajYNVw+m2VdihrJ
A0gsiEqIA2BoOsx+A2+Jkpdncbml4SfLmD7PpltFc2/c574P9evLTNujYotxN9gUaw9T2XpxTtaj
CIPRgmVB23FYLtjZzDs68umD0h3k+rFqno/BTMOpZU8NIUTO86mLyvQL6r7C+q00goZcTikQU+jy
PI4tmXiDnDbDFj6QCN/Vx+6HJIkDrf/yaNxP594Uyn6yIfswPHw/ZxpZVNs6lKCegU0rucWFcCIo
QBCZx51LGhMxfBA3XS8PBF0m37NK/P0ql2y9cyZ8EcRgUjllRFATle7Hcv+FGPN40O63IcQwRipf
bXbrZwSkyYYxe7b8wGOZc4oNobLtRJSKW6ZVCAmS2GM0UMlrDigSKDzcXdKc3YDnRpmxn2HO03/j
S20V+0UCt7iH/65IkGqm0snp4G4QUjBZaLs7FnpDApvjgzP/0Yjs5HHrTGNq9IG8/5E1YB5RO1fv
ALrkc8XitQ8P57HIq6KGH3v8ha+8B7WWbN05rysqguxqUh/6o3m9GJhH8TCy+13sDBdK6WEKcic0
gBLzmx4HYnYs3H9H0Ckh9wL4vuEJwW8mpE35PlQe4aYS51BvDi7GbXxOIg4Gf8T5KVgGUSUmbnW1
fYGrWzvTuvuebRl5Ja+TgD3bRnINh6ic4kTHpjzSDXfBPM5kiGvox+37qDOWL7vUheYcjnIyECa3
/VFahmXgsh9tYl1eF1IcdBef6Oaa8DRg/B3xctRfETYy8nboGY7qwYFbcIRWbSm/txSTRVMYIC7f
/dRe/hZOlAmBw+ba+ur0H5EOKhQCNKAkyJr6NzfyaAQGGsRMBBTHRFtP9O9rhwgB9Lw34O5nEXkE
GqM5aSUNTsr0SMrYZ5vSTDiL7ulBy0XN67r+9RLhIx11t9GMFetI5L39ylyhfOv7RlcsJ+cMUjiA
jarjxGHiKGO/i/LeoKammKPCBFv8gAIxf2cWBM7c0LZcqxzNm5qf1CZq9kDXgBAUIokIHnn+RPW2
wOQGxHQ+BkJytuxBUSt1kOCbeQoULbM0yO35bDlpYgBCCv8ZIohMM29mFakFJOpLju4vAjbjNKxv
6y2DvfqLJHzzFd1iIGCxtTyF0XJjNhwVtaXyTtm6LkJB+Ee1e3iEwN/qYmvFZSm3nk2M0X+TkTkV
0mgYC2FD/+agx9ytuz/7Bans8xt2x4T2lyFMVygCHkPstURNlUhWnxp+ZeIqVL3gP0jpuq7fS2O1
3VtUyuNMHbnHwUQKSNI1OGBiqdAFwYSH8Rk34jm/W3Fjoq1u9uYco11KR/gjAeXjzoS6qspmNhfC
1cZHjGuvHLAY9VdNXE49/yK25TdGOJeBfa3zrlZYt5rXPeC+NKDJ3XQ1L4NjnpccVAgRtH7Ob5iT
ihX/1yQaT0sHNHzNb//AwBIyzjXli9i4vMSssxPqvbFqp+N9jCNOaY6ZCoculjHOsbAmsPJBvlvw
yRWBfZG+vVOm6dPTnI5fnkroy0Sb+8JXUxqi+5iBcivl6dG8Nf3cz5VHMSfo7S3yHTFsl8KfYlHO
Yk5wR+dZWXSNtmcNZIYhRcz1x2a+oqNojo/yGIvr99WGyVwbsFQvomFss0kG/MjEEQhXmBXavk5d
Is7wHQHjDlMZ3UFtymUt03SYBEa5sBRGBO1K1p7DQrJRpCPwab+Lonc/PlcX/pUqtkGhCIpfSQtY
gf6mXwXj2jQ6T4T1LO3oRXGIMtrKMsO8sTj5VQKIYXnn/1LNwusatkjsGYBGrVV20g8K6TTgr6gq
HjHCMiEcCJD2E45lKomFrYsdA4R/0PwRb5hEe6lXkQ7Y9CNmoEKu6XvQFffeoKbDRqj7pnNL2I4R
TdVcNDCBjJrOD1O+F47YamIzEyq/XxebJv18Hf6XJ3+SYIc/tOKqgb2/Fgozm2yoOeftGKaeCzBG
YnoZmQ+s2oX+DJrgVHfEIgs9uaNGW/FWNjdQDbI22MGuBexRGjLM5OxIumd+7/Z5Pt04RZycUPhb
38U/gKiJIu/yk15u2/qoE8cLWJ+vmxkbnF+xJnf/zna4CNPD7Vnpudf5yXhBsFiWtxV14VG6gX3v
l9++Cbbq/OBTM/UAuIhZ7886AAq1TZw1m51E5L1FhqvYVhSzDp3h8p74kHZuCMCVbOzN/CyHP6Je
kDJeJ6Nd7XZf5vw+VCVy4XfnWRPikEl8veGI833WbIEUB8d5FmkrwoEbFEvGiXYcSsmBY/j6266b
d/PCIX5nD6NAGKCnAl9QXgvvkZa7EzXvuugi8S1Gkd0T+sulCcIere62M+JI01RSNdAma2vUajpj
FEtHxvxakdczhhDMJY+OrUarsVoOncZJtPzrA8VlCioMZb0oF7J787uCUENwUQ61XCCMD6bIyvIY
a72aROD+pmISO8Y8CtMjXhD46450pjxVfSI6morTmBNksJKvDS+5uDH5gnlN9P3kEQX2z3LWHc6C
sauwETNrNLdOuJOxLdtEhWbNXBJ29NERDwJlsX65otZCV4jrQzlLlBL2Vv2ihKSOHDe4bksjqNie
f15geWZqVT/wKBO/mtyTrd8SWlR9kU/E3HcD0D2+gYsiNtkhGgHUoTGFlmFmyMsKsPoQCWxwqebJ
oP4ENUCU/phGW+O4bPHq8ZsP4YJcZ+eNaanX3ksjIFhUQ4zLZXDCER1WRwqC/jki5NS7/tleDtgt
jA2gD9GFY/5Wq2AemPuj5qYTV2hnlzJXAsPTDTPjWFrNlHdELklmUvF822Yd/5wIYazw3DzKtoAZ
tEWE2jpv0TETivqIlrWsVJBYvjK6nM2BxEyiIBTSZYhojCqro4x0FwdMC3kVs9uERcK6Mitxp1uV
ABM58DiblDBt/9gUujY6Ku2sgHB9g6N8qsjXJv1cOlpPrUKFW8LzGUsaCBQytmm4AssqqRBIMFNk
R7YZvAOXxrN94u+M5gH/4JhiaQLC+of3nF0xokES93X6dPVRGnywuGdXKa0uN57ltjZrC8Gymm4r
pweYQrOYUbiYFyGeKKtDDWgo5S1RtpLjKokaq1a94VXWHUUcZvXMBEb3ZaOTJkbtJiutcq04EIWl
diwGu9VfJyjyYl1QEU5XwuTywCoEe4MiQSBDZBSd4ym+L6MuXO2iyUOZ49G4zjSYLA7k+x8KYacH
zQOK2MWid/6ZxvJLUXR7Oe3WF9yo4YINobldfI+IBwRuakV7bnZW7JpanhF5Qj1jVDD/KhlnatvL
44LnY25ZFBDBQaKEzcwTw2gLW6BRuNwLUdT8i+m+XyLEC31mpo4ywUrN3DO4O3X4HuqIBD/Bz2MD
dO6po65qvzT8fy68ksHoi6aP3aTa6ZeWDHgdVbpzoOigc+YBMUbzzcCMfhtljSthKWUDVJEBMj4Q
QhzqsRzVkOhbrV9FPBH0j0BRyhIXM+HBUPhUcXOZhUJhzG+lYUE0HsLhWARV9ectKGiHCAoB1Jqt
WWtmdS2GxGMtWVTb/B3nokKSMmN5TNqnDVCLORcV1vVpZSt1/2jPsJFu/bPbc5io8MNVZqaCKrSL
ncVZBLv4+ECDZi6xwRnEywvBnqJwoNCi7ce6s4ecLkDsldU8SW+wefxywrHyMvyHeqUpbkBoufxd
W0tXRfCwZSCL9C3SsaBD2bZz4bmyWWElWRG5e1/DQaJncFvBYZmDlVjXDmE1uXpoBoMwJ0Srdq2B
iNc0zfrPJ+ssnt+WvrtAg6CiZyMnE23bLTATKp02U6A0Wq5HYBj8ZLdbTfvKpX47BUiKSEg0b7zw
sb6sZJ8QBNJZ7W8ooeAkTqChitolcZI4pk2rQIdnA2RjrVqB5KJsgb3cA6nMKygZNEmOWNBmnwoO
bAmLexGXe1mR4CRnPBKjBYa5E1UHs1C++QpfQ+Zygk75hvRDSSATnjd5AquVhPWNhF619bm1mSx7
l4YFpTREuAokNXqp88qjIDu5HIV5G2PTbo5bRhp4vIIj29ZBL7oDE76MSP8uPqnm1Fn0PVpsA94y
ut6SFl9imhZmkLQeVcFmCS08Mq/5+XQaMI1ebErXEFX/eK17QXEctSwCvKZvON+DHjEkeFvqzXO/
upY7/0rJsbsBgzcYpETFVkE3j45SumgV2RvdqqSAp15Vmi8eAhJ65ncSYqKsPsv3mV/OFLmhcqFr
bMKnOoGw00eWP4DXAJtmx2ev+wm7gYSzeb9iLcl2tkjzhoZwxXjFy9ubK4ybtr3x6g4g6VsIo1sK
9YGDjUfQM7cBT+Ggz9b07l8xutlLDBCYMWSlTVA0rBg6/GGQGQdJ+2ZUpjqxBCGr389wbthQcY+Y
4biQX/zSc8jkfBnrvWpWCdFRM2CTs11A1mvvXbuTL1JxPqtjSuZoAuptkHntZUUFJ5PM0U3dTZpa
EJdihGax2M3dJN2jQ2/kbIsIQRT7C3QNp3m0AfC9/mBhDAKvM6q7g+cP6FRUNDPpl/SrKQTOSB+X
ZMdOTRCC8ARESFslWnL3HQDokXpFZeDzWYmeti5pAtQcb8Z25I+WHTz1ySnstYgevd7k5MGQmmRf
/QWXA7UfSfKRWnxGCoVjfRD75mZfFUow/pgJJWtQtW2hA0TVWIgd5dK1lEP6FLN3euBc43mwOTdf
6smr/9fyY4ym4GST4/9xB0ZRn9RQX+XR5tOLZCJChSS4NbFZ/msDVl8hoKylGj482dpE3pEAYmKB
xiLlLO4ZEyiHmHH1oc8MJMjaJQvB4uK10/ara9c+CgZEO4UpwIGyXvZ4GqT4cTEX5LMxQLdm2Eqy
jkcNpkwFdtiE2eXmduSqLGk9IapSwmDczHGs1/5/MiblH+UoGNIx44wOtNSHpr8/s1S4tVb6N/l6
HvxftjnNGxvXPKaN/HXwA+SZzludDZwb1PXbcP+S2fyGVEhaJSrej7rT8uMk4+0qb5HxnZtPMfAs
sXOTUDmo2YzcdHzxWqow8wZ91mGTE/41YQ8aDPABjrciSqYLHUnGZNGp65/6tQbmXiQQdNOCc3Tr
oEV+E0EVMWEpuHbnSwRXYHM30iW0A15JP+GKsi4CZS8M3ph/Gk4r6JvTkcJejFVWtyhEv7uO69hv
Kiw6RaqnadqXqrm0hTQUPYTSjzvd9FeN1fuXY8JsMTrzwMoinFqgzC69QPeErMuVtx07Bh0Tk2w0
57espIR9iGdcENJQVxJMyI+JNmsEhZK6GQJfV3aVqFwuKBrJm1sVxe7RvkVduF16nR/qf9pMJ6Dw
fIXlSZOPzytqSHTayqTxjMYPI4tI11MoODhyY/wuuD+vYKpvdEsYlPLYuJBch8BiUn0LLZAw5qoE
4ytT7J6NjhnNrxu9flUSkYmZR8AjBeXFXEOvWR4Q0EsHbzcV2ZABqfRZxzlT0qYjuo7fsOoI07wh
8UowlSWR7BOgQP4PC8XVrN8CFD9ek9823q4vaaGORgpUN7/4rImJ4L0X5GCD17YeBvaxc1LykMIf
uXwKx6KYc/1zHQY8oifMoQBg/zU4B8YMHsd3c0xp+JnXTFVuamW9Oy1yz1FQBMprPqSW+co//Wjb
9Qt/yO5im/+rQQ8Ae8womvAlWBogHXuZpj/jnfaV2Nt03EokeWXJCJH7P5ykVE2XGZNsM7/3OHOC
iFWEPZrW8+7oc3X34s2R4fVHMCWcCLWa/ZuXFyzB82hj/wjPOIVJJ7MoYl00bY5Vv+5jCL8yr5ni
+0vr0gIAWLkEs5VCGy/fYoPIO/BvcuaSXNrrSAQVhr4mzJRRlJWPv8jVlugj4XOxYku1psDDZVED
n1REMEXLWRfzjEICXObiGhuMIiHO2PA2Lph4dN7RQZXPhafElIX2RXXodbNp6VjTUARlYqw/w9+x
8f7e4FFkSU5LdOia/rw3vwDpQDTrfXuV0yD+0XE3C8+phEmSvxtgAOQIgIIXx3By2qQbDoXUbmqR
GVwXQbecDV4LoWb2mTAb3YMJAIkcJv8KU4nVZevhesfjng7sRcJIrVYfiWynHm4VmhheLjGyi2S6
42M0K/wv83aRlIbqME++CcLcRoCBFfrt2JFaXOVK6biCwbasRkL2Fj6s2EAnOjaKxlJK74rdWjlk
4LAVusxdYP8a05s9HYB0ZPiUPenXwPsJSrE2XDiyiR8RmsfO4fRyPvWXhFe0EtXhRLupUZH6ma18
m1HiBCnNGh4AvDz5Ymem2aTX0qJ+WCSMHWm2U0BpAwYjT+A/1voe6gPwTcIPuz9UFFR+zuNSol2k
8EZ10YILKL4PdNCyoHrq1BOFwpGG+ULuoTTM5u9okqpj3TxtvjwvQMMSAEWi1lKkQ5TRaiUC5AQ/
v+YNrjbdpeUNa4ElEKVpZRqeX5XHsdqJ9e+o1yawPD2XQr6o26TYuGZtl+YyB9WuVGsDre3/8nb1
GYmLQ7uaH3jK/KMnU44PgickXRUhj/z3kxbQ+SH7YnYooUAR7v80o929uHvtN6heq+B8QT2RYROA
Zoa5C/WVl27EgT5NytzH+aiyZGVp6nPngqQLogg56B0J/glHRtx2GZps9m9kHdsXgLY1QyAuegSe
J08Wil6D9N45VM6GxZRstU+nGNiVFMaQFgSrwTnoSnmuXHSvfPUMjMlmt6osrN+JYvLb0yO7FRx5
lu44VY5NW2JZZi59Zg56QJrB3V8rxoA2JksnsCnctVBBu02Y5lvgsvI71f5Gs0NGJSdab+ps2OTg
Td/N1dwTH3+HnabbpouO2dPjhjPljHWo6FHWfPD/WtdZJN2SJjcfZs6gJk3CWt4j9zbvDnp0520i
QBbx+Va+7ubXPHi+4OAUXAVeNiUZyk7vzm7r3WhcnTdQPlKTBXEhFf9vNvFI5E0I26Hx1zfPSzMX
q9q7OJrSDyxtjp5hCZ0dkgFrYBTHvi+JHthrFdoqe9Gb1H9W8HucQGTu/DNiTZVgEpBXAFCeKnEZ
kd24fh7kVF0HfU5KatcQ0DvCqJVaRWbVttdU5hcB92028oaFGWoEcJG+WmnywEsERzLsj0oAL42P
TyTkHSdEYENdFP/i7M8hPAS6zHEGSLYkg+5p9q7OpMRrkQp6ioQcslIEu7XJ6VKp1+FFEelvWPyi
vpyLoUP6chtb9PmR5PGI2yzNu0BY59mqNfmg8dOQrEgR6lG4ALClp9qVNQFe8ODuq0daGduuaBQs
GJLY2ImgSyjIXyGI3lga8+3+xDsGUgir0mtGv/qH11jTTu0DQa8L2rKqoUfh6YDY9isvbFeBPGIq
YwQMbp10NvkpuMxM/+gCp19AygFZ9modyFuIboJtzfYas2JmQunc9IavPWxeUVlGFws/+Maak+dm
URGGAbH40H5XwRs9zK68FAlW3ODlDJqZVYuBreiTCjI22FPg1R+lBIVf8osXwu7v7fnRucSzOj3d
cyYpAVJ62V81a1K0ZJfkOGB6EUQy0Bq4QEx5mjmVsLbmXlsXFuZ74ExAEJagN9Zk1MXi5J/6OGo5
/Sc8nUnFUoDXxtM1w8iwFbcqr4xXbpGZ7xfAGEBE1zfJDUI2KnYdlauGcSdXDpIuli8xtTGWOIdc
E81QB90gFE5mbdHlFz0pTQvEUFHfwrgVnyVYE92tPd0gRBg7GwZ7hdGyRplLTKKk+pDghsWjDATy
uavYuaDtBTvfyR+qAAssjtga5UQogEXnB++n91ZDD+oBQbtijfHEzxKdDo1zmutPojW6RrKdIFqg
vyR404odVdIiVg/rQh6alugYYcMz1ocNUTKPiOV58Ns3wWnPLf/76U7BWlMp9ClJncYjl2tJu9o6
fWxC9NVY7f8OgRa1WX2KJH62xy+Wa5O6YebIM4vOVwphq9oqgw6O2JvkgHJ13D+WiTA0vJb4mg0K
I4F6ZXB35qXhUtDIUPUjzuYSBiml+XBrencCsfs/2raOEtka5KP4gMW8+BxR579nWbWRbpRGsZY1
LPSCahnqqwNNUoAzzlnYpi2ebHowdxvBADtiBVDBjgvkDuOarqBKE5YirtVLNkLCNtT3WLzDeSZ8
5yJ84m+MEEBE55k/SFa6OCVnkaXa0UUrtnnrMgYNs9PfveI1pvPKY0pTFyAzRfdkMMuU2QwE3110
DDZ+Tjd2iN+7ClWDoZZHAIhR2pUXGwSU0PdLoOHyVzKFdRtxJbqvrlZuvlMLiDG/yIWgO5P9M3N4
+DyVwLudUpSxXTT0zWpTzIm2eutezC3e1moXck6+HLc3qoNd/oHt+Jcatu+R/uK2ECkbg4ZPqilq
V0Mv9f8ntjmY03nP+yltU7Lu7fQHpvVRqfCJq0gSaEMvcDMCFYXqivET1jdFgKAynm5/45lP2NXv
vOrzE0FfcFzkRCoexkWN+72klaLZEZGiNT5/GMfhl3cObNYZ9MUp2ify4N+s3G5C0ZuvUc2c4+qO
ca0JzLFC611/7/SZ8qSuOSOoc3TRgMu9boiAEca1rS1WQ/NXeEiKcD4dHn8AimyahX4zQcoZs/Z4
TUy2TrO5EMxFnYpc6otncPlCNUSkL/juQhHHSNZ5OD9ow/3NdqDAdT/e57ioOZr8G+JJeBS+37Mi
8fBNAM2r1JBazU2UqQchOUN6kt6VFL2uuSEazpvEi58CchauzM5xMAg7/qx/7eG9rRUTZ5j8giND
l9jiLjjOsd4higisQ0Rd/YebrXFoh53nD6YRI1s5PlhRBXUkOUntJdZvtiN7atrUxggHDZt+Im/P
kPz6VJeMx8hN1lueoscXlWHx7OSlXuOLDebgMrR6h/mZbDymF+2Hw9EJfE+YnrXcmDzHdP7WzYn2
wQ9zG/wGvkTYHB6Y+7k+1eeUmNb/dQkkgfFZYuaDBtxkq9a/IdJXnKu2WW1k4LcqiEa19L4KkUNF
ykCHdgSO70vVOShf1HREHzyt5RCXLqcnbSkaGc/vXXCJmEJOIQNJwCoKtgb7WoXoOFTG+Ox64qxp
ukWHqWTvik2etjVIZPkxN/0/NCRVRRVmRgV8vWN9Wanqigi9OBAIiU2cZBTFkp9YyNqJqB+Gwo3o
BkTwSvZ4Oa4Uvnqj6h/1ohH/WiwaoPvYMfLO5/xtEDy2mpFoME6+RqnVcp6d4q0JW0hJ2MWbGrqS
cXpEEeQaWRnszhFyu/jhIcj9unF8z47BrZV3Ix8w8iFJ1klLs4ILvOwN/2ZUkeypRoep9etMzrh3
F+j5XZGbqvWrfvrmj38pQamcwBkX3KRGwsRvmYxnKa+YcBEzJoqyzSNZVRqM4+HgUlJkWs6ihjHW
vFagu5YN3u1ssrB/W1hq8fmyRLKrG5Y+Uat+9iZEzB5C3J8QQZeKt4d0GHq6iSQXWKTRSIUJLVRZ
tezXP1n5RJDSuXS7SwnOYh/DUwflXOsUCps2B2gR+AvEBsoYWIKdX+FKPb+sagS2IzAUTMqjm8pv
7dKtolgofqI37zBiEzv3xV9MIY32tj9AorqPE1fMfX139t3aAXL6zHqzOwL3Gy6JIZocI/8VOqFS
e68Q/LwmE6DeYVKvsozFNYVkeMGe0aNi4plucklnmKQSf63V70Jh/rJZ7Rqa9Hg3q95kao5OZOif
gVscGs9zRwmAvUvZSi70LJgeNtUtTMfVcxhfhDrwG1kWRfPg3hZBZlQYYBuQNtcigw3TSRnwT7c1
OwNRVNLOsFwJiKo4bX1ZUUmb8rfI5O++Emg4WJCyGt9gcIVtS869DPWbLSRF8vkenheFl9nbnbpL
DJ3F3CPUFSsEMOOkWxjfomlZcI3wGb4XkduViFqmzNTbnyuUG5k45Bqf9uNGL6xRRVxRZke65U6E
aifLqk/NclG/ZqV8XzMSEPlIIu1gpsxYwIQfxOEsZs7bWLmQhjD8i7gCjrhPWqTSxzfBNaxc2TVv
96bPBemqRn56klDP64pYoqq+h4FtvnXdKlUwsV+j/r+evk48BC/5JndduDCfIfmUvRh9lRb1CqcG
sWocU6UwUjQJsL5vz44b9Uh6bPhmQi5uYcTGOn7gg/p1Hxcqd3RcsKKJ1wFdk4XXRIiURqMUO7+O
b7aVov+VuE9FH6SVYLj2ltpOJtnU137xLj0t1HinLD4rIORQ36iq8DujEuLuszdvROajwiNn3bjX
HEHbFPMLx2A96f7ouvi5ykHHx8k9NhMPumY2HDxvdeX0I6dGccanj7CyO1w+qRgFZkEh8d3u9ZvK
jZ5sg3K8fwzAS3xBKKvUiJnGL+89+O8apcdfdCKj8Ok97Ndp9pN/0dcbHSRJCNutwsAZOC4xkoDJ
VGVS12o5YEBtl7UJZfo2ecvA5blH+0kEe4GwjX2U3YaRu48TfeGMlZ3Iqs3P5neUXwZAUg/36sKt
BTwC3n2v6VOjphLN+yaz6rUAjTXU+uuRuGdNVVPlCUjbOHIrnjfTX7xuBF3V+wCTqrZ30gaLXkVt
BnpIE9Llneei3qsaUPMlNonPW55W1vUOu565TmS6ecPfQs4ZLje4nHhAOAxAbsUlZptfQWpvhOJk
ZhqfTwN52D9yCFFZnIV5mFNMAw/DRdH3ssncjdPjAC9as6ntbKxaJcviyaGeO15EWyXHY1w8TKMp
NlAFU35cLX4utnCwO/lFlUz51P5uj3HSY1hWQ7hQrTD5yFx4nVK207v1l956kAImxMtpdBDyQspl
2GriXPOylhbzjOh2gjBUyrjSDgYy+5W2OsuHhe96LdrjByxfb6q0ZTkmEWeDUG83BYFzBE7EmuUi
gEK27BOWzJYJ2D4YzhacAEu1UYgxkM/TiQni9C+fqFhiqTO6kNeaM0ZhPUXh0Kg+ZufZ0M6lgewH
RFHNvxZZw39zctGG8Daijd7DAcUXuw2ybocpPHW6c9lc8FR0oAtlZ0V1Et5qbCr0VI3cjzxACHN2
jMyecFG2730c3c0vNIbd9/uZybUUuW+qfjGG2SnYn++06gA3/TRbC3MaNJjYglOGFfc1eAiFLWpX
mn1W241mIgUgtNm3YRoufs8BGj+oFTHqWwbxWbWrPISr1yDpzZjEFKdWl1cooxMs7fjW7xfTXGTX
orF9lVU01rD1EESB7ZGBii6pDo/ldQmTL6JG9w2NfSHKMOHxN96SKtneBNMZXxn4wFq6Lnzr+4fh
ReDlvq2YIEgIgUaVq0neFCxx+TwFXOQlNK/gGbDsvFPp+STNph6NKMp0ButBwbwpscXLa7FwAbJ+
YVLKJKT3NnQIivSKufYKn3Z5bvHvz28TYeZi2ustAasTgACk6UhfceImgFRFnkQsyhFDUsO2U5zp
Jy8yqgFEQdrln3QQUugtHX9W3ZWOo6z/M8D/diikZkyaJIF5ppraxjkqLlNEusxZFAyOuExq2QQN
b5p07GMlMMQj+3xRaeDj4xdH6VOfU3CWjWrghdzWuvDvoXZDb5PJiZsfbO3jRhUyS1pc7arcr6Nk
vB76YIhIs8lcrsZWcu7lGZj3CBh3NOIeDpMSlTTs6y25Fza41pzuZKx3vtectbyb0a8BYNKz671r
/i/Er0CdwFuMHivl0QABU+apBEv7RqpalRqEz7JBV42AZ72u0blL23VSMY5QaT4oYCy3/5+Cc55H
vM4cMXeOVynXDaGMYrQAY7XNlKtdD48KmQNJVlwyzshl7DZOnvFgYWVvFG+RqQyOWCAxpG4QRJlk
LHeKt9VEdT9IATLydRK/WyXzLdIbpVZutLUr+FRos1mmoPlBHQ9RUmF9koc46bfqHbjM9he5Eu3I
zLio39WyZJ06m/KkSXErluSq7zn5CkRqe84wEtldl/hiXDKo3oCkP2CkIcwX9xj18UA0y3lAkxW0
a+QkygHdKo/cr8hwi8nVo/xgrZWmfhHtlVW5VVwAMqBUdH63yShsmfiOHBAqRYHzn//bz+nW+BoC
UOQq7O3f37T69CLj6WZ9nx8W7EDOUWg8LCoVEOQu5liHdrVD8abBCMSeiqO4N4HgEwR2EkFS3sGp
0tajNrz+U6ZD5xHZitV2aZm6QMWMObBVOeAcMSNaBG/w631BdPBQznqxF9wOr4D0/GxVyuSxxj+K
VJVdcV8rHl1OfmfbviV5fZfCHvoprvilbhMojYZWh+VQ2BvcNaxhCxYn2NgABYqhVghk0d5vR2YX
pjMjBRKsCfiE7eaaMJMheuuRNP6YOe/z7919qPwsBSptmmg5wujfJX/X/QkjHbysz0erUGgDNVvg
NIW9biklfTGdmDSYGpelujQ0MfkOLa8y+8SJWpjPd7GA4W/NZplwKO381lAY3LRVxuC/Tr8icl31
pyRfGUQBGIAldFymX9qLxvQShkgilXZT7gkU70pI+dumq9zmezEEH0kSeWVm2+1AWA4DD/AJzN3t
MK0BH9GUlA04fraKVGL3cbZdfAMlhZEtyjwfH8LdBMkejfsZZx0RKhm8vVf37GIEeQCGswp/PbDM
MqMzWkCHd7mCapl+LXSaLDCm6Xd9rAfgpiMLHHlzl03XBJLsQxA+j7Pnhp9WdFIntD5xhg6L07Pf
i4QYeOWAq5JeyzqsMcit9BCbwOWGf4Ziib+66RYMYHg62LyQ71hF2UQQvbstIbr8/Rtnz2mqj2sl
ZEi5z8BhKM9VxxW74KqQOezdM4YLFAejV4H3Rz5cll6+1QzHPtdFREOOzn4At3gVn17wuKuxEa+A
uyzG9EEh63L2VeZ8pZun7DkA5kDOwo9BIp6U8Lg4mAIxdBkIBTrcLH1AVTL+fPFHyRcdIIEJ3hMZ
MO2o61TJzWHghmqbkw8IPGZEhbPYbcuL1p1cwA+BnsyNBAz1gHrnwzzxgyon7EXjLSfy+T8N5Mnn
qq5gmEGXqpYGNquXFjq9YcNjOw1WAXjVTSiqSLAQU1oAbp2uNhuaDw6eVZXi8glxUI+drvv8v+Qv
66MqzjqPEbk68f0Sl0q9uD18nndKVaMs43lEP4uTl7nYnQM9N40egsiB/1sbUdhkS/NiH8Uwj70p
tMlcXPfovF3n8xCHcYHCtlzGsJqX5Uwh2CozF6Ho2xRAbBKMfpbY4+Afbu5xSShgWy2wQncAlYnB
Dbak3Vp0Mh5dEQA7L9dogqT76X4WhH41sh8Tdf8Y6yS6VROH/zhMSa0dnxxjHfcd8xd7qzswDgJZ
PQXJTygME3QvcMsUykSclb4hMv7AvcU/BiSQC9yeW1AAcptuI/3xiQCzpAXJYJoOp1rxa0cmBCpu
xiljRe7q3NiYZiK+sJvlrW591vEasHpPsnuqpc61oP9Ry35uo/1Rzc3uSrK1oRynTJtEBm/llYu2
QCEf0z1n19qJeYKt9vQbW8YVpEdOLU1K606mGrxIbd1jqwrdy0CQYzBOT9830PvYlq05AWv9H/HR
5ZnnGbLLBXT4qPeRH8FvYI/fEgQuuYryMZYjBJC0PgZ7vfWHGgPMg3V33zRpFj/yIuVGAO0Uyyeb
/SzoC0YYG67ZRlmSDpxXDsebmJXHSUS4xE42MJQkf0gGG9igbGTsTu6wJ8S3GfzJOHGu/P7MXAvH
RksSGpKHK1Sg1slxLqyR9XQjJXzvLNLy6O4mbbRX07M0UInrRmKIreius9yYx0p4L9U+WnsaaDhA
O7RKqy5D6mUzX1Zr02NmIC2CriaWpYtkCZuyLU+IhUr0w97aVbhZ09GbBH6A4HyRU/bQer9IzLNL
gnrJ6vvxDs4BlIO5YV9ePeoePLWJ8Wop8UDEfWFd64cgbnG0zmX+hIFNQdiP9Tbx25W85gwq3IvH
rFLEWwqHf5BKQhBFQ07d874kEEnOgp2O/WztYMDkqCC+pyGQ/H4eBwBvQ06axOzbLCRU756x7cfw
MODHdWz1QYBbT9LrHmLG0Y2g2lCo/IOlRiQKjIt8wbI4XPLYFLbtJVCSdOELKCkw0V9WP3m6wFKc
qqmG5MLJ5m+gTiIjER0OqxVY0pp7YxfMznveVTuA9MWSkeH9HOTLOIp+Ax2osrn5ElYQqdO9WXy8
owVCUJFsnyZxoK7MQOF1WoqP5lFwdml7c4M+JcICJowsOTGuoxQPPlK97lShDjclFRNza3aNygjQ
9eB4Nm7WFQIvjXOpBxHBTipgqcN/mwSRQcWPChIZq0C/oFOfvbeWQgxxs36dirfcVk0vkRaEV4D9
L7t0T/zJzLx2P2rVDiHwptINASqS+iRT89qTkLExSeY42BShU7wn+VNfHUiveD1kIGBn9iVoRnzy
Mroe5MWCPuNQ+KIKmYlIMTSbKa20NJ75HHzuL0sfeSfV5z+2JTlGezP8zh/ed+db2dBY/JXOs0Fx
le0qLjPSj21OBcBvA2dOHSsquAdX27/jld4XMppGEv/fQoRznUvo+c/JrRhTh3xR+nj0OMROfQDm
LhLJS8suA/6AR/qnngQdQtyMKSWNNvv1/CHRtUEn+2O7fq47edN8lxH113yLwZ+KvGH5Z/Wnf4Mb
bfY2XoWO7k++ddfRN3OtidMde5q+rMX4tRgqgWD4jNpClv4oMVbZ2yAYGdnExFo/zxZYjGvGTVkJ
pdkbYnQsj7UEs1q6/VwcIIT49oqjNyEEFso9aMV8Z1KxOUD/r3iUVC29kfpktk89h+mTe0Js3YCM
ZN3aet1avQkYnVTbEDxlf0sjVkOVI4nkRZ3/NZ01kqVLnrU8oH71mPB15cE0wI1Ow/PPWU/7IjfJ
5AZMhn5uACZU0oPIBUNtXN3KvrLrLcPqXiptJzAcgki38kUOqVad6eTAd1Je4SgTR+ZpSKDGphiT
LjAf2ht/hUPjGSrOZVwVrndB9tFUSQ72Rth7EfQ9kO00QlaW548tNqTYwpKnmnyhQkwTbOArnSDz
WKR2LPQ1LYg0f/C+0y0CGTlS2CpZwnGb2T00waeKZmP22FV2j/ES6JM4iZNYS9K2PBFSnOwt1+fl
4VSj3+D4BH+YSSihRBRMlE0u7f5/gAnspuyPmLOwgnrr11mIqBiccJw+hkU0SUh1k7c1oQBhfopN
9gyLvpjLefGMRIks3xVHWpeOpAF/8LcNtWAvav4q+CvygW6vkIMGUT1GBaexFwd69sf6e4iEjxSu
Uy9it3ywos1yRvL//lYG7R+e3R7voReZ9A2dLudK4Ww7GzLnBSYIMDQzp9gU2GzM+kVxdNdEpUwU
SR50aC3FhIy1UrNwGWPw+2n6dWKa7Bidp5+ea4+FbZGIp+tdNsDabJx46lUzfAaFPQOtublHYVaV
T/fE2Pf/HRbXBXjBjfrSgYSd+qHAIQt16cxBWmePiAoFA21KYxaDC8PN9/aQX4wGnvy8vhl9+wLE
e1U+yGsYysxRn/AXTPrHNzexx+JiyOVV+58Xpz31C7eJ1GydRtyLdzQNgYhymV2aj96IVloZnHWX
t0VU5CCsYHNBSGfFauaztW9mP8kFwM7sbN+fH34FHAfyUBA5RJTEBo3aON4UxcVk2IhVD9uRPllC
FVQJc3RkA634jXlO7/r1vHnPt1+DqlvjDNoz9YDFthmd41PPuKNNLiZOsztru+JrJwBNLJrMHLJC
csOWz1Jek/2g3/hMcDMaPFNaWKV6pBDKRj7pGhqu2ARYG+ARE8Uc4eyTg9ODfXwSWBcfUyQ3ahcr
C7QPNtBvmzOB88VXFanPfysxk0uiF2i77usxsQs1C2zpguDnICXj6+N8q6YhTaZVPGLpgM2eR9vu
wf9uTboXqg+Z3LgICFELVHLVKPel8hinw2aQOgtv6dIO+2fw7HUum78VjyVo8tzmgYJdrLFMoWWA
M+YEIIWECsyGUj/w9oMioV3etPrNOMknF6vv/iqADJdNNfsygI4VPMHYVDpDY+9s2TRQAdR26bZQ
RsXNZN6LAwFPubV5Q+IL03DaonAhKCd+zTNWVA1WJUBa8IL5FadTj4mDcROVL0MJd39kWAcob57R
31sDvB0I9yPui2m+8tbwQOBv25Gp9rFPF26Wl2l9A4IwwyuzC+xlr/WCzpI8hqV3KbOyr9Ne66GX
G0P+hpRTDd1yn888xtcwIV/WT1yJoGN2/C3XNlfEASTtDtTqerVx5IxVtrL3fekEy9ifSkGA3aPV
RCSMynmWM3KB7KnbHvYGkiE61bba+CIKRtYuKQNDBmwj7TzmykQ59ssXPi7M2S53FyhvS9VT9CF9
GRrW+dls0aHnJT9GIqiOIZIbpAFW2vMv03iTNYyPr38EG4VetohTd+9ACeTtigfMD1Dzh0NSpp51
hzQ30GpdLpoAr4rBe28BRnHDrz1+HS7Ct5oDD/2r/AbZbh+P0viJegvKz/F3PEzdWu/ZLS3VUM56
dmHYpR/h/EnfaCxwBU8jtCLl/uAQmrCCKhnrTZ43C1wK+YQC0VnDv4sNV8Vyo8GZslJj0Q==
`protect end_protected
