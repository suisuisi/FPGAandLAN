`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RopYFctZpOGKOvn7RsciU6+/8clWn0fLqM2ciHsoXHboWiCwtWV1HacodlAF4c/EeutjnFuuKf+e
BOUzM5LykQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hEpfu93c1owsglRxrpVUo8cP71+Ijqox6+nIxRg9+JC809EcNvYGuHI3R1YTVG1CWcghWx48fTum
s3F6tnwvF+5mAofn6TKff7dEvpo162cG2ZnYfl1lCuuJ/M04EL8X8f+7lQqZdROKMvjtD+4giupU
f0vwCaVOeGL6TkvuenA=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q/HcacaLLjlaZB/BInJxY1rPWl3qAjAmt8yeaqKSpbQvy9p3gOU5dlyepcBTTPEmJ57U7mu9s8ep
/fXuqlUoDM1RZT+zc9F8YLgoZ3p1kt2W9Rluk+CHtBRsk6yvLFv8GqJm8HL7r5O5Oudk/pb47fRM
QhvGa23VK6zKBwE6HCM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HY6sK5KbNAaVu5j5JnxQmzYdaXT/ZNey1CF93PRyG6NOxcnttuHskrg/EbaO9bbIObzbjae2vDDA
CAH7Hb/qVGv/CZjSzz76gMRlJADwY28yP5fc414ezgCW6Ddhpr+e7HmWr22EvozSBPDhNQJxK34T
P4jGYLax2yoEwM87Lc/ptosGV/5vngZeiB4pmGgyeDcBcN6HvIv3IMiLBWvbExPzWdSR8byd1HNn
WkdqWKTerJSXG8zXHp/5m/i7afkLIjztHYtZa2i02OO3nCDt5ddwBkl20T60iNrfwq/KsHlbxmYA
S2lSJBrIVJnaJI6MQTCuxuoRQ48tJanzQ6MaIw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mL3RKXswakw4gob1//loEP/FnJbpyuu/Rs1zoL3ywf/YLHH9FJ+qfkCAHgPX4p9He/3VFOUKtUYz
qWr5QVI+jW56Kg3eVUgzMADNlgufsbeOS7KrRO/YfVCen/n6kcd+nfQKfEO/XSyhycf5iVbm2ko7
jVar+Ek7RVKu2xZv0uAwfI2qOStSsVwe9/zhvoqVUdQBhzpnV7BzFNZ3SNKr4wg7/uKE2Ll9OBQt
H/fG+Ed2LPwZRgz4gbpvnWfUceTZMC8f8dUZObkARzc0Z2A9encr8Xag8F+pefyUrqbu4e5su1a9
A2Htia74sHqVJvEhdj5GByml8XA7LMT3rE7oKw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SKnnZmDU4XvTt1KUZLATj8pfSygo0T35TZZ7OOCqFuA7eTGVwofl5+JFFFp/ysTkqwvxsJ5dHyYI
ubG5DnTdPLnaYgNioP4mPJUZxRWaOykLvKRMQeHvhqUIl8A5D8eqDC6qi2naRjyw6Ml62RSI/bP3
2xd4Sl2MU5+U/77pL0cS9baXI/WDaDpq8emDzNev6+MEjlMxZhZcBVSz6CiCC/nM+XIk/aKa/6IJ
1iYFCS7Dkqyro12a4hRMVW20vA1cSeCMaUiw68GRlgZYfTy6XqIv7ZAg7GFw0nxqOKbl0LsNseCI
HbKhmI9DEg9AA45zCMYNaJDPrXp5PUIdGNX39Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 779472)
`protect data_block
ZnNvRcgmhEZ8QHU82S5FT5Gy72ADDEEUmMxCGcQxPxU1LztrbpiOuGteXuQRVXfuIRBH/irGW+Yv
LQNHGwFMKrU1esvg7MGD8K5+csocmgw9lbnyz3/qEhCilMWSeke0V7xFYI0XoWBw1w75hEDl+b+Y
YUO8x+hXPKHvAkQdH3jPytc9xAotF6XM1gSWupWdrt3iakzYtjPuO29LMtZvTlZQDzWTA7vK9/C6
dCt9SmQeS4+0cr7LRG0Sp9waQQ8JzdaR0FnVtSz9D1HZJ5QW5S4KC6RGfjqsPnrqUmeyyKRACVTv
MeDSwXKVfX9X37nxB7dAklWPmn5sm055JbrddpYgiWSWjFx5vBOJSpTfK/XJysQNL0wavjaWJ/8j
kMcecm3Pp4UfrDaZtRyRtF4yI0E8eXtVMWyO2ExGfTjxC2NS1Bgmmn98NcyjASdKUrszh21F2GjK
HLn8nSKt5C06zcEasb3D3MlBZXLoj1fwGfId7dbec3inGUilZ1xg4KPOx3AMHnWTtN2/+nJP8sW9
2zNULVyU1JkKmV/C3sx5t1WAvkSrF5JsTyVrCV0d73eVDihZo/griDbww8Kuu27CSvr/bI0085xu
QVGRFx3Ekl/kkX+AXZqHwYbtszLUhDO3lQdqJvzFSPuZIaGXMjU8V4gRPZJkXaFFuCSUaKKOp61B
WWVuWots3fLO6DOQG6+yrC/zBdYbGfa/lJgyBSf/5YkU4/PJvPRYJx6lNWrY3QMLNYaJOi6/hQik
kEvq16OMFhq93yGZyd9rJkwY9vKlZdHBqHDD6sKjk0FJq6wt6hbQVGDsLH8l+WujQo3DUVCfcLbX
/mba/zHoazPr597EwpC7CkBgkt3wJrXCysLHSgxL1qmRj7TLqxdITEs28WJk+gYs8xlQ6ruHmFVa
p1BwGTd6bzhGH/JG0H+AT1NR1ye7D5pbj2A5h0adqwInV1PyTO7cOJX0bNMhS/QKnoR03yC9ZFJ7
OJrUs/DQmkI+WJG7/2W54oIIQC4AX6mfYnbEhH/04l171RyIMPG6/FSr0DfZO+usP2u82YWl57aJ
2+J8hEWrvaZCIYOCVE77p1ndTeHBCRoPKNXpDKsDYiU0Ek9aVjMTLsw0GW6swdX1lJwTpC6CxMtj
0qT9p7L2mS0kZQoxca+5fqW61b8CKEP3Z1RIAbqAvDegJtT4gkX94EjJdvvLfiOeyL+Dm/8WPDYQ
qVnOc9vj7Wt4Hlu7O7SwWd2i1IIhQi1TW4a0wEwE8htNTtGkYeL6s5KPGvnp2c+4Gr+NJOidf6+y
Kz9dNeYDVK9eyPKrYVjzrufDasRBVIf3iBU8af9OCCbWkBLaHQ3OcbMhiqu2zlLv5g6EKwhG//+m
J8JmWaf8f7UBbTKDM4aBs9VfFcyDS8zBYAn1rNJm8ad2OqrPvoEUCpgv5kPACM/00HpVdGZmYaN8
yCaxnv4T2N21Jlzd6gbTSrsaiQZ8y99hXw57hstHOoSeYhn7nt3V8bmgM/gcBwNdZlTWUPLnxDlA
HH4repfUMmmvdIOK3KjBgd06G/HyR5w8710/FE/zb2SZeCdjXfJw3Fxi38WKjCEz14gsiRKnmRB3
Xk2qJ2o6KpGtrbrGhzSJs3Z7ab0n5JZLMgI/hJl+ZFPwOikzu/0PUtPISt5ESBDneyKJgPiYQHtJ
Qr5iBZt5XvSfLDT28TH7QnGgsiq1yG95o6Bi+u2MV5rhMOkhJDOgHte1C5NpK3meNhaHaPLG7sGi
nlKQwWEE99p6WThfVTMlTMqX5EIP8A8qcgqK9VIlyc63D2B4eLrbhZyKu4nKKWRSST+tUoWapTmn
Kep8hlj1A1gCE5LS/StGYFnL8dJfCEVgrE3i8i2pp9mTAK5v6GsYIVLIW/qWcRoUfDpeFtCy+lJT
JiCv5SEkWiMG39hA19ZKDqyN6S7W+k/CyB4s9hXly+lrL8u8kndmdtj+R3flTDwNsvfIAKW5Utcy
RDY/Rv3pOwKW+CV56ShZGPWSjhj1b+DKqkEL+zjLiovAs1FuO/92SO6kX0FA291Aev0X5LHkInxx
OfeMKWLGAQ8fNIe3DRVUq3MmYzBUuOAhZTLjLfTe6erai4d8LNZxANXHWUEHZKndOsFb1p18lQ6N
v+PmOy1Pmz7wz5VvGTk4VJI+Mz8iGZ+V4ahFLPywu550jntBXEQmutAESgtzJtHwEmN9aAYdV5Ii
/jBX+pYqFsuRFRihS+frRXPy0HM9fVcy/HBT1VB+P6haGq/3G/wRRQ9BSNeZLw/TAoAqL4p32dIe
B1CfmvzfdKs6XShA8AWj8pbWyJYcY9F3F6tGYI5WYpq5IBoEgqCQ1QSJFr828ME+iCrCw36Po6cg
qWHGk01ZjccBwhLOaU+9kzPIi5Q8J2SvAatEAir1syyJabPe3iplHXvwo9sNJw80zbsQ7QeWuQIj
6NKJdWBAH91VOxg14AXJ3BLl7a9ieMGBooOjRTvPJnd+cpeIVRFRyhDPdbka7mPX50xLwHL/6r0t
FOZN1AXmuoyx102ugCcsGis9oAVXx0Wz8ep8dSgRRpyAxQn3xWMWgXg8wI8Z+mdfqTV8wgEQmciV
vo0hK1xu03fG/1KJiMHw9oUPA5WL/TFSZZnW5WrOb8jq7iyKdfaqdvaQTYBCmq+ALWafohUyCAXZ
/1zsoi4b2Sy+9P477qigmX9B6BB1VQGfiHITj9bGIcNaIUsSjSXw9D0gjEiOO4OXQoe3BwWeFZar
keC4z+Kk9pZqVilNCyz/XSzVgLCu3f1K9WjEWyO/xsQTxEWIvSS7106XloLN+96zijxjt2bTf1OI
RZEfrFcsHQG7VfkzHFCS44TgPMZXWy7gOwg7IiV/j+OSO4i84okC4ayko5W7onZsf5FU/C93WBQq
6j33dGMPAIzP2BAX8mqlfIfVLmISNaCuIzS1wu23Yf3VD9kYuHVzXmPgqzj2laShuKagdMONFD5L
+zLpE5L4tekUGG9qq0Fr2pvsDUI6zyeWSndEb0CAejB+PEAa3YPH2UuUoYGeDNZ8yJjNhP9F/vlB
gxFQ2b1j4KbxK5oHkIzep8K64pwqoIsTStcHFAWDIXcnBjJSIQiUhmzudq/+XCm7bQkqBq+j3Nu8
4pmZIC92l3FyOUMRikrrh6eI5Vfb9o179PCQFnxKsvt8KGBzXTWZBzshPjitjfElsssgrcuuNI/V
Z9pdLLJ6O/75Gx4q18oev2HP3LAufaA7YGWGr9fkgdZwFnp+HumYyFRUizsd99Onea2WFqGSgxi8
GTXSFgepkvEIR6kmbW736dlXz6ueAGnoNlEQ24Dy9CTrNdAvR2P1W46buiCwm3eWijn8yEOn/CQ8
gnUGKP45ARlTEvdvZ2Kx68Kf2KPy/4V5IokPbYjlg0xf5NxNV0NxrVfT4drBxpUfGHXKt+I7F2c5
TJiYMnQSD8U6hYmqIxZjyS/crpAc6y29JgDgDj5I6VANw0FdBvRaOrqoQnqMG7CNSayA7TFulctq
uIiH8lpzjYE7ISWDZOS27zjaXghGDXsvEatDhfPcBNaFXg9p2gl7G+JF+Y99hY9UP0/YabAZKP+g
Bm1S8U/zqZUgnEwKIgAM5cINy9C5wqG/K5Zvuxur3+aGJ2bEYv2myGsG3673naunJMfGGmlNUtgo
hNzqUJ5b1OMi1GUKvWdLa6FLK4W6WcuiwL+FTxM8qLhmI3jKPQz3StR7D9vafyjinxEiglqwYOsC
QDQBe7W9hl7BbAoB3wuF0oonyjSY2vxRQr/FEbx4XSO2Nhbr9zXeovRC/IcZl5qk76oWhVcmAtvt
4T6WZ4bgn2tbGacPL/ih2cQ1rv7jWZdS3PX/+PvnitQCjcShvXgULV/+s2cGSltRlYTNN8lQ4Y/T
FyXpECUOubm4P03L3Z8o4c3ieloJ4GYJeGmlDoXog4S1oEVn7G60FsTNcCKK7wmnZfT4DIBWb39M
SnLEWbbxh7dFTKSaxaPCAQdAFLPqXrhdNwXKTX0h01U5yqus9TgKXkYsTgX327wh/6m3B75bYxHs
CE937AeUlxB7maR0yNLZBCg/RJbdrp7YC62r0K7kGQ+w+T4YZd0BLGLoe6T5Ll0EOM12MbFPkf03
CXBWZgad9Sn9E3bHYj++2lQ6UHEJ5i0YkbGgKNA12PTH35ggL2BJFUKZVFfh9YzoJmkD95aUPRm7
KDodGrc+BVtEj6uDNH18kpjcjfatPyNxXdOSwk6R2XLvtVNI1hAoLwXYybBpt1iwZuONOStm1sB6
iimv5guEEswPHpmf/8mUv9n+fcHifCy1sUK7lc125dZqbocaMBTd/zsI/BpfXParDLKbPhlGGRhx
D3nyvYM5UAhMKN1cxRfQNS+FNgVa8yywarF8VBoVKsUD1boke8lWH1/mGrHofZpZfYpqapK8jZxo
Y2v3mnIjdHdXdrNPVcoBv1lGL0h1bXdagejf7RCWcikRYJvLpa1aUPsTOEQoWX9wwLNFd1BAPeEJ
0M581hYeLslhz1EAzxDH+dR2rcr6QS3eya0Rb5qN9L7EosJv/iBBC750mxORrlwAzbv4kakkt87o
dyuQX3bo69Y11sGbo69233kh3wu+1JJYWHZnjN4KrSGPW8VHN/D5mjsrEbhcehIeTznxaN+1O0wQ
rt353icHYYABx2Whg1AnsEXtdx8w3weDeOmji7fFQl8HGr+8dVFxNg/K0189m6dXLtg+D9qniKni
6foyZWdyAi5kh8MoodMNuOu7+30boS49+vZMj+NpPFe5DtReNbas2Lsq6jwJ1tBbigKdYJQtq9sR
Q5LHDZDKiVDAIi1y18QZONb4M12ksPVMODk8rd2PKgNPT7R2+Dp2/EXv69QGUr+VAM1xe7uBYWZi
24cHxC50UM51jUwbMQpB4wo74wYQSEAwnwx6NJ9ChdrCSRiLfqbieSaGdFbn6JzNv0B3GVCyvdrZ
OCXTXq8cn1EzFi4Qw8hiG22+pfo19Qbk3GBb/ovkNslo5Hbd3hrnHfVTzWMP5v3n21YChfs47wIb
IegNp/f7BfYvb+TwJMITkexNysdXTWnDbifv+49qJ8cCAsJAfAbXr18D//iHonmuckFYIuYQgOnj
csrixHtzAJs8GygiBTbXSP9qQelO5KE7gOQmi0RRnPcYIbx8BDk53RGKciHEFlg/+0Iy1lYHAGju
zGnMOb23wRDYy0nrki1b8vNOdHYhvJ6PCGm65DUlf0MpxCdwIXQomWkfkaOwVKjtKC2BFRHotPn3
T/NNwWURCHrctPxAdf7oECobVUP08QyQtUJxZeo5M2HHsUeq0bSYgQoM1RjfWbv9S8ejwqJG4ATG
dZz9+Lpu8Ke7My/Ws4VqewMU1bsLbcX3T+vNN1vCjeqExLA2W+fFSGG0M9cNmfT4ciQYrPbXipmL
4bMffW0WzyojfIl4tGzXTsAsVILwzFYEPdNWCDsGOn1Aq1Ar8ACWZdBUT02wEFsRNHvM0aRQj5nc
l6EukjzCGfLrnzy7eNtzx4CaqwX1feoRAgnsDR5TGk9P7w13axWUr1gsue0ooFYZ9HUpo/mm2NNF
3X9RKY+QlfR1XK1Bz+I0eDOuytFp6hpKiG2tfgefV9kPWE5yNEkwj6Ot2+c19aNCTVH3EVM5/Dd6
ub3LLr69L48416ajZzN8AI+z/iD5avy4jArX+BLDOJGkBu4YQqK2VS+8U3bCPauqq+Q+EbqGHiuA
+xe6G35kN8FeH2zp5ha9LnRfXjSVG9TTBcwcLcqZajjlCaw6FysIH8/GHxSlxJJtve3mWeQ041WM
eEMUbNn4n09yFAQvP5f0JwcLJ7XuX3iQszBt257daS2qI+1/rc8CaHUvtJ0mtoy/FiXiiEScvV8x
V/W5N+AGE/bkYsn8NW1Hltqopi+FSD86ioSkKo0fpzxHNS5jqc8H5hMdtCOFFh0prfV37+ddbFOW
rLCG3cdEtoFs31veTe2VhwPjTLXfVOuhGIJuNUQi/4ZmiRA2Y7XcEyyde/ktOjDb7HVOwNOPDVdQ
N6FWGiezjHg4pyxLiootaccmAavIjc66nAnXz1r92cupZUz+pZeq0L5nBX7Khp0FJ7oU+5cRinOB
gxqOZsmCan1NCMf3USi2sCmGY7e8HMTvN/i8kiyeWGrHjUdfl+1Fl+jAKTRIie/xiGA986hAmWhT
I5NcSYiU4aAVBdhpl3qKb3ikQ6rrGOiB6omWOK5Z6iaNCux4TDZSJe1rzQ4DyqS+X0womwAaFVWv
YK4zLPqOxFgNHlbioRCvGpFbnLw21hbmoDzS+L0iiKdusBw2oMOHW2R8Bgsos+rWHgBNNngBRJl4
vOK69J/8k9BUdpKdraMTS/MW0brR8q23c8wQdGtjZ301IlasHOdZAv665TX2bXaNu/EIw2W5W9Lh
siMHaTefURosEfVITeUQ18BQYqqfpKpNavlj03wsWLwBkEglKQYkBof8ggU+Q6ow/fNB8gF2fYpv
bsDu6V0mZna+KacsO6ta4T9uE4wDuPJxNRHCzHGQttiiDpXDJ60G/qeibygYFsQXYn4j40cbUpHT
our7W+MXJu0ydydac228ML1g4zVJnivlXjBBPa+Yr9LmFtsuWQHmtdi43hdilUSEWdo/ltS2CfwF
wD+2jPgKPNC7LwGwp1lELNcfq2MEyOHHvV2GQhcRW9WfC2zgWWrUEd+hnsq9v1MqkW4JJAVK4Alj
Dmu5m4ss25HlP21I6S/FdO66BvsOazKrHmBQ/h6pkx0UCJ+p1W+OvSR/BIcewYY2+ghnu63PfhlB
QlfAhyF2e6COSX8o/9mNI4S7kiQ0FhPmDxBamf4iffn15v+WnFNR2DYcsOAJvrkeX1jxYwHjOWrT
Ehd8aXTyQlHIqGEsrb2r/UA0fmHmRDeqltn6uHJ4NqIhfY42jHQbxZv0Dx8wibABl3SzcoJyuhUu
iVxxKG4WSN4FLWCfCeyQD4qN5Pq996Vnjn0Jysa92h7H22pim3ckP7ofVIoMcE9H2ytDTfQmfGFE
BT1HYehRq9gyRn609wJo2OhgdBrWoJQ4ZwxjH1u4ECIO+QLHhIk8JSYAQz8Dh1AWHkvPyTcDOt+R
blDnpxlyLEt8zG/1Yvzt917S6ShxaM48Y2eL1KcHHON+PBygm4Eft5IJHD7UIOYMg9HjZajr2QxA
SSwe0Onxa6+euZT3RL7T8b8/JQp0ZaQwPWm7ZJWPPQ/tBCbv0iIb6S2M0yqEWYvU/Ebyh9tfYx7F
KVsHRkdW0ClVRNgV+g9OORES6m2z+lSv6HNTnzgyLweqrhjx0Ya6wUEM7/do1UJb3B2Lev8K9VGw
SVjUtuILeJNgAKtBRIER1ojZhcLl8pcohSl63+T5PEp2hQypisCNVt5oF8yHEU7jzCbs2Skxn5Jk
n+cOj6/q7saFcyA2CmN5Iw6YBwNEqaqUZLR90/sW0BskTRfwNpyjjb/z17bPCaHTDpSPbVqDnV9I
3EMg9XiJPYSfPrs9fRaF8OBe4T0/4xn39ymQvnEKck+GF4HabZmtc1+2PVV6zG0Aur1cT59rMMZ6
Pqoh1v/5k8EPrCSGMGqtThw4wVlLGzvB440/KI9CFHf7i1hgTz3CZM65GLkAfXT6FQyK3xU3JQsW
NgkNwtJhyb3o/nyXt6zfzTl/9ybNYMzql0wYJRO4LBI1Fya0ijBexLb8MyZFJlF8yeVhHpD6dHMh
QHB1yNYNf2AeWFBjaB7tHr+XfxuoKv3r7LLOFYTnNS33yu3dHjPmROiuDdGZXoVcGIrYhpMl7drP
EV/bJtzVW9iUM1t3C6tU/e1iOFKE7PIRXuHmC+jhoOKHx1UFqIU2hVNB5qaW9YYFRQ1e0fZQH1cf
c8e7j3D2xskHyiHsJicKxX786TyZUCGXc8TS7cFVnqfiRDtWGhG3wxAOyg55UQ+BrlVW+O5vtXcm
JgOv5ZG3sGAh0+ZQPhrfnlydtTcRclaGa3xF4JJBLWLvjdN2bNjkpNeKIABeugXzmywImpSXO+Fg
5SjjgfB3EMPTTyN359jvzWcNKKaSLLFWwyfUdBLUlsMO6Rm0jODi3UGeit31DoILIQePlIceWMMR
QyWrjWrJiX4jENpJFCyyvBWucxEwldZeCpaZXo+GTEQK+/DTYz/lCN0ma/qBsgm2pZz5Q3Go1Dqh
nbI+5c0Lh0BM1Om8I1Zg86gCxs4MMKr+vV+1SIplwnddofxgOZXsE8c6Hq+V3KQtIVOx+ECBn5Ek
ZesUH6wyoyZ97lVekLmQehAIiIkZkZLf/ZorzCP3bdhfJ+fUxpCXc4ztN8P6XWv6rLgxVtvBEkNz
ariOpKHXweKwDcd9rGpScfu0m7Tx+nklxACcisw9fZQ13glhP5e3XoRM3WvUye+j6TCoSNM6H2vJ
NqhvCuWfdxOjyjruAxBGbIgZTQv86IXlzorRGhHQ7kW6MzMOlfltkE8htx9NWCA+IJ21VNsSXxHn
n6L67PfY9LjFZbiC4yu2Yng0ZUXVXXOW39uV4As6OGKzrMbK22fHH1kElzJ2oFqp50lS4TuMg8nK
vgm1M2ihrFOPiSRNiG5JnMUwlw8IUuE+7BoYwiuzyM42Vduzdij7ZH1gviOI30hgRXozv8ZS97kK
lnCsOQRX7j3CF22Of++OvqK8MpF0uE2KZz3aj4CypirQIFOFiVr8/tC+Ed5fmmOqUC6JDI8eVd1O
y4D+6GNCjucX5Z1NQ59JYIvzSKncX6dxWsw9aMZxlu0YI0B/PNnge58AkD1PPumY4jnIGl9pAiyw
koEr2wf6DCZG2sQ5KPB+OgGvjePbMR4RUa+HtTarEHyk/SXFUFiP7kADQjh8/1AWeJA9UcpafTQP
6WPSxmN2WXy906P+lq0NE3Khf0mlk2BCC+nWPpkP/prWzf+02aLOxP7FCescaetLB1aGsIxGa2L4
oOHpiuOpJ6cXuaUovV85m5no8Gu/NCiAHgBlJPuXsfPq0oWbeGz4/aXuqfSzgMkGYgPq7SgD8Zdn
ZvSJUF2EnbVRNicERAKeVJA6CJAKQfA1GzIao1e7PEOzSrFU+WDpyjR2HVBxk0aBjtKG3nJWBN2E
hemVRPNC8t2K3t9UraDT45gcS7GguLdzS1RP3S1cSUePgv3uQoELoaXOMQEiyQAY5uPw4mqvaJoW
z36n6OBUjL0vHdX/cVYO4ZqHwMdDB9AGvaCh2+rnr9vnaXn+cENNj5XdFqoLNxFV+WJ5n+G61WBx
HEWsMw3wioons/BCbkToZMIY3jvWfxb4h+nB1LABr477UAWORUk956bPh7HQLKJ0EOLpBAZEpbWK
W6BJEHIUAzquob7frWHjZPuUFATx3RVNXPCghc3qmMxbyxDyUcH8MH0lyyr+1e2TPRaGrQ0vFOHR
vKiCjfZNvy7KPurdaRj8lZ6FHSlBdbVW5EgYXB3isys02+VFWf8HIDNeth/iSgKSdEMt72sfwUYe
UoMIgREVbj5XJwGdLIGnPwLBwf6/EeUYwk2GXGkaUQ3rC53Ydc120T2/5djTDPNcwTjjmTpkpz+B
EVdVaK62hXOk7VnkVjgTUlqodFCQ+zdnoWsBOkbj2yRrs5Nn/KxYqVaHWIzKuBImDbXdArr6D4e3
qlPB37PaBiOUpPYxj95aLU6lqa1KPuX+8LFnbzXQQcBvuJ7iJ1bd/4Rp/32BQPqzZabrXfxBe9ui
6NfQIrHe3aeS2ociqM80QlPRY8BB2zw7ZNV5Jv71kSKE4Enc57mlqfuNw02tSfiQPkcFv9QtpzHT
HCCJUKi7K4D0FYlyG00SM6axFE+hL2ycNVKBTgG4s0JlXCh1r86CmecNs6gr+3oscNwbXN6pc/f0
ofJ2C9awhFQDS6GLckxK161b0lZOFhoXdXXJeploAMnGFuxrERL/3/2biVBfE6Ef88O+5PPAOE9A
vjDKPtp61IfIlk5XEIT8GRT39BrTz2Dx+9kv9E9DKxiRTKgAjJcOvIUD1FfhKRDDkLEI4Ma0STb3
mGRaQaHHuSjEKWnnCds1zHbOqh0wK29RidqT4I04n6m2ZHJEsbH8E6eciwwPHfZBwl4jLZJ9Uhdr
3XYFBcd7YSv7Zjm8PeYOoZ/E25VlD3xOM6qBiRYGcBNMu8zZNhUcmQLARWJJzg9St1V5aaGF+g6s
mKpWaj5cobXPO1O8YxSyPwOVz93q45CXO2G18jE0Fo4LzVUReqIp/pma2PKFybv0+FfEZw1Z62UZ
uU7+XlTUmuHdy/haMgAP7TdioZtivnqBapLnmbiVEksTCMzlXWGXMlLEc2ZuBHYW5PyU7Bme4jgy
O35WKRxawa/hQgd2wbDN4yvBaongt2vlsJZLwSvXComWc14cskxBIrZyyQi0vmLSHkXGfJ+I7UpA
9ru8eO3W/bFnhR9LJ+WMu1IJvUHSHSzoOBOqRYuIYg6IEmX4s/LXrjjmx9brboulmr6n9uW4fg6F
LkQgLa8MWrN/6Y6N+dm2ucGeXN/svYQBCiu6RCVKQ3OsGTq2UL/h392UXF64JX8d6U9icParyPIz
LauL/qkxTu2NzZQ3Aj8JntJuVPU3f8wdlo/A/QnddtfN2QJYXsx0bkbuitATBBY6vieb1F9NKgyE
Z1+w5YikY9CThzFYI0HSt4eIZTris30XUjkL4UBhYNB+/+bzE3X6K5zY6IYlSsKqoJmAd0o4z1iG
Z2qSJTKLREly420czyY32HVm62jKhaps8gRjGA82PdDeA4o/MPjrmGXM455aktgDgS1on+9k4qyf
bB3oYIWOgu0jW77lWPwCswa7KYkJnAZtvjcYUFsbqziStKc5yWBde1Yf/RwX+/6wrGNjUK4eHdyh
UoK8AiWx9xK9b8CINyUlQ987If7q+B0S/D1TCFvbJqSExeo8uLU1gehJ8oVRgWfTBRmUEmAL7/zQ
vmNl/pRDCM5rxsq1kmqDSwyW3SnmEyDv2gNsDfkRmlta8ykWKmS+RQ9UNe2ki7WItAdKxAXLqVIW
JiA9T9fK/nLgIEqVd2BrnklogqP2xKp04cnSh8a3Pjr4j7Z5DRFGdTRJ/Ksny7JYplIobzfHZcad
9bIuf1e4IAeF3BYJ7WYHWkEXko1RogRh8cLHi/B+beJGSanq3wGOPUYebkY41n5kXflbUMsuSAu/
Ovqq0ZqyRNEHoWdcK8bFeaNWB+giFvBJowMZtm6e9ZkreSFw0zFO4trPJV30NCfyjxtzMGxE3AK5
5pDjCix48rEWMrOYphXUNFju3rkP40thPeL1l+dPQJtpuZjPXRgRqInMYgz1qMwbVLcBTUVi31oc
96NXBmYWXfsyCaSahEtbaHhuaP1V8qcLJRlhsYeFSR6T21RRZr83kKjknaywEqaOwQKOFPc8aTPH
Yb7CHZOPB9E83SMbS4gA91Pxteh7XrMtP5xrIdfYF7LRx3o7yuMymIHqAUO2Wk2gXIOHcoYMQvu5
KYLC0HrCz8DZNh65e6WDlrUR1V7Q/vRE2KfgsDlRLuTWuuOB89XgZpVcuSEJfelesbHrE/f9TNIj
U1eqnJkWTd2VoLeejklCHtEQamh8hed1MeFfLj4IKpRQN+ZTgGLcgHVeLBTiwX2C4bHqTcCzWpRM
pkFwbXpIrDBpts7Cuwr+YxYZv2+Va8oXrnqxQ4palVfRdrwIVHJeBL1keXOaUYgIAPH9nAKWkehC
4tesxUNNeyY1ehkSmM/NzT42HFlAKsD6ZajMBPNwCChXIFVTpMNNYcK3V0aahMJLEjztovVB0akH
YQNzeGAwjMsflgtz4VBnQICB8Ak1QSEBzPu3161l14WG72isO9o5VsAt71enGmxACqkqrmVMQCK/
/Y+kK5eAP9KaZiGCwNutcBet3HjR6Imu3W3pZK9QlUD8Uxs5s2Tc/QG04QM8lq3htrrNRDHEoxJn
kNN8jIiqOFdDjDMEXTw9Gl+82dEbABtS4oUxsYwctb72UckV8+09OLRTKvSOOcoXyIUurenJ42IS
1qZF4yQQ8I2u/DCkUQmzcV4OzJDWhb0kIlhKibM9mqsLfz53lN3WI4qr1PYOlKuVGI7vKozZPz3b
7wwkkAFMJB6epylVYbu4BqECwi6KaGjjxYhF8/i7yOx8MMAG10HwG1mFxHjy17T2z3edhSZ3nBXs
j5h3nD1Hv4hcqPNrQu/qNxYTB3eNRmCqAnkZYvGHJdk0grBbkFM/eXGV7jRle9lShyI5/z0IyUcn
izeaMgt2wkk8dfY9ijHPo5MnxQzvPGsnnmY+mGyluzmY0ZJzqoZflc+XE1UkeyWycfjMNi1UFk3u
OKZyzESCLwoFTXMIdexI0KxSgPEyMMZ5+rAI/VZlgchfXJ/RpxBJuo6SeK2wWmzbbBN2BM/kityG
Itb+Tilb+xSUeU3V7EwWz+I63gDBlwNR+YnEECeAW3CrJAHqGpdYvMFFxLryJlN4DtCKkFIzbV/G
mW8DQyXM/ndqfTo5CwzTwGa3G1gHvsCq/d1jTfHafq9oBSCK8Ctj1JGOxdHBG0/7lM1KtRGZWU+M
a3HPskLWisp7l4QHc/UiTZnsHUnkwbPo0g1Lo/7R9SkqAnnj5AR1aSeG4IFXZKPksqY8uEyhBCRW
OPNnpAD0VFBr7e3rZwRWB4AUnM/PImOqIM+C+byBfuYMvsdpjq65frS8oh5vI8+bkpnHRWmuLOWX
CpzWYxnTFsrF9sT9GOW2dsV3vkEXjQ+AWldng31MTkoUWMHbkb0mQqSmKLuhmoXklSY9Djk92JlT
1AUlrkX+k1CPLVVa717WUjHJxl7VNkNvM/LiETO6nWUO3ncL5o7KpduvUd3RbMV1n3RNH0lndWXD
t8+BUiIJxsC3z6AFXiqY7PqNlHwh7LsUBbIjhlZNlBr9m/8DbBDVT0WXWm0mdmCn471jXSWc2CLm
3XXrK9KG1DNxS4vRnEZqavnR3/VIe6+UXIATgtrbU7sSOIB3vuGcE4UerOaBFdZ2FMzw6EI+XuYI
XomkmLo9Yx86/3rBd79Vb6NlR9r1Is/o1jltltJsyCAAnPnirJcc9DC99Up7koHdYQfpz+O8y/TR
saAqaFViSQdpUc6csvXJJAoaoWYof+QSrERW0eiCML/QrSdPAzJC8PB3c1+AeLLcbVZgdjMibU77
o5QGz53nuLFdQjv3yTvyCH4lfFIUKI7SJfeAPDn4A/eWX+Xir60gIG3o/IsDa+mM3uhMh09Ja9Ld
7WlCh34TKuN7NY1BTfLzPFRlQMtaGAcWf3fGUluIL7iKBx+P8rfDqib2ay4toRxAxLOs2I+hKTBy
M4zdyXFYWUgSROb2MqiCwk/1xFyPz5iVO0mIOKRvphONAp6pHdQ3AXahHULcO3UXlCgnoZThQvVv
O1fFEsn+lwwM/3G9QZA8G13wWG46SONanJO6EOHZrVJSaQeqPgcKPSOgXJRLBSQN4EO3aN4+ThZT
JGJczlk/K46tnx6TLCEPgLFhhH2axSNAzny25DcP6pFjK88eJK7xBBvIGKlYQkpROcGhIwLuKHRr
fpxfGBtIXy7pOTi4ZE68M64GWJ+hemE+ZKxl8VOZspl1iS9lbjUpwoCehT4EdQA8p/C/U9OQLLJN
rA6t9Dafn/lbaajsiiyvletn4QIG3E/9dFEKNP6TGGrnnRI7INcEMJbOZC+f6Cn0VcRSSrbonx2R
NYvZPILxAe6TBYWLlDAU/TWda+Zjg6l5h2FC7+r8ArsXN2Y5gtTmFy0a39nSt5fFnNSWlDqUnPaD
KTRwdGnc3MZhTGIwK9Zik+wsbAgJJPZ4KEztnzq+3MYxSNrqh9vwAec9E6JWEZLd7+0D355F2qp0
Zp6dKAhENQ9unS2A8ckS8u5XeIKGXF1gYb0A6A5kpYVmm8f1NH1qdC5ZKA+YeLYb3/AKwVrQUphl
l8GvOo62pAGlStQcIeVMQp44xnwIB/Ue2HvhsprGn2J5J8laR3GyS4X41vcuHK4VwIZKj0jCh3YX
YSbJ8XvcS4cbvjcbXS12p6jQNqk6HAEeBiiyyAJKbptJdmnCY7+E7Y/5RPdWtT0IE+mudvMSYdzP
ywTzR16vXxXDk4RYESkbmRe5BjSvnPNe/psHrjb0lFI+ND3oinj0CbASAiuo1bRM5obrSedzaSnH
iqc4TSIX469sgvB+rh6kahrVJ8jYtcFotH0r8x9gATndaalbucJAE/SkYWp+Qxi6MoiN6CvNDSyB
R+3KIN8gk9C8TBDnkduDJs2vzFT2YLfSXz4YRtpopGX/bfze6FvGphpJmNT2g73WX4HAuRQCDDl9
IiLS3epVoNW46htGbUDT71+LUoiWhNDCUkaCbLmPiquVNjWaI8Y0i0LnNNVr/BnQPxUK9N/JVd/c
aS4qDlGDAUmZkve8HXsiAryuQ0bbBVXuAEyYFoRAT3/CUcmXJXo9/ur0MSL6f9+paedctraCoOB7
Ys6KoJdABpG1+rQliVvp8qFI1QLZcTSFJ1KWmQe6K/3IVvg/bGocX50wqqX3Zs6Pw/p4DxJusy7z
7nGu+w/LSGmzeQl+QggJQaBcN7M9fbblTiVU0+8xOHrTJAuHo4WTIfUkf/KpqI871Y267eW/UT08
Tys3gYZLC1enVq1z6iNJr5CJjddVZUnSXD/yMH+n63tGJ5Txv5HU8PhGE/3HmEfXlU/vGnqWEuTw
3kPoqevPKSSUkHAqUXyT+J/pq3sVxZCNjuWnSME6PKgKnvW8AsBQdPG5rxEadJVkyG7jcFcnxqCW
s8oSwEyyH5tJYZJ+u/UkMwvYrFwotJCzh5C1lNOL9F4Wf8ys24BjwGJG243j5EZ/b4fNXQZK834k
Pd2wifyDOMmRCCn/caSLAk56cqgRY0ZMBcJyxTMY6foFP0JskEDJonZ15dx32zy6IO4iNrAZbZ0v
8CPMZfjLrh4xd/esFkZdKCzcz+CGmb4psmkeOAbOwBiRBJ4H/PNpnmZikLCj7AKmodrzhhZv8j1r
9zhOy5GrAWPAzg9H+YnWTdlJ2x6tligBNE0ZD1TSXnoYURrG7+PiDP5z3GDhLGLYDhhFm1QRb0MQ
dDDguC8rHPirT0Ea5y2LbywqcfeslRaLeGLOO83+IVz/qKEDoMP4FeXWIlk68XxydRMM7JibR71O
gKFRfr61bTJJJudfPR2Yn9x98MsKLpHgz8YrFZdtHnQmxjcoYzWaSJsnD23nULz4yOvBH0AfmOyY
ttqRI5uPOqYohPL9/f+tKkin8K8tF1ChddTyUpMGmt7wcVfhpeAj7CT6pjrzWQ4bM3x9iZtt6e4y
T0SU2zJRaY4QH2a5QIrFaU5Ro36en1qLduCXBQukwgU91Q+wmVI817iWv+UzTugcqM2/0T41QcUz
2zAKV0nav/JVqdto/BkBJ/qYY1jiktOUidw2/HPraT9UOWwe5FCEUr0PtyvCgxR00ehOBt20cbhP
mA4+XhBSAg4F0UMcxguG5qFpwogQDHwHzrcClkFsBJVX30r4ptK6zXVBkm7ETQxd199maSW2Fark
JGPT2/FV6qJUglYIQV+T/7QPFB7H1ATOH2BWcU+lhN8IroxnxucWEDf/tyrsIpLC3xvFR8/jVXzl
ire5TwiFBwk3KntL2g2HAnbVd9NEkaf0JqkOQzizw+u8VPXsmpuoEWR4QJBMIyMjuNRRFfW9ANmq
g9jc8xLX51r/thi+F01CFdmCwqpxRkJOohUOz52r6tqJpMZbCtJa6r8vW5eznE6w+HbjhbVfoOXL
xeTrKcwsD9gZdOEghKLlb9MAH76W3KGNGWCcvNlhc/IERuxo+LM1cMO6C6UHuoj8BUsN7QaQWlRM
G5d190D8v9Uc0kt4j3G7wB3/V5Rh68p4FUs51g/ethUdRx2rfdkjhoZhpjtBWYZ5wtlOaQ7Sy57V
hTMgVM3+wT8Q9GXm45x/jVoGtf5MDCXBCYpT3LryPvwM0KA7YB77pWny15Hkk91FSIfy6Fu19j00
mMYbD3LcPrghPbgBh3v7Lz5w+NvVTLWquMf8DLpO8SmulGHKZlg9+MD+39tB5l5Tar/91Klqwk0o
IUfx8XTBuKqIDIEUt2hqHk3Yej3Qk8+gCQ+4+HwOq2CbNCbYFnpBJP6aWjpPTOiD/c6INQu5EWtM
uyDpKqT8IWM7x9cuWDtQguvEf6ertP/4oi1HoZwYblP44GtPr5nDNuUumUGK9jLMwx8qf5lAdXpO
M6FHnHyyAq5QlOG36emKc09dtDhe/2Midp04sGDE8hjJOihBWWxg5P9wbMN2EiTTyVY+gZt+4gph
YVV8kVhWJcbhCdTNg5oQbKWbc2gnr9wcHaUsScOeszwq4xNM6mxSnz0LuuXsPqhzITFZBrrVwVmg
LuyzDZn2EIGeK9CUnfql+JqL30LJK3mAJr8eh1LaRip3n27O5tfCFMrTF+bOGTXnVfOphqQAOsyE
r6z2jOnKvfBNdEnL2rDJyUIaxVwutdAKRuzj88NxYO218ZW+CshKZtfx3TI7B9DpRsRVXKcq87sb
JTjtJpQIdnvyv4dbAFCRI6u7fVz2x64C4RToqTB8D+n5j2NxfGadJBqcXtDLotKHp1U+1qxEbibX
lyPdFZ2n7LXJig5D40kuAYVZEqCzeI7AQfgsTP4WJXWg2ltFgRUHum0a3D9koHKy6N2W/V3WywhA
COLdcPKRqX1MlcxOrXfW3bLF4KtA9C2V+4iB9MXNo6rz/vCET/FxNlTixcNHw6MKnbeqiJdeUrgk
FTC1bMuWW43Ck5F9Hm8BpRftQYixfqIkEcdW+AYTDeRkHeImhA1CLfjvKkyl9nb6XwkxRpvSQjmi
g4kxSQ3eEx5p7Wax0R1C1MvMif5Bxjl816n10Xtl57CMRF3Q4RfqyTRj1jPbajzHhbeh6eNJYoo7
gf/N6Q5iYRsIL/jZ1FNhbQgxvNSLNmf+VOyMp+KIrm8NMjCCTsctPjayVTYESJpdPS5o/HwVI5nb
A7luBRxMn1zukZBuaW3pkf4J52nJO6V2w1KD8ghY6EP7jMBgaKGK3VBfi9JVpT3c3hu6NqhjD9F1
QoOw7DGK5Qim+AUy4nXHgozWsFOxjI12Ece1on8wSUuW/9irk2pVQV2oCNUFwChB4OkFciWB8t3l
DIgBPngp0pstpe4VxEStKPmtDSzLGL9Ql+fpWMc2XDlQtyGuIsSX6EMS9meIpeZ9f+Mkt3JPdUAN
ySiWWik9LWrL693eeqWhEb6IR0FIbnNZLIFzD0J+8p0pCoMUBdD0GN3LsJUVswEATN6APvZEHXUY
LvffZbrHNmJOGMaLr6ECCHfuH9vpd/ii5GhDlGujGA9/Mt+QeufK+wi51fqwwFGyKyuKwKSZwlWP
F3JOe5N9HxT/hynALqrXqYrUKUISm9ElAy7pbtEOqvwW3T0KLWLhzjxLt1fMrzPtiEHk5q+faFyq
KBb0CR5A/F1Dzf6dg/pUQNI4IZ4TuG1Lln6UIF4CZSJZu1ApIHX3HreOv50XCVn080JJXTBfVKho
2V/dqCsxmOe+KuZT9SGTBUvII7wZ6CvZfHZCEZWfekXCsFEPWVM/IUJnl4cQ9tkD0b+SBPRzjel+
MSY7eo0JiYfVYsSJ/+59q/zOtqubhTCY5ILnUv7okO/U6G088GTp+aQ3EBvMl35mq9LATQ66utH5
8F5jiDF8CewByi4Phrbh+4kkpqcHYerq8Qocm6voTTZOihuhbpilmamI/CSgIRkyOlr7gn1b2ivZ
7EI+t5r74v6xbdk1LF2PmEcsX0VTydeMfJ6PI181X8QzNwYz/0iBUeR5hQMTQverWQDgG+NU/e4I
7f1piEyJ3CZfyAqOrADwZ77rQgGgS/nVYdGaegAC2ZIRyWLO8AGV+6TV4aXG9c6QIYHXcLisQBim
FQISte5MNUbmP47W3EluUssngFCDqZGI7/Vlvl+fyoSBeZMvfypenjo5TzWgwJn4x0S2UlcqsncH
iP3zBdJ9fEqkZ7f5+Xspj+a4QKDQJjemnXQcZsDqZpoXNLD36qzEnc90onjxzg/GfDVS8HO/1vol
5pkdqag4OkOImh2q3PnVVLBSrEBGUr9z2q3+giWMCZAVhaDJ26tVQzW3tjiWbueqDTGQ1bA5v7AH
ipYSKUqn1w5cITQXD0SB61pRgNPHr67tngO7OpxqUyYMaCZtSf5s/1CzvrEGyj4GlgtulqCkH5XV
xsR2lNkVyucZ06W+5PDyoZ/EIWXgi+vik758xQhHc7+bNYo+dJ427E1xwVVefj+y6imzmlN6K9+p
isPEh00MNTL3voU40DGk9+YiQBiUrmW5ArFpqihBC5Y97jb/LO/KiiTunre/r6EEde2vr9jzqDZr
czIzWZO7G4HXIfG+6MTyoJQVUO0kDp/M2m73fvBkPeRCOrKSA+LhaJ2k+XsaTBNOT5pamBA1zi5z
TFA2iBcpD32JzYEPZuA5kBwA14rmxA5y8tCqH3ttu61EY2cYQi7ZA0GOjaS2g8U12xh2w5lwLsdF
XRHkAd+VBCXn/bvCakz5EHDplHr6VzDUCRzHKvfREpzjhSTpkWnG0NYWyy+KLaKVZMNcHBkPnmXT
DsUSL2dWGhy6K+m/Gv0Gy/1anzQ9Fb40FQt7uA7KJ6p0hipa1AeQcK2Q45NwoZgCIMDhRyJwgXH7
J1RXsZzaNUN4cizFZSdPVktKeA8e8J02sQQRK+i6tNlvuLFD6Dochg9cYOjnpvW8KMoPvFl72PNR
QleCAsvQs4CW4vytRS3TeCeEqKvjeZGO0diKx7eoaRJ82d8N8wlpc7JJDcSNyTBkdC3LN5BA5efV
W/Ew5OydODCMND6IY87XVzxTaNylrzTGtsSwDhb70V7diyfe78LEWFi73qsnpNmdRK5NO3dfrl6J
mi5NvOsH7CV3uUvzs936/EYHQOcnYcBfE+hkH/UcnWeDMHGoonNSC6p3QYMlyuGKQKrW3edkshgI
tW89gH3sogVe8yvT3L/XfTbFFcJRP1X9RbGpH4Q9sVXawBS29Sss0M3BHFPN/MfJ/yvf6bjlHto4
PHOnldNLJ7vwt8PzLeyIQKL8gv/aozG2upTa2F6bW/dQ/dRE4G9fl+XBBMoBrL6iwklNKxcgbnzM
QQ940kk4grSlLxRIurp4MkBXxUERT6lGr9RsDHOHBp4DpMLlSJTkR7ENY8H1ED92TrlIGsVhEIw6
QsOoNC/kNcQpwmZ6caefX40vXuhPTLiYDS2hFH5r8F7BI9dJNgQBPmFo6ug+w7WhkzVcVm8jmk/J
vDqieo1LWAWvqyacQ/Ancb4Z2sWmypkkOLqKZwcI7uT9q/36Z7SuThxvhpq05w1V+qwaNY2tuqv9
AakkRFgJNGvgwM8zd7+bZeC0RF0LGTJRww/LeUpLPBhFBgIZnJdWDkRZkeNsQEg0qAVbQX16cD2w
PJxXP0E8payFYBzvjwX5MeCBtCZ2QSMgDmb/vEY3eTncnXZN0/Ey632VdEJwNud1jRdKe8EUatu8
SqYKxg31tk7eWEP2rcjS39NU1Kr3kf+CErbdDfLNeeBjNqf3Ry6hS8UXczoBf97bFonl2d29E+8m
HR3VMZwwdDOQz7QAybKLqFzLeyrjM3jN9A7ZSZFzEaU3X8KJp0R8qso6UkRPmMxdIHbLcGTRefYb
WeaEXBX+PSxVqe1UgL4oLb6xfSEgGjUabW+QsSKrgFISkcK21Hcjh1WlYalHEebRU4WYR7YOCz4P
3EHO1kLtPt8BoQw2yc2iKTMO9W/ks1xaVurA/xtlekEIJPc9JHB48N1Y2zM3Oi2oHWwvpZLPe3NA
iWha7PuSKNFDUXB3ZTuPVOOaN+BATOl9hRrGGawTNWrD0oazRYxeHOxhwLsPu9oIGayo9gNaCTnx
hYqAKXJzVL0JywTD1LrbtE1CDD1Dg807oku7sGLC9GWbBxBhZpH6v2wsLoYcKmoY2cSazSP3aeYR
eD8IffaABIoU6ajxVL6Rx8+yIqXRYxwpDcJToUDMYCdd6ABr/HZzudrR9RSOuR3eA/mx2CbHN0rB
oIG6qF8Nze5QJMx7gl3WyTPLZYF2HFZecD9f3321alba0e+4LEfkI08UQN6xAi7Ett/aSO4ZFLpO
PIcKWTpIV7zoIJV0w4ePeHNtDtCHTOptQnP/ijwGoOp3zp0oa4eL54IJ5BIG/zaqubjTBlg9ATL4
8duSgcL+kh3uP7+RdSUrEHaj/VOhJ6xxxKHp+STEXKpHhV+9qaci2Jec4rp3Yv0RY/gV868cUHWd
pgUFWJY8N0PJRXla1lmtmxyiT5JGNjH3FGeEFQJ0NiyDK6ZPfu67VyreXcHpMQazSSRt39yj9fFZ
2jPahuhfOkSNNFY4RXLLjqMsAK37bd+BSB0FOO1XoUtulnRCE+0AcM0Hz6YKthNdYLaWlFCpGpjb
ua3WZ0wmGq4vhsTzuV+Alz5kTfhp+9H7+hTCUkXyAWLNfGdquax2K0oThDPe9bU1j9Q99lI58fic
TI3RD0cVfVRvHupmIiDZB3CzKYx8l0NwrIGvnd54MsdMIkj69MxeWhGzGhl+T9eCn8Sbm1BMYFcd
1MakPfK7BNCBRXknkP6o5hIP6hURLJ9rAR6kB3z4tNJC4pP2VuZ5UHEFWIkU3XeJIv7UfrGkf6ou
J0w8FnTzG2o2knZMZCfQeKeWhUk6PlSzLrDCRyvfmoNBddPwaanYZHMMLZwE9lH4MrzjqTM0e+9W
UjkMNbLRjwAiGbYLO0TH/xwP7ygQz9osxzetk3qJSOd3ZQ67/HCZZH7KycFOGoB4ULdbDzjcYOqz
aeiF4PVpgIjjy/WB+B1KDMSKJhQ31doQjf44WFT+PwfVjIPWyPrQMzpuoFciJljeCNBhJz9l+/qx
IVektqqt4a66HXZow5VIPvkZR376xzmzqFKUyyK4K+K7aUJI1bUYsnLiPFsYet5fxSxhjqGu+I4t
7Nl2pK1DkJRiHnJmRUfIarHD2YncU12WWZg2w7k/h9jD43NU9oj+59ThxPFJ3npNgs/Y1f97w+al
2vTCqiTXFulUYHkVsfCR0tA1xFzSqNk5wAwoxlTG4TYtiPwVv1WpCQbxrv48wC/xZchzHue8EAjl
CWd5N4bVrtcuxAZSnkuNVY3h7uvr9bD8O7XxCus9+/rHe7kp9sUcsCDNlqmDOu9JJaXaTa/j381O
ZXKQO4noNIq0XrNyYoMlreVzyP6iGAZIifC0Cxfy+m7tTE9V30uAZ7m6yvcNrc10XsziZswG9/KU
dlwi/tGkAnn1kl56/H7mgyuDqszMpIMh2Fx1S82FGh3mMu6MOa0S5YAUbxj4Htzx9LhWPsPoTwl6
VnSkvbvRbbojnlsJIjya42hUdHDDHsT9A/GfocbCjLnvMh5tZe12i0Gslb+tmk00TL5BgbUOyLnk
b8Ze160SJrGnq29DncDAfF13hQhfZZMRsfRJBstNap+MfKa+qDFl9aRu8IzavxjW++F6gDwZyfPZ
Ccet/KuO0OOASTVz9YDPlIykWoGOH23ok1aijnGbaiyjpZB93rvG14ONgBxnFNJwCxLLrd8CW/GV
N3RotAsjXrbgHynoci87HKRlB3BztnDUbQDlUlt40xhrGMXQBjBIawWXKkA5pYfhKi1oJmj7YoKH
evXxA+3EAehR/AC0HxpG7RV9RHGo4vjbQmqaqGpVPBwt2BRfrZMR3p9/BjFoDEtkAbDnLn0fPS6t
/vgvnx/uLnIcxSveBBFKU3LdsEAp5MwzUJatjOyc7kb039WgJXV2ozkarbEjE8Mq/BS1tFP5Vpww
ldM1R5xhYHL7F1JDvO+7XtN+rVo+0A750O8og6YIzuxHO1Ga5LAdMuqs67EWVSmm8ZtsLUoMDmRj
DnYT2XAqCIq60esYpxMh7NO7z864RX4b3ATwxUqCfHetaH0HTI3VExkLGPRWnxxRK+OD/NxMTGNr
iUXRqNp5kFOqHFepWe82OPlZyDDo8kx1nT6EiTKBD9vOZhihiB6Ar8b9HURLQpW3KGnv6yE7D5/s
aoR5nT9qpydnOw7hDtWd6I5i0gXU39l44z3WBVXEcZu2OUOMNwLM3Iev8HQMjXjBnyrcOxqNhULH
nINPVMVqR1zmJNyLKrtYXkwM/WyPtlme706Lmo3Sq/V/quZ65co/BYNo0O4hCBRI7gl5nmgCBKbR
EiLNzICP2UKh6hyb6b0u70jHKP9cr/7hBjgITRYXWZ1fHiEuSdbosZ6PfAXTg/Vf7IMOo3VqCWcT
MuUybZg30hrCVPq5iTq9wXk7XCJQNaI1LD4SqqTGGAJdykmsNCbrJKRwccgsVf2GztAJqa0im5G2
TeBh5+ip8lG4q11fIbK2OnQCvwQaLm0Qc4jR9dmq+38zVrS6wxVFwXNXq7kh+8lRfPSQ/seW6aL+
tzY4k9PEsvg0YrrdHR3VKhCuYPmMrjKnYQH92mt8rHPP0r+68BON/93sX7+tDIXgmNR4Qs9Exr1S
KtG+L6nKC7xjPlUjkAJDX/1xtxhb6kh3Kuxjn5bXKrwVlLSZSFi88Yhe8erDIsJgpeEBO8yTl2EM
xolkQoNkywtV2R80mhoHqLqCVN7Irvvbodtiq1klJQLF77olA4DCX05eW1j8x05M23KVDbmrxX+0
xoDW0sbpFVhe0gh6XCXIzaHdj3LRNreUi0MWv3AzyHT7jAdqm8qzH2WZ7S8vxX3at51Y+V6V0AB+
RtwjoZadZk4c2walPnmpmllIehXG37LVJBznHnOD0dfJp3qKPUdIJ/88z/aRY9GIMoXG6gHG+Wv8
eyOq8Rt/ZC+KAGPv0lf3DGeSd3xplm31g7yaoockUllaLpHeF0NjGybAklQR3LoRL0OKEkhHIj7Z
6t4l5+8f+AudzvNLRS89CTo9Eae7b2rmsowcU9uCKx5JnKEt9NJP1eWvGeSkso6e9P3aBaX10+vd
OchxXh7kist8uP0S59j7cGXIJZ6/ofGHEUgax/ZYANpPsXp57cJwXMJJ9CmCTQS6s/KKUtmxCqXf
226mr+cKJWeF6enbn7SAXQWvVaKivz1Mv0VPqAD8XaE2RvtcsFwtuXgfNWvHr7ByFP+b5as91Jpk
Xt1QfgSC51ANRuRfavqsYDdZEd6cm7wlbkrrMNMDoLf1LQObLl0rFaw6cR/b3424nb3KQZ8A1QUh
kCopjt7iXrnKijOc9Z9vsok3EmFN5IFtL9IJoMdYVhp6mnD3MdqpNSUvNtldgr6d0gG3qiNjLzpG
iyezE/KOnmLQwcMXj8XklnLYpyO8Wii1yehBwHkG0VpsuswTkpk5NmjZEbE1gV7HlKUa7aR99gfN
M6i2jsqUEiE+GH2wFj99QYgV92IQ6mcS1YzK4hcpHl6B15rFw7CmM5rxDzxDsVKWZ6hxv69lGM5Y
kkoeauoTWm13IR8PvNrjxMrAjXvqrUXTPXRsgaqJ7TR/D7KYhVoUIaWpc2kvaL5JrR4ZD1Y/tJEH
A/ciBclIyreCGvJqiEP7I1Exgi8y5RpiH2Nhb53PwfVzmkMjZ9NlPJATT8Ds1oZZ492oZ4L7kt3q
nzanremRODkeMIAePinHaYlegdomuSSP7/CSmkSCgE9JRCWXH5rvgP4rAkDbRlRIrt8C5+2h6Pqd
ZPtjqmBBCeSHhpyDXkWOCh7L3PZ3z1YSsq1be+1mb+3pm/Ba0Nw0oe9Y3HnjUuBRjeiRVYDszQ5/
nXC5MJUpCy5g54kmwLXsBYwhOwPQshDEoad7iejE9R1TfDp3TqTkGEafQbpyWLRdyG+N2sh77iPt
GZ4Fxvh3BdbxDtBXboNt5crUMKPG2GyTHcdt7sFAycC7MGfAZ0803mD1M92i3um/iFI1wpEz/pj/
39qcwgUzlmyeNkwMU8e1aBFvAnitQgYnKidOsp1aO4JHljETPqTDPyNI/KL2tPqDQeGqxEinbCDU
T1IFzlhOaj4tuq3cJttZ2xV/cLGFBn0Tzw/qzXiBcfgAj3QevcVJy/g6t0M+cdY2bcY74OaaxUhW
eEymTVIWbEArkCS5Pdjw7Hh5GkH6dYspDjVv57gNQse3YLQnIpwQm/10jpqaKFgit91X5GMjs19f
3aoufIFGHeyAEpMQfWdNkq1bjva6LbG2dEqfXBWP0XoY4dwz3ntPeF9YsIQxWHRH9OOeqRe1cwhT
1kI+e7mTYTFs6acsLTNrd6arR/QpBPg59mGWwyUHKz3xeTTmkKFQfWpZ4QIG5hii0PX0NbeO/+Ie
dHk/O1/Z7b6OJa5ad+CNGG0nyT55h2QHTjKxk+WMF+wKc4IoSJEMzEgNqOwJj7NHT1tgPXNhGluq
g4teQ2Er4aq8+GbXOGlThnD9ioH+P5YqVRk/P4MmiwJXSYtntd0UMoDYcxMvcKUIOhq9oTZjuItX
2Q1Kwh/XCwFQFWFiMjPRCOGky4l/3FZ8QoLFFBPudHrAd0MDx6fiqnszd8vJ70fvo4Np9Q3Qus1n
rYgjuXqQ7iNogpRPaCDgaQcHirua2Uzfja93x8cWiJ4LrFpofbuAbSlvJoj6ntmAOuV1oYMGCzeE
aCzEVhHmvGiPm/fJY/o3tYqPylEUpi73syN3iT8U6pN+FXHMGeYTbL3K7A83uQPLKe0BxiKeZP42
lzxcHxGL3nRoiwIMYc9tQAYDL32nqrXh+Gq9+rTL6vyrdiwTiys1nXbkwY+dAJpXhKZ7oWhhrrqs
hlhooSKXGP5/lEieShHbFy+LEBJ3J0jnESUCNZ1VBpxENeGOH9qYE6t+939aKwTuhAk4oTxzN7PX
nVg+qf7/GzVIf7mSY/E2CD33xPOVNEj3M1REO1n489zRvvdcaK/hUsCdFM+TbFMACPuSyZacT1/O
YUoRZYKA6/w5g9wUUWi3UW+m4vgKzLWrlp3akLVWMh2oQryWeB4VBvm4F3tAK9RIecqZFTr1v4gZ
Ebj+23iQfmxZOKuQtUCjnMc5BhF/slCOEGX1Lxjv3NBmq44QufPhIwCh6TpYYhCZBLc7V4Nn2ZTf
jd5jqqIa/O6LiQcwMe38ym8G3R6TyA++A2le736Z3wxWz5W2a+ApQUSWWp5lZTRlCNBwQ5oKcMAU
NeajftRqqOEo+t4XLdbRDu5toO0Kl2KXVge3JX0AuakuIPx6gITz+kxkno62ueGTJaJvlY+dA6u/
taJeyjp/W9WUZjGBcyCLL7YqPf/wJTsuLA7/ZfXJoQjGxeGZOOEA7Yh266QHFI/g3bwsnqrhcg3l
oqPCI6yCaNDiSu5lsdCrtYwRVIT8kS9p+rViA2RO6A3KER1y60EbcflNxi46YiYI5i+FMM+xGIlz
ApGMsIgP+H8vSC6aQElHi2txESTegJtTUG3tDJ+uJmqW7J2I0Crd1puwoe/0+vWgZ4JZ3VvD2myo
nRalphliAha7v5EB27+m6UoHe4pBuZFxaUIfPWVSJWq9bQZK0WFAw5q8dTq2emcHxk9+O64CkhtF
gjumDd5MqCX2UUW00Ots+wMEtpvlvUFUsyi7o69J1kQ0UgNZf1JO3WZ3xsLk0LfxA5gPvPfLP00x
SkdszjbflYEbLY1GNpI3RuZ1SOclAaH7b72CHy4hvxahFb3D/lg25BN0pAwVQzmqTwAZJaJHQVOX
rMCcZd5GXW7Z0pwUlE7pRTqZe0ox3a5GMsAwALqDqvo1Cpo+Q439+vpzwKscdKVZyYqrYHw0TbAd
KicBe2xwPicJAwaCXxp27pvnAZPDotslbOVT91rtu4vCS0Vh7PY8uo2FJc6wMMEi3rHPwmBHd4A4
IyUG0G1wv7sOnoIMkxkAyuMznLrqjWiAWe9gCsiuWcGVR5V8FKYU+//yFgrb0k1b4s8K4uQW2dI2
sdJeIW6BzJWS+KVukyRLFlceTXoGSdnUbuQD24HRNy+OwporiCPDUjK/tzfmrbxihXlxH1X/4Rq5
aUbUvr/U/1UcaRostye2Dqg5bv8GYYRjWsUTVmT3COv6cVkT3phEz/4rA4iGYJIgnBESRSD2YVga
iM2+DkfD1A/pJ9hZMy4VUsf+XLLcuXhWqFmRhh/AYf4uizbxll27A5PqyQO2vsbYRKrHyRmCqw0q
L69kJcJJLUifds5tw9Ixdkl22Gc11Wc8EQoCqNxsdcLM7dm8Q123t5y8zX7jeACgLQE0rgSL24nw
loU0+o0dBVZ8dOvTa/wRn+HnWBzbWAA3OiLO58joIRMfP5aS+avnKw9iA9zDrviDC7GNrvDa4xVg
vJxewHlSsz6Ypzh3V43cqtFfS+v50u1cLRseiel9ozdM8DjGSseBWo6ataoQ9FvefZIOOlJgCoj2
HbcjPmFuam/Y70q2P0arlDAIygf1idHy9UxCqE3xAumIMJ7B8Rb+IYYLciUH4gKALZ+Bairl0d0m
vrJBG3fja2GKC4PXLH+ybeZh3q5TEX8lanEPt8JxIctOdvOinYqLyM+JbPzPku5H2fAbHKkIjeTZ
RXgOBpLbRwNHl2OoEvJ17lE2gdhnaxN8Zw3t11Aa6B+weW0TCuM53BlrM8Tp7dsQR6duMAcvN4gE
Opr7eEmucFG1NgzVm1DPyhGoVOA9/j7Eexz0nKTu/aBMxHbD+vQuddg9CWPpQ9ig+OYfsgqvhxbs
rWOKFXF3OXH6PGAZ8c68q0WS2LU2i8lJ6vkgtpCeFH4fupsEu+xGQjeoCnUyKN121pqUwnsl2wc6
MPVSdUYZ8o1dZdS6SYI366UW7o/3krH9WE1tJc7pWXl+2ddwAkQmNDXuBRwN6uvSqCaAIxjr9Ahu
sRgzVpCxnvpZB3G0BDQX52sXwO39ViXDhSBs4Co+3XdW+bDxpXoAFiGuSVNLIwhq6sxkda6XYBhj
IxFFj9qlxMq1ld2vKJXw/BaWVSJfmYAAYfYBmD0m7TmQ/svISJKKzRNVXRF509/BXaDQ16FbSiMJ
d2RZ5pu1Ypv2R3slm1i5LNWeIKUFb+V3IqqG7n+R25O6Uh/ULrocwKn30aDK1TkD8ain+QGzObcV
eLTom5Jf3vqqDmt7ou964d92q+tpraoNhyFJVPI3EuwHTOaWkUosP5nMaxwrcVdDjWzH9mKgUi9L
qjdD/N+cWdjTxGuNLQ4PZ6dx316+XqIhGcVrp6hI6yQO2UiiY3TYxs8wq9LURNNyEuW9H9K3nzTs
s81qVwd8SEXmCQ/7GoPBM17oSZBDBp1l6MMbbh7/hXCiLW7+0erHbFNpYeW8KRLQQOEXuQSTpnFd
AdBog0X1tK44HPGLKwY129vGT0y1gYEHD6JdDrIpxmfjXoY6QjdjVksy23ENbHg55qheJ6mrI1z/
Q6g7uQvqTBYahChm1JJ18aSP0EzT6dLWBKfY+ZJh7meoeXk/RmQnbiqpv/H3tVYA5uQn/Fn1Xkj5
3sRnkmpmp809YWOR7H2+fae+q+X/24px7qA19cDoZ7Al8AvR5zHk1rzkW2iFZJ4QyFk2NFre4YAX
WMrA1UScMCH76TA4cevxye7yoQRkWEtsrBv9z00tyfgyjRO9sCXETIixid8jBjfNhKI0O6Uo6/eo
K2sIWaqC3h2G5FS85kVvgm0Ze/WD70Ip/7bU7GWjLsJv9xOkoYsd2kx+9tCx2g4rkLBOcAsaq94F
GsPxZl0lhxMZcex6BT4tSkpgvag1JDBISqBLaGB2tRUTOvABBDqXiIDsSjvvfA89R/sNnEiLPDEx
JTkQiv/Oxt8rEmXPNaa7AB/1R6Ry3UcR+Isaq5KhVfU1V1RgXZFC+IEYvY3OCuKHB5tvmGAbkV9O
w15zjY4xQyi3iJi/6s8InGKe/jLAyZARMKFd+XHlvZoq6adMpsVlh2nRQ1f3C/GcLa0eumHVzOMY
voPsWtbBe9wygodtswWAbP4IhZnSGwmUn9T8uUylOlX9LchQvQUXnjEk+t+zjXBKe/mQDQ1/Ra6a
kpGpKt6lMYbn1avdhESx5yHJ4FVvRhfHs2En/BGhwWq6M7GQyhZvqJ2z6tZZyek+VCPS1g8JIHc/
AagdFhDTOQdByaXZJEUpmF066HbcL8RghdmV3kRGK7/48HAIJIwVdI1C82+rrNg/ow4Xd8NsVQ7E
9KmF6dDeJs/QDeULy38GQAJWZOUm8nobe6YsrhSmr+0k12BSpWQ4IrNtRBOhkI9NfBxCUFyssDhf
HXpozUAbBwZeR3XetY3KaqxU8zx+Ttc4TezCveppVs1KXrrb4CJkxSNUFBGfphnJ/X41FUQdI+yI
g2/cdbC8HybUrFbhp8dB8+SidElhEP+t/LHEqF1KMBT3dSyqCY1SeuyUz1wi1AzG077BJBZ09W60
Ms/rGotIDOVnji+wsyu2krhSOpT9JxSxbWZgD9wZH64wuFNfBOOC7wfR8ZLb7ytV4mljxuippBeB
Awy8g64OQUw9WgstufrjED91lcN2y6HgBLYpQNnsSDvyPbXsA57ht17IBkhW3t6Kz+V+sjD3H+co
5QejWrANil1SsH0x94Gwu0HUxHv7V2ao2FD5+i+T9THuWER3pQKED5ZIdqs0iXkLAJiYeB+qhbZD
nea9kS+puWfwssAL0wu12hXo/gA2sW48uNW5LFtRuTrem2+tMMsyBixWbua+SGnut9f9K5ISg0y/
8GzVLINsjFLZGm8xL3YyyJ8jCWWboWbR71KYFv/MxbRVDzawpCjrH788SohNfgF7OMvt/XOzE0wR
HXQhWKtlByHuFWbO5BjVPRP8NV6q5cfYHPgvRney/zMKisQ/OOzrO8Wg1XD7tDxAtyF/hXaSoQa6
ARTqGa1f/FUhkX06WGpzHSBnJe5BP9dRJm8SA4zMfFI0UnX/ugKQndRrq6sOiRd9zz2Lcj7cZBln
Feo2kV2HI+X8qVhp/mB35WiImY+BETB2HXhrQwgvK2BcToIAK1vGZP24ywAoxPc5YOZIQ956EL9A
tjux2U40FSZkfoIaPP2UedjtDDN/Gu0BbTasCft0Gm4n9qr+4RTv/6rXeQyJXeMi9rtIIh7t7Cs3
OcoWsQ15IrIWu+gvXP3Iz4bpN4a7d4zvV8D0enRvVTw8SMx+T169/G8rz8Kms86+VXLkrQIiexTv
1Gn4s4WdQ0E4B4NVZjPs8mZOlnAncRkuRZuaFKstrb45rO08X8Kl96113q6hFRDfVDdbviHyvBVy
i7VUkf5VxoRxrPnENoi5ZOrr1wtzeQamt3BuV3GXBBRxJJi5tAb0LBOxS3cptK5pzdG9gITvusQ3
90d/4l9ejAtYR3uE4oxiSAgHgSMTduVXBkxy/1cFiBawmkUBA4tLLStGHrMHRS0w8qTO33kr+P6h
p3MF2tfjpL0kFrbSO5cyUZsZJdXax+vvPUjUyDE8eSiLZeNnQe39SlBP003vVal4/CU77PQgbkAW
H52E9P7qWTAmVG3WGHaKcSfIFPwFL00fs4hN3L/9c02ey04sKc0Ed1bbNbFMGSoV/ThM5sYkBa/V
D1upv35wSjBaZCVBublYdWj0U+E8U/BS9xbYICw5Tek3daUdFYtpZNo8Ddu1tja4sOaEsVUfzvqi
6p3vVY9ilsDbV02aO1dQuGts5o7bzrc7CfcLOP1HkAibehFpuSojdndHIBQRPUCmovSeEItkkZpP
OP3MsypgMiB0obMn6EjTHN9J60qX4Hs+oTFzF8JDjOxa/Hrxxehrh3llwqaYYVCOJbfLIpRQtyeL
ZPxE87Cj/5J/wPtlre+BDbVGI13y3a7jDtT9pGDbY2dT7F7Vlva5IHBtlh0nbhvKoofGHzhZQz/7
7rnh/0Y+RlQdyonkbuIjcAAJpQu1vaUHn1Xd0n5zEbeq4ArVsg3lHOmRp+K34VkILUTNUBwSem5C
UrRUIhwQ/+SwgjdEUXr1+ONX1gqHACP4bJBotrySeaWPIv/R34KPY/T4Pd2eJfQI2ccBypr4JBm6
gMWGiy8W2EN/59zz7P3PZodfxsRQMpaM0C3qreZKSxJk2NYdy725PxozQ6QhjH64WVz9v6Msqc9J
EybxJlzBge/zsrfdifSKrFXXsNcdA934buYnoxyDZe+NVviYHbQREjkQNdQxOoOVKa2l0TSfJuSs
r4J5gv9EHD6/dmGsMHyflndpVDFjCSutKZTCZtckN3CGL1qxwPWZiJQZFD9d7XSI5yg+PhFsPFz9
mXClq5zzkNPCNZ12rCtdaOY/TldFNnlDeGm1QA65w7gZqWuyfotPUZ6/nrVDmxM4jDXLKPsaOum5
FkEFWm2SABcpom4cSGce38j8t0UV/DNBIi2dOR48dPmZe7LxVrKSzt9kLcKbzrEKy3xcf5MKF395
jWuDjpkeAq9fmIowER0PLNHV3D6S6x+p1xuXDS3l5vVQFwFV+6+D05+Fun/6fbk/3yorDg1ljmYE
HNnpZSejmc+s5sCAeusbDRCq907XaaNDUuEi8dFU2hWbMh9qn8y15yT+ypCJ8e5vgLc7FVIIufRW
VXf+qPvLIpDbq4LuKioJjCQiRhBuryVzUl67eHnpKCsGyqXF+hX/9yzTdBwk3HOwehvizoCVu2er
vSKy/v5LtDxiYLSsMI64G35FJ4QU2HGaFxAmabvTxJT21VVp2zg8qR9yHUlKfzRHwPY2GPId5W4K
bof6J4py9PQdZBafM7yEWP5BpHwY/6OVZ6tqghTTlX7ECP73iyouqMiR3lomBvQyfj1V5VQLDKxt
wINB8gKOLh+Tbe8EMHEwhPUtO146jeQb8EpCkyDkkXdERDqxB/tTG0BDwbx8qaOxLazjQI1aIaD7
qzELjKcvzW1GooZAEeCghrKLf2RPtlapskHrdaOUHLga8NomoqHovVwa8+6a1b01WbQuXj5Xi5jL
otB2fu2x31Pe44wzzk4UbXe3PtIyittLaz5NAKqSvxETgUldqpE9YZaqG3cB7jsE64XNCE2s8FHF
3YhGOD1mITK6aPAv0bxmBYtjQBWlMxnAcFe3F7vKfKi2VZ76G78SZ/ajGW8Ww4i/BOU4mvNL0lf2
bth89H4n0y6NuafyXLX9+YuXpSHR45U0XGLws0wQ7l4ET7QtzDAZNvkiRTByWTHpg2drDTcT3Qps
hyLMKlXcw8s5LFRFTg6jQlfj4kXb8RSVlDbq1olhSsXO3vpSJcmTSEGrwm86BIPZ8QEX4bOofUtq
4CBDvReXHPgYZAH681bR8cyEkMzn7oDsMwd0nMUYQ5fGWaAk1oN0EYBWMK7dmbr+vEtBVuabXXAM
5WjeTTFY5ooDXE9OzazHFBnrzstQdAL4DzmicsqLh37Fg1P3454S+Cfq86aZ4e0v4dNWf4Zzslmh
SiFxLas6HljqBwd/NuaznxcCtlryQJlctce40LrYLLd1Wk7zS/xPaPFyvBokO3+CYqXV5IvVN8t9
n61DEFg6FxSL5fxaf1JyiY6ajJ58INvTpvagGFT2yeIgxqmv+iorR21sNUCvfw3FQoM+EBVhZzJu
k5k+bxAmRMRUhHkmC3xxoH3OLFVbwJdnD8uKSFe6z4NBE8+vA9y+dI7eHxk4FUKBWXUhtO+3TXUn
1xskSvD9VeHDSm6XCIIVV0YcH7QY8WfsQNTyimeO1Aj0ku8lwCowr1JwTBd8SBiwxc3SqmbWl6zH
bD+87ewH0F74YXhc/aBll93P9xFelR/04HpGysD9Nw3AYl2B3g6RDu9EyCRuHp/JTz8Gj3MZsjw8
17U15rnPhnkXvwwXXeaIhJKrXzGcUasVv2CkvuYE0eci+2hn38oCsfsNNy2TVzHoFPsetm94SehF
Z48Iliviy4jalwl+zgT/aKcyyRE4cHktQRxYTSdBr+JSx7l0Gmw4hfLgRPlWryofzLcBQ6mKANQJ
hyNgEc/B+GozttZ2pmxFxRuLwI89Kh7MOUEQ51SjbaAw72Oyy6ZY45nbDQMSNYE14trk8cniY1S8
YpuIxoOs2SziCUxDi+7Go4dOvTqC9gqnwlN2GydXKERrTW4UcDSPEFHVqrfnsoBrSJMsNaFP6M09
5gL9avzYbW3I5Go7qn+ToaKYIKzcPQAt5T7EtH9Qyvg5toKHWhrYNzIS2fihvmClI23QW4EMkiIj
FTzkbdFRn+UonBu/nE5E+IlgHoT323yHaAlhjVU/6HRqV9Gb6REdXRMgxKD379zbHcWpC3shVL0h
zPiaW+1UuMTY8b+3xy6i3hglzqx/N1b6AgHboV5PxfXDkmgIltqsf6iBHxlqq8yJ1GchM/wE4RgU
QdwMyvb15PR3LWXi4xXYEv0aoqg/1Frr/JY1BiowHXetQCGr0OnXwF1YBHfGPSK0ylfKFcH+J5Ru
jcrP8r5AqDhDJp6p0kabSIIrNdxgInjVC3iTEXifRba3Sp3GLyKaAH48hdS/Nw4+j2kjPM0oce93
GjXHnuH7GCH5uI3EYiGFjGHxg2yzfv/B2nyDaoztkLEoJDyXRUbyvjHzjEBhQTCItR6+NBUk1CBV
acxfkIFmNEMdnsQKtkxPl7zlhQ+JAKC2/IC3axuwt5D1bs7N9Ao/Y64AgKs//oGb9yVUc+8TRXsH
CHs4Zki1lliutZ2YAV5ACZUZ7gGG8HKCvAj8JKNpxj4uh8AGtJgAJPn74AIvEkdhArLUqMDcBtmm
ER81HmGzL94/ztHo94sJW7ffqv2EHfHe2ijkk2JXOkMlY6a8nuCGTE3ETPyb6vbLeO/Ol4lNO2d8
oP2TLEwVuZpmQCDfRf0dA7UqQ25A7uHWu9HOdnTix5uZ4sQhfKePJtFFuYA28wrNdIbsMJFUUIg7
txof/Mrxlw/0kI69v4F+KWM8JGw6X+JQiNY1NLeIJTm94Mifs22dqvJ9BTKJNTenu7dBLL0KOUiB
VOvqdD2QTUWiRRaIGId4VdG6wyc/6qClZu/xstEA7GUa30ervc6QhivxSiNxQnjsYDDL2r2qI8TX
0nZURShKB8atFR8Eb6xsgdSYjAp0ul11hMxFM2IAbAtd47Whil6N2dJFpXH+glzJO4vM4ImFaBtZ
o/okFEoutpKuZeSzkrtnxDM8hq0BbGtKfOgU4q+TszUr7OZjvZFj88ABc0LlJg9HSG4cWagcewLg
MvZCcyIv5o2sI3ZgnzMJNoMOzRX4jEuWNjBlktfGs5ue1CEtQm1cbs/Edm37vE69JAW0L3EdDEQy
ArNVerHnknlsm5RY7WY2AoiywWjMPAX7Awe9gQ9upyYURJtNYPUWaf5uVtUsiDIyg4u+gGGDEWZo
P+jy07Qs14oybrq7NfInB1LApKqqyqDmDXcvDOSMRnbrHqd27XWNoLufFN4wDJGXrAxOLlsAoUeb
Kj9Fu+9aq/IbCAy1ITTO3nZEWX7EzK9DsEUuS0irvlNIivqqdiFwiQorF/XP9C4K2PDy2wuMWg1h
eB85o9ZIINLScOFDZ4m6HMWdRUH9wawoDayG4sJ2ycvpxC0Bxs2o/AsLH1FHjUnyHMZRPD9xVXFL
5MnL3U8zspO5t0KOa2L48PfoFnwmRXyq1GsS+AAqvM0uT81rvVZgR83gUUieXgdx9+YVDr0T1OFv
50Pi0tdhr8HiPsKFsrYPUksR5VIkDa0ykdcGvC900wc4+xxTECMRe9Jc3u+28lA0RLZJ4IRRNqc2
mh00plBlZc1Wl9UrtRMolg/vARYbzMTIDueLi500DX5QO7fxjFR8ym+vzvwAQHMRwfGtg9xtNSI8
CZAOFuGYyn5IBhRhme/u9uF4kAal88qOcj9aTnsAb/Ajt1UQdVKl/wKTOJyP+GTVUASAvE6GmruO
eT4uaBvfy+sH/a7/zwHRGORMadXOcQJmTzex4SgowtO1+0VK/HzpWprTnS/a1gnZiGoJ82WHWWXM
ENP/PTT344j/QXLBha74kwO7MQA4prDZc2sYbcUD0s7RFsYJ1nNzUcYapuPRf7+j2fnQw0xGL9or
77/O5l6qmU/KCnl7MvoR8vfhvX28SQJ/9eUplJd+qdwrL0lGbx0E/Pzk2ID8eCnxdJMQYhXU+tlM
v4PCfO7XfrOgXxOvhEqAOtpZ31GgEugn23cLN7hLFgSCZMGvPmJLssuMDnaSMajfKKd4zJQt6SzF
xmjMd/T/3G7CcYYF7vASvfsd9x43EmTpU2It20QP6uQr1f21u0i0aGc0I9lxllT6fnUdACwKHCfk
7rKV8VolXBTMRb0Odbdzdx9PL9y057b5DbANvlJUSbGPFhM9em7j885sFNvCzQYG8aEcxMerj8yQ
xPW7EYY181HA3+JSpovC68Mgcsf9yBezyoIiBZbDLUz/sszJsa7f9tKEtuJVOkE7lkGsrsh8FQBZ
77PYhpaBcDCrNGv5XUl9n6/3rj+/mgVp1LV2jodhhZvOHXjYuHLBHGTZJJyof5P8nEJ3+fzNMA27
m4lQA9WsoGcAcYvSw5OmgN+9WUkLbP4JYWOL76FCutv2DGbv9EQ1UjuisPY2S/NSi7/Sf8bM0VY3
njlbJleRx9DnBH+yyzgFUai4Dza3sRNLBkyQ3QNkaEztZg5Dqj7BkwhAaMbbOloLrFUXD8iOUySn
ZUR1eioORBcrBaKehGI//geDC1I/JkCmPSOpme3YhKO0jf6aiQWWQngwXhOvajvSigpaOKc2QsY7
MEwZdbS88SmAf1+q6NK4zQHk6HmTLY1pA2g0HNf31c9hjTP/dE9qavP3qHCoDuZLnNyBLC/+yntT
XgrtRjpQDew+aCzi9kfFmhzEINgDBdRQ29V+vxt01Kvj1Hl5QCarI62j+lBRyuSsxavqSzZOefHN
Vbh758QSHU9FDqHVqc5EWGnxZlWKt5ovULvug8hNYvvshEK0lXmqUCQ8kT0L/I+hkCq0HZ11X0wG
E1uGaiNtdE76k/PoZG8of4nv4A63MiBekNE/nXLT2N2NoZDvTA7N4Quix8383KbrUUnSsNBp+coG
ne6VWK+gHZYPQsKpHwZIcwxW5jONI9SxJ7ikgdySTb0E6XyYkGkXsJele4CUNXiyoS2z8l8i9gGL
9GNMHkG907S1S4h6nRsJI8CMkCsdRCI/ENR+ZuJWE3MP8H/0/0y1PZhrHby9dGIafXH+ap9t6NI1
LrD+0Rt6k+LCqKs0ypLyzckMUJ/ggXngImBXJMWu1OgDXT+On+vLkJSAfYio1tOAJ3FhYHBjD1Ts
mlih8K2pYZV5VTZuGowGi/ZecKJME/R0NwPqU8F0hsQqojZ0aLMP6XNIRRDgwi27DMMPMwaGvo29
yBacsYibx5Z8BJGnLjX50TBEo2fG3C8UKhOFkU+jQ82tgUNVkxTuNavET1DVoikzsS44mJbm08ua
2XcD74XgtZ2BhBOEQB3Qpmuq/QWD7fEk/6ku2JDRWj6VZyUYCCWJdQlEjFrWgjY/E+9VZx5MLBGh
WqgjYypk9tVWt1CcOys7hxx1pWvJ1wNJLjOYmLX0UkkTX6yXeevj0SFRnmSeaPX2kgV8jE/eeEap
vUXpqQH4VjJCPbtBzQpdazMoaMnCj+VYQxwMCoLQyhapVrA1H86/qsAFFQvbADHnsbNgmrTO8wUS
EqYwAt/UP0nhJyEqiiWvRNHYkklsTIGaDDWcCWbV1HOMjfcvK5EzyQL5GY9h917xBBC7U/NI2IZy
QWacQQhm3u4sPLJ+6OXtYa8AL9dUfSmLLdVfaH29b4ruR6Mc6y9YdSQ8q77tJNaOysTs5je0050Y
m/om3RI5cbJ0ZSclUrD0FjIerAf2gu4l9XVelwWm1dQqyLMZXw3j8hKlYlJ2u+/kUUhZFSooctAR
A96HzVLFIaQyNcyrwP4cnj0VimapJJzfwB0TlaOxk/7QmAMn5MHX0gVfdywy0K3aCJY5Lo3JWk2O
Jkp6T6UHwbi0o5Lqm1x1xsIRXf+c8sm2lsXJpiiJ7tQhEDGon4WsX/EmcBDworMcuGv0/N2C0tWj
uqdzcWboIH9huKmYdrhEqt+zoE9cSSSTw1oSo0+M8fOP4joDjI3Y30VXOnUdCi89TFNA+y3Ij2oT
4tqRu+aPIFPMwka0Dz80HRtpRH4UGHPQEQfoH3AVX2tGk4gR9Y6sZTli8tAd/jbprwI+q6XdyKAf
wIvmlX0pDoRNzCFWaqiYO1iPNTdqV1KJnsj7TvEAjbJNP70ffze6HH382ppD2qR7T88bAwLE0QcE
55rsfYfei9c+g0ynQ/7/bqKYbYoYDiHiGCik43VDj1UO8Gm8pZbraC9WXotnlBToklc38ftAyjxe
uLEvHyPHKMYf9ldGDCKaRSgGWMFFeBprWidpfWCIYzUJ7rnDCavZO1KbBJcrhPt23n/96qRdL5TF
PRyhaqMeXmaFoyigfK3vnGV37tP6Kv25H5TTz3MI0WZNsZsaOBgZ0Fg1We1oiXjr7Y4KGTbyMSvG
4U70TSR26Fn3qgpPBMNi/8Vvu9DNGBpOiGomOOF3XvFJIXqYyqiKYmWkZurpIkWA8aa7aFnmZikG
NaT5wXToONQhM0iZCbfdS4UkE/cVicid5P3Q5wExoHo6+fcT6KIPcivp+y6tWQeQoCBkGcd55C/I
PMZspu5AoljJgxH76FTtqV2OhfJNcfoAnrh3+i5S63wHOqF0BpTbbXJ9r1EMsTlQjt+EfN6eJ1mH
TnPhlLU5KIpUSyMQndA8Tza5ZV1VEU7B6BxI1S4riFYSNji39Mj1XPV4hbwAg7Vxpo9ta+/6C2Ip
Cs5iC4Okzvwpv9IPEGmQrBxkiBYmrz9ZEbLxfAePp38iAuYZExgX+XytbQPWdvpS0V+YWYUpE1+T
CdgK3q3bOluGXDta2PZJD9ZPBJP11JrzWPj1Z9hXXNRgOf7vXD8NNUHuSIRKPmzSfdeLc/VxMkEI
aNqfMFbNge9Ymh0GQtfKpp5Ukp/08DVOumz6NP2cOPUXywZP1G3PsxiTNjiWRoq1cIReKqI+wx5f
18/sn6sC0fxi8ko14sQIoVxic1yMFAUzu9wbc9HLBqf7/iaoF+uOn9Uey9cgimsRs+6bjpPl78EL
aSB1s5sTTcWIzEK69CfFs/tevUFsEVTyv5abcwg1QXCVvdX53zRFXiKVBMyhZ2KVyPRM84GqQREy
BEO4MV/RTxtZD9mm5T/EbbDPpiowwyA5XVuqJBERr6M4tgao+iGtfi8Vb26ySN+okPfLU40Mc3DB
DNIZGUCBW8Gq/VzCQLuQ8TrZhz6vUYVt33bkk1CSS1+Q+hv4vKzibDkNTDVvTmOO/RubalEC6YAk
w0TTnbAHeb8dnKHlwwFsM0vrmLmVtg5Kbmk36VrY5R1XWlZBKnj1LVMmNzB3zkaR2U9mEAlUedWR
DWcFF3ob5GFPfAZMeWmZaZiAxWr5HafU9EhqOqUo8Ciy5nwNYb16YVI8SddtcUiOqJuUMf/yTqRe
AuvrBZ0uqKTW3fe7eZnS8c1HLYh1y0eJZnoe1RXuu8Wlm5kDKD1W7kauCGfswkgi7w19xcb9Zpxl
A4EW5ht6KR9d3Ln2sIP+iq6MN6UcLJ/7YNhnUFdHlQ8pyFPgHePsdA4TI8RakjQZ5yioXXJ85fkl
d6Nw26PA+DOGCGBYO35FCpfkytZSYCVvT+RzoMo58xoPB2A+EFHku/ZHLqtWZiRJE+vNTnByteYn
BjfOcFr+hHzOVBl+180dW77YjoFnfB4zQHSDgKL7vRC/QMket6G88cxff4Nu7ukXCyIlSP5ya78D
0mlRFBUKAQZtYIjgo4lAt+uemMYC+305ly3AKF7e01osui1bVdiRMgaCm3YHsttQVvOsuULBuGYM
yeYk90dOD2RZaoWLQjB0dxpCAFTNRUdPvt8ooECbfhFp20u+WqaYcIu2L7VQ1URdk86ZB1lTyJcw
TB2gJXOaiZv+RuT+ksb+KGg9c3McJWDWSB8go/OIcMXLWbOhScjTgHWXQaIAR1IZxwgZSVu+uuHU
bvl4q/ivVHVuHwjcncMhnHHNMqj1HaP4Ktnp2LAgEybkiexWcjvQZEyCoEceOoXXsy8tMkQE91qQ
/xInejLwx8FTCteUT2OeFLXVQtV9Fc7uqGf6XL+svGxBJtK2tuMXCzfvTu60F9jLeUVte0aC+vKw
o0scJefkTv2pBTuaakNhJJmCIRi/jjPP0NjqxseIX2d9NdXCUMbBGi8XiHbpOiyNHusImFB00Iqw
hYLd0x6yFDa57aRQ/No5yuL3FEXR+abC3wCT4HBqM+42N7vswrL/yVOf7iJFxu2yJZunC4gkxtDf
Snevo0KduyLlh9/VKBDJNEEos44XgPFnYLdrtzbJ53wpR15lohCGskKkNn3NArY+xg11Pw+nXb3a
LCxBe839fsCcp/K3MimbPSaMPOqeq/nDhUdrmMb0CPbgZ4QJ3r9k5rl/qM5hmeHFEGy8pZizDJrk
EsKRdM6dzlWS0rbo5DLtsQbLuHI2u3k1wbXMOtt1J0z4ezZtWVVsy2BczS7hDp5NMdKRsgeJNpph
DKMx/1VJDYt70yvFta9aJdUqmNP2I7xtxvleg7ZgP2t3CTZDyRUF6fHdeU+7tHld+nnHDVJh/X76
+JEDbfXEMH97mUN0cvkDfgiY8flspkDAEusDplFlcA2GipQpCbOP8doLjfSPtHBVaum4/718hWWy
RHz1PzT03DWz1PLyDe5QfduVBv2TGwEnQT+SwZ5qmUUq9Vlc1vvRSbsXCtjQxWsF3Ee8CC9Pkb1I
oalGUmtl4wLFzCuM7LR91bMLO9hjXO5wa0yJvr5L+y25HbFnIwA2eaT4L1Wnb6a/lAcbRa2sw/rZ
EtUI34GzaoRVgz+NE4CNKmYcews7rpcID3h65G6HE7n5X0bDkGxoQfG10QoWHG5DvAHrZ+m2QFM7
eI37/cC9RzWbchTTlykorW+JudHFLFd28JLVmEaeW1a18+LBHZ4ZdxxsbAske70NdHnBNhIunr+6
5qvGPbiJZGwbxSbejL2rpzMKFZYTOJP/X5FSGxi8otAPNVATc26M0cNgQ09JRdS/cJ3nq1iV6IiO
3zxddrGHdDO8qW7TjQXOX+rK+WdmKV6tGhqA6cLRCYmmPuZ6rI5foqynW2fUiaNU9JfmNEQs/3EG
9QFvI8lOdfqlhrxu4cPp2i6Soa1FMAOrB7+ZkC4GcnEg2hygvA1AJxzx775ReqT4czYRE7gYYZom
3umsn3nT7raLbQNRAAXIR5gPv+QMYTZXeOSMkBblOh0z9UwXHKIf3MxA8hcDZ9Ycx2aQFhCukxg9
2IOsCTZRUfwln91B2QMNZlSbh/U0SvhrS1lIxlDWk3DStPv7xkdk/xx+JFPXCQLA8GwjQq9RbKei
evRMVbWJgsBOUyNQf4JEnnV69//lspoNc5UCCCa1Gjfb6jOyqGvE8VXlxXZPGYm6M9ASG0TvrLnH
wHmI8iPPtbTK0czJ/jD9b6gY84/3zTsJ3j0MtRX7qsGWZVNTkA+8aDexqLVA4hSvP9rnrVOnUxuG
ME5Ma5s2WpdvGQDRLCdIRzJY3/waO/mLSH7PacezdA6JoOnskg8fiZfhLS8/wFaSXOgupSU99w4t
B2nB3Ko/P9AYVCQ7U5ZGrvxcU30oWhmH7j8i5F3XiE+yy9QwWmdu7pwolY0yfmOlF5uQhtRPpRwb
e06e811i1XMbOJrAiNjE5Dc8N20/4LnVWwB4jvLRLRjbejsqjW+lyCOGo7imJLseGWE79mcwvcpB
KExC9Gp9p0dSQxgT2s5IL2LPovpBp3Hhxm24g9TGwLYwYrFliKhXHN0Ux1xQ0KCQ9X3AuJDhtBvk
BWEyjnZaJuHRD47YvBkC+KXj9ZnTn2yOXquEAwfutcsko3TIl/pj5IJCvB8J+bu9Mrs68ys96rA3
fwEiSsyzrGVUFLIyI5lfWeNkTM+olVZPOv4ilB0z0OP6l6hirfhb7Kr2k8+9vIWDqAdYUv506XyE
VxmRjvRRkURjat83BReVPriJO8m4VWmYeNIRqniEMoRqzoh8jCerunb85s9+DPBdRZCtu8w9cQcr
4XA/7nA0RoTGUssclpVXC4Xhs1qRAgMEnEwzxKCY79jMKX50WiDJ084DIPOXDRriAk4cSNZbjCXf
Us2SkcDvctAZ79gPNiZaTpP4gUcsopSModdWKSx/dftS8jijI9mlhq0BAhU7dFPaFCHqVJYxm3ph
P6teXWE8BCCxahn9JAQSRokIXarzPeU4kY29f4v7cluGV+ILzBjUHak4Ojn+XIOTa3370+KGmygn
LV9m/WWG5uHpn9SaH6SE0PYv179P4Fb1LtSTzw1SyMfOO6hoKoKpZgmVbPsthF+OGJdjeD7n04zo
WrhMOguBA1HsDEptc5zQWIq5qeOF25OeE9z7WVKTStNZP6S9PXuQJXKC4VOspNW20mlQhUPzjybJ
m1DlpvK4QKzMA64f7BKTzUTv1LBXp1YyAJC6jW3VZsfEOfl+P/mbDQDtNdjO7L9TcilPWX9USTAF
/tGwGfpDJkcFECysKQCzqoBnx8fZF6AFqYWSWyBgsWqFjv9pm8ZPcVfSV7AUUVnd9HMerMhngrX4
NugRgFDKvsnOXKaJ1b3KFhGBjXf41QNzrDsrtuJEmWY5pzJmIXd/QbjfZQG3mVqur1VbuFIPeViM
JeE8ovYq6DNzTAofEaR9e1zRk3TLRQ22ZXY3jLFzEG5Nkkm56dF6YXFKDnnXxlV8KluvV1ahr4KC
VBltpllyeTVwoU9hIxq3sfZ/DJK3R3sLVBVGGjeVRn3WfBdlHMfhfbOUIjj8Tb/aGDrnpSxx+6Fo
g1enWTqLYpG1pthhfUE7LhdpHiUObobncGbK+TwX+FpSIBhxZKnxwfZXXTaXArHbbUVtTgexxfTF
O22eQBJRFlTbXogipFodcEYy/JyXOKsCuWltEaDR0uPMznt0CDpEOKKHZrtoCD2i6iX5DLm8Gwbp
4sjyCIHrG2bxMhmczzFMuQOzFgE/Re7rCs3g63Y/waq6PKXM4DX8rrawT0RSaihsCBqsFo2kvU0M
dI1g0HPeDGCqa8fPy4iZtcDh7Ub8C4DMlP6+BuHxxFKdcihK7LPcv9AI3rorYfJmnyXV8OY/Rx0O
Xe4YWiHVEp0vnUrV0Gn6r7Ye3Vq6tbsd+c32Q+c5VUX5eBfkVthkbOdSePqqkNu/GsM3wlH5w3Lw
T/uNW4/ob/fx1jzVI7VZR2grlM+/1qWzK6W8MRTRST03nkVDkAruMvMK81NN5lzUaWNTaa5SIit/
CDbbtkTD1FMSpgvN7iUysqI7qNnGc4AL+y02aKvNyGFTJkG83wyF/9jX/xjFrj6lvg5YSA7zE0WI
/tCQ3z3L72w8FxGrOe+gXkulsOwwVwaKjqriB4jHA48zHDKC5fWe0nncUf0LMKNNbP601BHFIeMA
zwXNni+7orHH7bn1O1PdARsQgHDpoofJtCrEFKXzwmX0sLGfO3KE+/nU2kQc00ij4sykkfPYRVWR
8GRiNyFHgL3shx+RMSmkKYLiJQGYBJsPToXSz1Zv+1Z4AT14juMyhRX1o3dSMPXMhLjsA9QIprdz
GGaoAoW86TUCewJGPk+h4BCrUatfy5oe8evxLIJgvqga+G7IWiHLkeCa6N32Dke7Kh6486p8pYfg
OFXNDJR3dC/Ib1ptBo8l7eR1bjujXqFWQL9T/5xZQuCXNiggR97hpOHOurqgL7kdjzYw2Uj0l3jJ
qLtJH8Eq3SJa2vLq9m0wO+gfzFMWbRYEi5DQOK5g0pqgZqL8st5K3BghcwB/4Zm/ysngtOEce7tn
SVmbfTyx0Fgiz1UiZUn5RiomAhF8L7TYe0/2zto3OBm8pVJJv3eZq4Nt3jminNKkuag9XEWGkB9h
LkV5MhOVM8RbrO9fUa+SKZVVp+RTkMu8mqgmlDvCoZLzfCuqBG05J+uBro6tOCYNxt8w0ICp5rfB
IgJgqwKrgs7YcPwZZ8QOzsf+SqX+BPEX6t0d1e5CtwQ3zMZQTArEFF2ZzJu4lmgRGcWtdBL1q56B
ipTOqDtvVCl+EqWRuWqWgY0KHgdXDWsvIbdHSOTxyEEtjcQhDkIgM4srwxwa1bfmTfiA4ZKIz9F2
CJE4rUhOgKmoLt/1SAyEsGxWhPa4DBIXqAB0AKATFpk8g5/OtiDx+jQMpYzS/IBIFgs4YCQ1Dsdh
jnxAXvZAxvCfjd3VOwBj+rj19CoUgnFv4lezUirYLaR8EdSUOSIOCqPFYa7MF3Jv79aP+2OaVTY4
3B7xe2euuO2cQcgP1xfUH6a8Jmu1MMvQDRo02V21SKxEkVY0sSl27EYdVrW3QSi7hCP9F8tXgLHL
GYPdLXUFy0MLApveXAwWteVuCHifRcEV5xPalevAv5bYGkYTmjWrvQMQcuBmtKPs9MaLgMJ7Si/j
Ly1xlFy+9oZxciyiJx6yqKI8mVzVGvuJIsCr5AB4+n2eE29ajzCbKFkHnjMfb6X10ZiY1Ys9YsKk
blvqj8yQbBP0BgT4RyABSXYdyXMAwEKpiIi5JHDTV95FzcBOSWgDBvV2l+P3mWn5QwWCcTY3ap+T
4889o0cK/wtzeeI/ti8q9+43gXpK1N/ffNYgnCUMq9qGJcCY16OVjWgVMV9G3fPJjmo2ja2CdHjF
1pS/KA/FcNcLeSar7HPrAlN6VPMcFQtqMOoaUQaF5VdSf1IFzogSR3Wux5jlZ/1BW70YoqkfsZ00
38BlQrE5qaPVnLutsTtkS3Xpaezwzed0+B07yAJYAKwKls4VcIPXuBYhMlkz1aDDaRuS7hlftJR4
R6MFeQSDNC+ZwUbTTHCZK+EUuwQhmIRaJyTvN7XaLeehBw5l+zO5SyEi/ZyEHdnca3/l4wyWYRqI
eCInCqSb8eal2aXJlZnIEOQ8a2cF7p7+HUQehtaVl+rRNi4ZGONXfSC7dh3FNChb5aZFektpbLwS
KxTWcA4aoZ4UvFTdFeTFxPgTSGkGvmQjVYsLeLKuXxyhP9XEG0zK+pgpEpwX5lA1+R3j4Kc1ZaGj
nSC6NJeZkN0i7xJ3j87RFOZ2juiGO+fRqloCWgQx6oS4LH9U40v0m3ggfNKKrubTZ44r7f47ONzR
Cf2Jn0Tn0gULVVUVwgDkGvOnO2jTFLblTj7NFR3V6s9goz/6nyHNKBgeu0mo6RVwODqUeCSTvm/8
JS7JKlCdyLndRKzVCh+LLussiR7fpcdYuF4M67qMILcTO9y5UsMWPUYmy9zqxCAqk9mk+y7srKbn
USwjuqb5bMPCImQBi9UX6OABEXPjAHlm2IRgbRIzSwO/BXGsxSU9C/L4c5O+weK9mkDzyIrxA3u1
3flZdyub7EEvhfzB27dET5XJ+IncjPxdGZB2oy51pmPOs/R+nmPsG3JHmCo4p5OWmhjjqD/+ZlJD
8RHNVlFYvHXVlEhOhV/S80uxd6PR3hrIo34n/3iVk86pib8o6bXs1pB1jiAKx+/UC0c8Zhh+5JCG
6DWiYh/rrcc8uj7KTtkSBjg0/SyxYWUdxDd7G2av5n1PRHFRvf0LzW2eCxQ723cy406SEIipnBE4
tahx6KEUFWpXHowzKjh1F9vYqq81K8ethpip/CZDWLD9v8LiPp/nzbsf7ck9G0v8dLqgTJiYV2Oj
msBAQ6WJO8jaSZz9eHA1OUwljBLcSOEj7V65r34kT4qumozoJaN+xyTsWGc+VqrZma8HDyjoV9xW
nby94xG2LQPQ6B0+JdpWh/zfgbE2vGuJu8OJhHurUfrV4PFmO1DintiYcQZqYM3efHsfw0I6YqFu
p/ujeaiYJWxiOhYtF0uq7mdgzAy+iub2ERaIYXQS5r9ncx92TEy6cQpCgm3fOtTtphtD07ke6xGr
BBIvHOeMW1grRisnNAnytbtdHjS9sTu0bOf4LiNPpRa5IAIBpKaw6AshMW+KEUW0rsfsgOR5KWqY
42natJQ/y6mARECRJm6ysIy9PhPEYUIHi1DlGO+aoYPt03F613j25RN120GY8cjyA5mqo0Sf8uYX
sOGA+PDF7vyAjx87USRQndKNI27Pe6fm4WFHWFVbgiq904HisZDMfLA7H+WVN9stWr+JzdqmSRAQ
n4VXsHF612mRh3urH+y1IObzdy5MTBkAlaidz3Rzvwij0lh0EhxsuPGMIj+mPut7Y9gGAZC9JRBk
JUMVqKVrbBHJA7oXZIgPCPXyXauVm6fgW/xf15oRl3IalR1uE5dr3dGXc+71sImEvzLwiBt6epBL
+4YMi/4bGN5H89uFN1WLxSlbkIx0Vk2Nf5JMcNkFOKXpNSq6xKBQf7SJPU9yoN7nOvA/9VJoht4G
PLx1y2STXApRJ4DB3LPXy+EyMYLttlQp6hOON107W8UaZJO1a/R8gJPECzSQkUBpPno/gQRXo1/s
eb0ZbV1NGqqGc15Q8z9OSbnrQXtJbQDO5T9E39DZBr91gaOpAduKlzkpqVoM2XMhL5QxIHC6CV2W
u1pjSA3bWUjc7TGcabHgc+ZFoERKIG+0hsuO+4RhAtbWVUKsSaXR8+gKGGpG0JrkrbzJM90poBdY
EcQFx1rIH/dSvz5I22KjkmBQMFFYpaqkdbPa2UiSP+OcS/4wShCIXmMsxsGS7vkv86oDv/mDtOfE
xp3R3WeZVilCyOeHXGt1WWv64C1KOmEAV6BPz3PVy0Nvw1NWS/v8gm4vxzsf/ONDBbhCdnq/aORw
qeRo3wZgPRm5+wQTLDdwSXUWxYGqf2EyPoNM77YvuBrnpGoq6p+1JqtoJGJN0Tz8gzwWOqmp1vJO
l/Gxs/0X52vv1UBzVpeYFt7JrMLQmpassZ/Fq/MSEbIoEuk3/9GXptXMsVwTEreVZKnyjh+u1jD8
BG7LxgHleSwBHUmAvr5zft6zfFYLsH7JjUjYMFIwL/mbPNeZSm0rWntwh9yUIRdPRFAtx348owjO
Gl/9UAPt7GPHUFoUVqmocJqD/NjnZrQAKTre/lZItrt4uu+xCBtBmJHAmu1A+9JAq221JQDKPCjR
FoMvQEUcH26VQBqEI/0Wp4wiGOI4QP1Pc6i4KsuuWKDUAlDvEl4NKAspRUXyJLvSWiLW5KY/hRzV
DR/XLxQ3M50zkRDJnhuAZFZQ83lIONS9bz711Iktra9k/Go+nkcyrtbl6/v2qadfNPr5sGRPEuuS
K1LoQawfjHpZVqdmHpqLklzvMrlNSiwuyXIH7umoe4lnUxfUtlax5ML8tgXHVjO7ktpyzS+SkymY
Vtt50UmoR2UkvSZKTNojNvrkN8TQx1ObrfUcanVy813mEIFXAMFPZxO7rWZg3ZhgmYY9TF98zWRe
CSx4c9i79p31KuuNDhn31Ds7ZUyYK6TEFn8TwHoEmB55nj9n1NLDz1Ka7yia7EMG03qflVeQOof9
6dBaB4fkDNv5C+1Cdm2PtE+f+Yd6Jj7PHDoCyc+Qjup1JXp58r1H72J+NaZOx88zvl02SWo818kN
K5HKPZo0bmX8deWzoclmY2EHlZXjlrrhKK6sLLhZU2xP4XCr/wTe63C0sHoJ6jehQXRIXtEwoJ+9
1MpKeBjVk8exFSq5HfKEiNrNPQhtWlH8YFCXIvIGYfxl0yXwDHkvvMptv4cEpLvfHnxDZcCOou5e
78UpTtzbrMdAIUzKm/EUGdFn0OdBTdPx1z+lbmv9KgjdP8joBToM3pyacvNA8Q/t43UXH2LRug7Q
yOHy4OLuDD/yJN0L+eK2m9pq1pz2or3KoM1Avbnbeav1q42nOQKhXKJ1WN3Wu74idc55O0tv0AVL
EA3eJXwXO/y3nXcBt+LkXLwFvr2XMIVPE+Z7in6VjoKOq9wDIykduU3LdIwOWDLjl2rA5FNi2aHp
7cjPseJa+XfgSUKwegAeMC78ZZiik/CuUp1KE7sJETWmpnS2wshbXQHArll3bMKl1xsKx3IXHQgc
SU1WkR8k/j16Yl9BdPrHmu1NiWJA84anFcj5G9LcSZJcmx3v5dOyc+4/lkrmYRdwAMb1nTo0bR/p
Oh1xaILSJ18kECNwU/+5G1uhuEyLLLoy4ZKN5c3vqSb/YhPHCp66cnAJ8SCYjraCpw84oIV7LQG7
z0hsQynykJdoBTX9VgJRQwp9kVFLc9pNWX06VM3sSdDcb1s5iCwivuNJCfZDr03RlCx7pSYtn+Ha
Z5/7tJEqSoeEFDjLYsE4riVD8+SHCiEtEcnQV/AiUgzJ7a24e/77mUNaQ4GMjEgD0C+cFEh4EW1h
ra7jh64Z4plkZLimoGqnCSI8ibIZ45CmZng+4aHkC73iquwZ5MqfDOgw5y6PWmvV7QXWxnzjNCuK
GDGohvAzZXAF4FMSDw02puBu1uq2xQdwHxojFDJ3KFdX8pie9TqUFZrH1kdXag6b/lOU1vVIE6M9
uFIV24bFWPd2ac9fCrGm22ua210+NPszrOjTmH6DcwCy4ZrR4zlkj2G5VN1k9oF8ayhJKsEmZYMz
FNdw7kCsrJWHW3afysODuYpNkRQiXi7YiuyTX/FyBqgZVSB2ZnzDMgUKyOcoqTcc78xWjRoxPYeg
WVDywpgdfvkjCm6xFlmFjCA5QEMvxzi66TbzptRcAr50gQws9jIlmdoL5kFr+J4gn6Ijhr1XtyD+
obcpZTdUAibbPpw/5zD4yPBxPzyqgom1SCgJXG3gpB87E5x4X5VmxavTbkN6FIRh5hB3m12bRMbv
d7KluFV2pFXSjEU9pIDHNrLkGPTBXgdghTAgS9lcZa7fRkrz9mv8eAm05KGJezq0Elb4/tbpOAlH
4mYuZmRbcXCJeb2tvaOUwt38HAi7Xo9PNz+SF9WfnSKDfyr3kFYkzZiVPO+S4qKeUgVvjELKyYTs
Bxdpi5bSKjxOI2C9EJ/ooWKr9Y6EXPs/FYrIKDWFWbi8+3AJ6FU3iw1gJPgEZhsKrHjQyuFD30Ut
hxfyIY27arqilevjz2G9VH994bSaCl1xkhZILVHPpOddx+JPJsXfF8w6S9bHZRqxtUxnkevK6LJ5
8N/BpJTb0ucg38b/GncXNhnyrvCZWzVjBdGP5r+4TksljlMRinDE6XGMYZmsr+GjG4loywW0wSMs
hy6QrY8YkaaocNaXFuP/4g7N8X0Pfo4oUecCCvKA1fQvoFFNUqVJTq+0RmZ7DYCQxWQQn0QIId/9
79VvIBCwMQ3KCvBJiRn7rjGQS80OJJGpI6rqgs2ChkSbHwOQPTOey27DLQEH/5dCCbGIE/WTrB66
2LsXZobMCuSysLtvfkb9GmcGGlY8y080WphOyxvYKKo9JOK3A6cYIXV+GXjeIWlsAE3FZrONlJFp
mGBegT0gGI5dY5+NwDBxIpnumaBbygB19Rf9DA1VCxSYsB4hh2BU6yO8k1hdhR1EjV6u78EujZHS
peu815EPd9qekMBjGMjBFOzFwrQPiptaFBFiIkOQTob/oVdVoZEjnKspObt+1IANmjMWKCz9Q0Xa
LA0Q/IOmYIJi1cqjkGnbWP8F7KyNPoeB1zQ+hn+jt9D/7QlM08AGF1UaM7sZMzvj66OhmLvIE9D3
7yjdgQWqGoJR8nBDUecWPuXpxAnG2ZUBLg506rGbHEYGZmdb4xNhT+0Q+A1eL6Sgt6de8PTMuA15
MkYbmCua8jKe7gTJgX6hUacD54P/ZKgR/MxgDnUUOziKAxcukVHLxSjjUf6ojVbf/o1RiUkv9Wvh
pO/mZL828Stp+C3JLLtXKJz1MabV88Lh3IxoxL8eM+BDvSIELh91xtjtVS30qH4ut6PjamWANSrz
S7VR72agDpXXi0bdMqGL0cDAh9lbExh2/AJsqOI+09faGt0vK/wn1cYZgFoFOfuZjb6DU7jrwQME
61lrzh1fjUdIZELz7IItVxQ2PExCRBDmX/olqxvR9J2sj4Jb4xxaM+QZzlDNM7CKFXZjjmQjzf74
qPDhtKpIdFMWWqUtNDkSsizs/i6C0j92jPWJsoeLS0Vo6Wpye3c+IJMLXMPwJ3osIzm2RbI8BpF7
vce/vGcbIgH3lsBup5GUFSwAmKSDa3ol+NaDWXg6YIGt2pa00LTrT83uUkBnoHNE9ilHmADkbshz
irHW6TncUVU0YhpvWg9lOgztOXE+yQiVkmvw2FEZAYfkU6GshXeDH9VoNErsu0Pz4S5ULB5LnH06
saiUDRtHOEtgFpYSgpoYIBjFAy6mm7fI3FHyD0wxS3/MT9qjfutqKA6FHRtUEBJ47kH7uHAIHgQ9
SC+zplwVx0kzSuVWG3sDN2VoCi8dkvDLj+60k+9jrT0ulO3/e1dsGeQkiOQd0U0yMX2lNi0Gto2K
OWhnB6SZ8q2VPetT3z5Jw872GmkXYlE+DZjWM6fsryHPlmeOMaKjmw/d830vMUsRxKCnzQOgycVy
yuGJ1SHlhxxoqVdnRYWahodOEqGUon0FzOajaRn0DwUcgAKQMoxJloFPS+JSa/9XJm4zksvO9u8u
wzEpAsYAyPM7ysrnVO7G7o8CpOSFGFWaFbrgx4EiCl7wvnEu4dhYAUdcZtcDX/TqbkOkB122taps
HgnemKjcgLzIqea9voYZNswVq062GGgj4PNU2lsPmiXSSdtKVQeI3sGGAfUkLScMtnAP7cJxYzJ9
Xa2AX6MzXG8YpFDLrof/Y2JgokY45U4z52kojMDZL7mYyPAOQrVi0MHAOe/dy4Sr8rgPtCUs1AIr
YhzuUolasuqqpBmTsOL0ntorSaedxdjXVZoxc7C6Hr2rKEI9zNpdfHDoq+wEa308zo8TTHc2uYxW
NAA/hQq8UKmUFLwOqVYGkPzrjGaQ01PAZrNbSGZlN0khwGZAFxlRczt1vx66NGKRHR7Vl1lwqJC+
nUUO0sPDuKLTpsErdzbrjUc+s6YIiM4SB7a+qivYhhalQmyhjYqpuveXI31BNvIZUGenoOCS8hX8
JxveLW7rv5Vh9OjYaQNR85/xsRdFD5Kqfxk5/xo/+wJVbQ+votugKxIBbu2iwTtJAHDZ7e9R2/t2
VctwCUeGyR8oOEdktWU04cfiE6Gw+IjyG9+cWq+mVan1UKi2HVxYJTNIqvE6Gwwq5Jt9DADoEt4k
doCb4U39Cw0rb+EPZGSaDl7FFOTZomlwjozGkm6Wq8MYkSyba9aH0C4i62/e3X0XAsoucyXM9vZD
qz5c1uIZOKhRmRiXG1DpaUlylFADBzlwxf4wRDIdqwuRbZ+e+travz7xzltRZJrL864phhwdhLVL
Uo3zoIVcJEKhwJI5sTI56pGAH/Z2/9HGHEQEB7VubE3+AKFzwCX9pgYoXSdme7w+yfJyx6ANcwYl
qVyw5KT37UfNso1ib3iuZR4Moh7xu/b/uIIE7x2ts3NKOqu1pSxhWsncxKSyO/q473bj//leYKob
dahRBX1SkL6IXgPiCvss3NFaSMk0+axfuDy4JAriYcWTL1uXaB7C/oBS3Hf1IECXT8oGqT/UgtB5
oH5bbLfR+YJKxSJ46Bhhc7xPCLpmIPfC8w5umxGnGZ/hXUx/ceVIXBBBSO2iQUe5/kyv+pWCvbni
CNIeoPrAfUtCCPJOdGBDDW1lzCtxpsz9+bvhI5USbdKacmcP9Tf8j5hplctOH3p+qZ9W9gxW2toC
zo04uhZzFR2uwbJJwbccoRB+bOXpJZ+A7lQ5pJ7Dk5W2xsWWgkuFTFh4Gs0Mh+axdq/KYkyPni2M
he0ntET3TtDHsmEM81VaSm3fvuRAQCEaDpya5ezVM+HtbVn8WEK0tzdzd4vvE5WPfE2XQYLrlECi
vkg9AXS0jBFLfSnqrzwaPZmqUgZeCvpxgJaDDgVh+aBGAWMGc4wXdGku/jo/hY5zF/y1hhNQOR+h
2fbuFshZHvSp83gn94GGYGZRpEf2maLb8tXlqBQqKfwDvVIiI0aAQ0aJYmV0Bjv0N6SXa4gtPHO0
6J8EhKeb2SfUtb3Q2nI1sAbEC1lfAaPU9fTArtM/z+sByKXXMP64PtwE7m6iRxXtPwxFDjP5szeZ
fKXVAqoUuwZQlT3bWjx5aUg5IHl/koe3Uz9pQOxw+YlLWl9RWe9pEff82HlC5k64n1r+erCAuA+W
A+MXKZtokHJ0sW+3EbKSHdpwPksjPkBIy2pWgjn/wPrSwQKS+iR0k/6wqQXiT9t+gSQhE8CLpbPV
y0zDQpex7aQc/boWrxqIN9h6ZRxQYlWxCnmU/wwz4/OF7+EGi+Nyj+ti1wUHqcP/ZrNPF5mepTHv
/Tn99vY0Gd2JWRzDfOqLEKfXVZNBaMZdJUz3gBPs56Y7/CFBklS/gZi1jIkN6pKsW2C4sSVAOb7z
2js21jXRGAmVspFACnD31xsUq++otxnsqgviLmp5p3RF571Z5OtS559cXsWrsnn3O+1ANx/sAy4l
PvCBD92r++On5CzAEOetkn+l9c5z2DMwblg7qDCeDYNsaZ8iWJTVcQyHkpYnvNwjrPtribC9mKXz
xgnVf5qj/F4JOK2HPwfgw1/4t3thnY+r987e9MgKIQp6HVlRIYrfo2C/c/S9a92VwUXrsfJsCMeT
SttD42+Rt5VjJX4VUr7akrtzE4tRbrPGMVvvzcjoKmHQJYhbNj2hh9n1pg5NIWpFGq9tbp5zL9Kp
UwWfdckd8zPH5qEEGxdX7KsidQJgpPFcs/VWsTctr6L/FsFbEk0fZTMeIqZ6SKUQg5WvJ2rgzAeV
yjVO1pJGEjHBDwg3izSq4IflB934pW3vbC1RH4XcOmbekoQDqvKBBA6/KBmfGVagyQmEhBJjVQC3
QIElR4M3witdxAqfopQW8iZ667xWhFcGG4VMNcswRaHI2sU9EmgjsQXoTcn3+ccUhzl3QbodVKgQ
/nzSXYVQ2fE5WDpzjsj5ZR1AV3kfRPE7yQ+L5goT3cUGEXFy2Tv8cBjuXlZIypFQ/kgSmpUOENJr
qglmxAslxVVWmnPm9IARvATh3kgDPcoHN4uCZLdFu0obZtTds3v6muC2y2OPfZO04/Ciy1qF9Zyx
dygaN/mRmOx14RfEFMkScoYECbF/5Fb/8K/txvsPCjFVwbw9j09pkkwYSpJ7oy2KJsRuU67BhJiK
lJiVvlf7KwIGlktUMZfIqFcVRSTuBmDVf+2u64fFE/BnPNrCp+hDtYWDXyb/ATt3NueijB8aaw+6
AfgjNLYjFfZ7WqhkIWkgperPR4UKfz+zCMTI0qJZ81G0RvlQoeBpokcmCORUJMVGwXtDfVzdwNfK
4tBIBglemw3KUMY5oLx2JiK0qSmXhtJobD1GokeXqTtJyrluVb42SjKU7grHD6AcFJTHSvy5eX32
A+niiwXbR+wADU8otrtUuEKRFCzaw2YLRnbo18tku5QDf0Of4bCJgKcD6YYwPxrYZl6s9infS31J
HUSEOhi5YoI+YGBry16NobfJPWNg2iBMCsimqcYjDNAPIRy7E2rphGLUWEj6UQgSkJhDFvebm083
G83AmmsBeMtjpUTFNbonx3wJqrrYEaP3v4Hsk/5FdOLU5lOkBxaIixiIPT2e8ajot9u6PHuhO+wQ
gQFvEqnjuo+NMelCqIdR0ENoOD2yYLaQAS+6AtFUrAOabqKjzbFd30Uvs2Z5NMaQMHArE0morGct
PUmnlPVWhG6Kw3wxIaw7rLYCRAQmbYCHGAP4FasxNSUgg4kC7ioz5avcMgLWvuI3ph52ahA0r9aT
AOgKDIyAuldgO6wie+urVNqisBAHn8tiA0JrQaJCDXR0HYx//Udn6CbuWBQF2mwrJ4oiI2p+zEXu
hgTJyYy4eXlwhgNqtbxcXMM3iVsh/9ULgsHxFLsmRXoQGYF3Y08Zq9vLMZuJydJiI+PgSxVGM4OT
qn9YlYSQYGxNbq7c3uHFtb5LzFKBnrjxwQ5BREr1PIG5fxk+/4oDb1iLhU1TZFFod3VAQwvVH9qt
bASpudW/57onK4lPA636hF2yOlNYBPBHMr2VBZFKPjA8uN2i1iWMU9Id3b9qntMk8fmC5H5PIGjW
TG2TTN8Gk7pZDCTCrwtQHXB7iQn4WOqtwXroYlTbGN6Lb0fuKCRS9dSAmDhSdNkS2k7ElEbyMpF6
V/Ku19dGNI45GPHAhHZovFPYsdL3nyTNf0nIDMB6S525C+OGeeHrSxX7uDR7wLNqpPfNmfn8i9ex
Wzk7uU0N40UbywlrxTGzwErYrYQLvNPhHxFQEBwiYToZ0C5ehNvFokD4OT+E17VNFGWeTRVRdUWl
JC3C+ZJsBXgrg4GCdDKUaEpWycyDk0OZHA1C4SIZJCna7hS6nPoxS+ovCfttHsj3GNKhuSCoFaUC
fAK6L2Q7iHH+z8QB3nBGaQQz6Actw+/9T1pi+dvq37pGV6yOy391Y2L3OI9YPYD+euqK2Z7r+SvS
BKXo3EJ3PwHkmjiArqLUN7oo+AAmcE3efyQhxZ7f07TXQ+b484R7guK29MsYdCpoM79gHHVL9+Se
9dfY8WaNm2q9LBxxhVA3oZR/FPjKRPAjNTWyNffpuaGkJQn0Rj19zm5ZxSZAnSxeBVsoI25GsKxj
x1CAR5jfYQFDt/ipTNMwkkAqXllJhwgrX5KrAr0ROwSnBHiojv0OIRDWjQ5DxfnT4PMQi1AZ7Mej
fVipLcqd5zoiUDkceoVPDr3aaubKuhljNaH/9uaCeke7L3ZGJk82VfW4PGQBZZ+/PoCEktiDj5Zo
rkuHSaMZMSljR8VUOwRTcU+plgjZu6ZkoYOn9GhWa6PvcXybLQ3QKF2PEQOZphJPtIiG4V1h20fo
alk6fQEovJ2UElhdyfG3c9YoyUnJiEGeKR8CrORJsmtHg+AsBDsZ1Yp4E6nbRDIeSzAADEqJH0lI
R8IwMZo712qB5X4pPN9JTCQWpU8S76cIO7VqGLQd/pgfVcDT4zGloapxGkI4CmC4H4XgfF/INXLi
5p9z7xocieULWV+usDQq1Pj/ugygf1Kiu/OnCMfDWLRjbgAdelfhn9tWphxozIaf4x99af5E1OC1
jRnj2rgcLbNO1Bgz5JtBp16ZicljUV63myjWrsASmcsU8V3/GsFx2UlleR6Le11WJUjsaD6qDPt+
HTwC/lt2FuTIqXuzVXP3O5g+QELEvLqUA3mB4NWki+7SXzu7SCoLzSKbT0NrGRQHg5FNRdUlIkJ4
cY2c+3Hv9+53SK0kQaTGS3xjF0HI02G+njgbbBtKLXziGrjilObkOrDVnQTm1ilOFlD8VTcZuBSp
BaNr+/xJ+XIC28QWJdxlb/h8HYFYlYHFsJ+7aj9QR2zgBwnIrNwtSVeaThE9kmfeJCys7IS6Avjc
epALqRSy+nut2rXPb6/rBNNuRxt6k7mqGC+fDy9eE5Vo0OcaBujYESVChCN/eY7W0RWTVJ8Hteh2
mmEOUXqqrruPikzV3BLmBnMMa+owcKNNboU6oluY608f5CSemfW4EXlah8m9DJipxXV8nxSSkTMw
2csz9HhAAyUsYNWCLiRC1o1Jqh2PXvDESUlkGDQdWgClLR2OgsLe2QmHgUkmxqPwUY3TrqLAuxiV
UCA4aapvMCnuiPe4N+QJyVkgmV0z5VGs/yFhXBDbApIy7sBPx1bI1xQe29k4edPtr3JW5NCh0AFR
GSdV7dXRxvPu/t0KVT86nUmLLIZjufysdaSRMz7QEzpDz3kJBKLYLc1A3zIixL1EzT37tqoQTCC2
qy87E4gCqy3u9GSapSbU87HLiuDXo0nvi8HFzx0cJOSe2+0iG99k2ETXV+fAYhEm/c2Tzx+snr3u
63eo65JItKuAG1Qm/ZuCzkK5F8z5juam/jfW7wgE9+kdaxusXpmKP4eI1WONLvA9fUyBN3jmrc7G
n7Q3K6TY9gKLv+qjehTwG4/VX8yGpszz//lE/mN4tjoxZtZ3YM4pcLRnMmJy6nXaOiyCHl1at5xi
pB6n6moVJhY2p2WaavkA/OSut96vubj3EssEdjHJU3UTjzRcN1napiI3TbKNNmkIc3SIhK8q836j
+cORF6TI8dxujwcgfDg4wapfWeq37PbY6itWgT6Ibt0cSd713l2d6+FkGgS5z/uglpu71N8ccCZV
GUJQBgpCJqlYVwh+BrmowSUbYQAB2547aHs8OTpcNK42xDRJcrJ4cFo/a/SkPZPp6P4vl058oL/F
xmyJ1xnEru+COuC+vOlLe817BWJDEa3Zgc6ZruOPFUvICqTQMSwnOh1u6oCtScTuo3ATnBFQU+p9
xZaprZxI+7KXb4PpO0TjS7iT9Gh2A/Rvkbz3S2UyretcCFKUSLsuEGxvQd9W5f/UgfRWkhcTRyfb
d8PHSxmdW/QEHsm/lakjRKOCMWosWFKZNuIqOymWKy0Yec/eHZRhXdmQkg7BTlUqc45/6odX3omv
gH4w2/qXF3S/Ogy0Xe4VugsdiIr1cBk7cX/pDBihPPJSeINU9RuV4VdPvh+oSZP6MiUkoLYN8qDg
L9PkAxqDTePW9an+137TcJ/QCeTxlGBokmAncfW7pJPU08tWUUWq6cuiJR9c67O14B9DWlGlkh01
bInfUqIgtc7Hfqc865FecIEuIfq2KLjLL2rnJCpYv0MnUM9LZMU/goWLobDURrn3iYTDIxbQi5AJ
Z3Y7WHmfCrACI5UgNSjS6IDyzBrJymm50IkVg0JCi2m69Yp1reeJ49LzWCHyf99TO7jGcVeAAWpW
3OLsMyMIeDDGAP1ztmMY0wmwhcmMDFvV88eDdiRtI4hP89FWvF/yZDPsEm1htEROtKC69/mc7k+i
sJrRInuBuSm4grzlvYtJ6Uqv3uBY8oQxfCShSnAZkEL4B8Jeypj3YdxM2sJJ7uv7BqG1tRBwbEuO
44bJ62vbYjNor8xzeWqtS/OkO56ViSTkwfYCLan6IOPW/vl824bAS/NLL9siXuGiLKt4uKYN10m9
yiYKsfBdLsijEwVjcIfyqT1e+cZJvXzCgJJD3Ywvv6mmdGpeONj+t/xzjmU5B5QwS08sUAU9nVRM
GpqQ8Wu+xma7M4v/0k1Z22jI1gwnGCwFvuwQCUo6uIAQBMiqGsoNQo8yeMHVSu/7LlkiAyDUHwWy
cVXxJvWprWF93dnq0QPdQ1GUmv3+e1RAnC+84ylcrJK9a0kATa55AyEhFORU8+++Npuph/LIZ1ji
D26rILyt5BfDzQUa/FcooCsObPRZILyqsUg7bToED0fnFX1Ck05Xy+FpbHm7PZ2VtTA+iB6zWk8q
4jTBk8K/CsRNiPsLa6lx07v8SzL6aVaQ5g6FarCM4aY/isi9fjh/dnKGQlSTNvcNZhtPvTPRU5l4
lNJZ4FV/qs0AXySjw4TBcf3G81nmTWc1L7LAy3c35AakA6TyRX+yw86Ki+PKcpXTReuKzSXhaPUX
auq2Xb64JEK0lqS5iCsQd1qM90MoDskJOoWUCr4o+NQwXHuXvc1PwvDmZEeQSai8qyhq4xoAA5Uy
iXEf8zOmjPQP/73yAK87pCCBoKBlZMPhUgqR/61x3VvokUdkVnYqemWuMQm9e6IjUqUH9DlBBtXA
8bpuDVtDHi71R4Lrr8YGXOXHPIrLM24ubk8K28rcQhM3Rq4L0x7OIsME2rz+Rh8xkO+SBOiZ4mSb
39xpNOhfpCAvKtFdWkKg2RAt6nEB1ACOCBsop2pXiXiajX334Pwjt6JAovFu4Ux2bpXuy3Er/aRN
DHH8oPGL12ru/RA4VUbYG5/m+0lrNaU3ZUH+Yjg6p9mqobvq1o9eMm6vYMhSADQATktjSgWtX6pD
wophxTT6MA5N7H/TEI33Lh83NIRjvg6C2G9Q3n5uHZKykNUYmA/6uGbRxil1uLt6E5PqvS2/ZDRq
IzBa1lYmiyDIy94dpHKri/qtZ4+LtnidRGCMrcE+Clwy+UiSmuaN7TfUOlPmrqbkhSMdsH41ocM/
cnwyx5OP+EgN7kWTPf4A2Ef5FaAc1W9dGf1S8Z0zXpoTYeWBlKQVBlE2MGNXXV5KxXJZi9po/wZC
5nshm47eNer6cdM4gesOgcJNB2N9XAAjRTTxUGV1fMqsHQGeahBf/ff3GE7k7zn8g+kLSkKKxvC2
+cv39Phm4VCRH2cM2Q+17MNooC8BEB+lYRvB/MKwXcFRNHHM1edsrPoVak2wfObuC95fwnF/H3Kq
P4kqbEYcG1tG9JNRZR6w0CMDzV2Pmxcur6SsibF0xd3qb6Qj6YrYsackAQpwv7S5k8eFLLm2MKfv
Cgx66cao2SJa2AJpvWOuTUHYJVjCjyvf4V4MFqshHXIcIj9HZ6+O4Zbbq5Y1bBDlRqK1cVtb6KaE
wlt3QJWDushWdrpJoMrSg3FzrdULc6YQXYvPDujw+W3l3JqECa7dOCltEhLLAjvJ6Fgi4O05pCtt
NWYfPjQhjF+TXN6DdQoGqWL98oG2F4NpOl4H459BS+EIb36fQyXE3iipCIW+Im+62NCeGhBQqSeq
wusc7veKAavDRDFqgkSW+ZvufMjEhXPjUWfLSHh6pwoBdG7A8AYG8BxfXn/BjdcnbqEuuG4ia51i
ShRAiTaS7J8sNcNCOiykUFwk4lAWWVGqqaT9BnUl1UgOIopcponUfsu2cDU9Fq1mgUufbIsrWeWZ
k0Qu51d8Ev4eIjmE2DBOKOBbIyzCwjtHIn2KQr2B9oK9O1A1PTQRuVWa9X6lJNt9xr4rHrkY3ING
eW8tZj6t+6BN2EnJ4YtH7eO1VbC64gOTxzjht0PBXdaTtHrmov0JAIkpRV6KoqjLse/MTup5+OT0
PXr2Coy/FnDboCJ7CkbXRdPYYijTcKK+HirLLMB7XbvNlx1HXxlQCe6Xi8wAKFEcoDUv09g0iUNf
WuzL5ionZ55Ny1kQUN3/3GqwXs59EEjhzn7A7xyZHDNqDYQH8cOnB9REMy+6VXW7nNC0xl2bkFCC
Kpg0KMWhyHC4jiknbrcalZKSgMSDVrG0nqOdTX+N6kSbtXom3rUBNbLKSGlDZXqSl6teuyzr5g7v
VtPf6NdX4JfMDnVCRLjfch22+H8gxUT99WdD1OAr74coC6iiGpgiTAD8GR3q/q7yOlQ/Kj48epCF
BflJZNOHi/KYq9DSn8h5cpy5Oqt0EdZg0PoCVSoVa/mnfkLnkUFg5P0Txhl6SrC0aj/VkvoIMNWg
AA679+innMRo6WjwvS6inCXczHkkBXR+b243QkJU0H4lI3r3WvNeDomdoE8Tnykt5Fo2iguby9mp
m+1L9Ud0YOINepWJJB6K4vO7Uov4Bh1joHcNX9t5aLhaj0L8odZA3NtU27tKKXqULq5YPlXCXIL+
CR+tYtIFvIRwEgKjtnF3i9sdGZHI+VwBfPXgRA8X7sulJzEganNpvVeHI6cVLB/R7UGgGkM9xX1t
AH0psgDW0a1DBOjAJC8JEkgKoTNl7yEnS+/RraF8by6WJofcDXHPX3ggF21vcZIGlo9WpulrrwlI
bhkH4ELzr+Ql5TiAFM8wEC/CN2TGBVWC0GeCGhL04kM0fV5g3qA+HmgMJxg7Pa5KXdPFVmfqym2Q
BAFu3cJfj778XW9VnyS1VvYpNEuytekMfU/7yeem21QgvdIXdUg7tsC6OAjnBrbRz0btS9EfSkkq
CfZ4ZQ40TDgnBq3FqlDOKhXVk0NjTIDSWdSAP5F62LKU3Vnl+hnZfSzGSoLi39uTxxRqPs+dVbZs
iOTJPMH7VUMEnj2nwvpgJKeUWxfg+YG/5p5/yzAFPtt5282v1RULKjE+8FwiupR+4QJ16CfRP2qf
E7WqYMj7sy97HkP6MtAFjS/iuHPGc/OsoMuyg6xcHe4ipAIGGVnDBxrw/grU8cotVC9yp3YotIDt
0tqVhem3zxRoJp+9BYMkUFJF8QFL+3kxW9xSvcmSCeu3RVzi4juJkgGOicB0g6FwiOljirHC9JBh
9ojQ+ETQ0KvzHOfeW5FCkv363IyHtChaKZKRU8Y5j3NJnjE/3M7Thbx2ok56MLiGLJK0faN/HbMF
63Gur2X89ET/LjMeyJaOvqCHBIB/GDLKFd0t5ymhs3I6xohApJvjsQJwC3OHQDPXzTmaNzIwToF7
4tcqoQ/sfDNWKAjIrtR8E45zIHFPz7Xbn3qjAkAgc5TyAGVl58WSP42KaFZQ6a7+ffuPhOYRi8mV
kOtuwQWIADRgBiF4vViVgXB+BvGDctCIdCwpa9CvCKMB3616UvfBV7pWOYviP/kAo2iE+jkfDJPB
m41QLGbIinPjZ89huMAZ5Vgu5QV+mawSEHjRZSah3brKN4gK0UoaBz11U+PBwbswFQ/FJNKXaSO2
DbaHJtE49hSIoaPV4N5PnouAFmq5XVBL0EeGNsD2T4pU1udOgbxsbT+yFWVaeWzp+5ZSczWyaAoB
+E/qAsqRG3rW2Xpb61Ri1HHbOIN7KWs7GU8PmFrNux64IfYto7Yln85393OPGEE1GmvWswq/Q82S
mJIE63hXMuuWxRHCwIa/IWYY2vBqK0paY0Kd4byYVI+KzX/gkEqv7ta9k3GzEjAotVmVysQl6g5E
nZRXLu8Uc9GKNvyfDQHwNaZ0/3HNYTmx5jaO9LKHekvjpOEuSunsv6nMaMppprTZnA3zRuyE7Ji2
UzIOVcXrXiUXWKQM7/wm1W7no9nfdZRpjs8dnDacFiShlpcKBJg+1Pg7ufH/fQbfjUS21BU0cQp6
489dsp3V9mE6/jlerG3fzylSNoOVS5yUJPB+VnJ67dkTnPWEtSGh0AdAL6NJ3f7yp0KOs5i6pbcA
QvUFaAePwuQbG/h9P+OweIg1+kHYZ2cD8bUeyL0AK2G0cfjmKQVVceWJJkinPFxx4QiPlA2yZVUl
G5Ckz9VjZ0aJngJtjFTHVcNjpbv1vRwAaRj2bVbzzOtINIIJiNCdyeWOSqVcj9343E0weqItb3UD
3DTRYOeXeq/8tiKnMGbYmUFmvStnT+x76SFtz0FJO8+BkYp5HKdk52qmoKrJ+YqfiISn5amXinez
CP6orG4kMQo1Q0BXhJ/2hW9MwJMn3yfUPz7qyoAATiYiVvYs+8yuij8DdyVgjhVsrLjRewFNVRAM
YS0gcpPUt1c5/xiYMnIe8sZb7UsDfzDIDyTy/bAqjibM+rHkXB3vaJPHiKbFSEm8761SRWEb512h
sfAj8VipVoaSZCOBjugT2qSXwiRrYXpoYN4LkblO8Duk9B79/vs4prdc4rK3mJlaNDj0EZwgP6x3
4Wid8JrPWQKSh+M6zeowIAflXwa1mxH+gITwemRszqLvrmjoEICJxS3vMikT3be6uOrY5loahXGB
LOicl/OOuKNKMT++j10bC2wiYTSktZsnJCQdCDKmGY8p4zFV0FShuFOlLrWyV9NsC/sIy1HiA3o9
vSXdeYzbzmBQO4WhcMha3C/vdpgEnmDgbg/qcMe+8ltSS97OoaTzZjhVqQoYB9JbEwiFOP/gPC0v
O5WWcNm43F3YZFUYyN84y+KQ1bES8zx/lXHGQ4oXE1ps6VDSuUcQ+D94CpL/4lbuGPT/dI1ruFWS
dPbYz6zY89J9o18+A+JIqSQG2jwl+Fxp0yY2dG7oRyFZRlC1hM7Rvda04vWBTbV2/XMp3HKiliSP
PlA8Z8dNjbDgciMuJX5joGzekHM0j0DxWjI8e+DeLHkONmMDlnp3OKCO9OR4hwOfhGOKlFPOUtUv
PwwiM/y4byzhKMfFvtHjE+DgJ+R9kfsRWvcQMVwPlF9d0bPHIoB3FcFug7wNJdUKJqb9v3/iCCva
xDBtIEg6QwDNrKk/7PsO0PYfntX73d5571QXZq2X/3Orf+qQVNt/JoXhjFGtRbNNd3Ap4cTbsWR6
hvfbnRe0qY0yTNqEPXmIfs+gd+qODrj3zjukVkztzMRJvbguvV6oby8hZZrJ3LUd7rdTiPI3Fkra
28l8iIzHJ+sMyop9e7Y4q7MRwVtauOXihsl0y3F/AJ+Hg8f63OYWu30rfhGJL4icqppAiZdnfqvh
pBvjnl+zBX458/k+6LINbjPHSygi+pm26c+RmyCqhljQI29g5LVRJXsrt7UEwZqOSQkWjiww6SII
VwUNPK/ocjBY+DVga1/liOFThgEfgabsyzU+c6x3WmzS8urqF7GgjfrHCUTTloCxumJQ4FJOCreI
dyFgIlTXac63PQa36r2QfeX2NDW1tDQL0RfyFMFA5tgfjZSluu7pZhuqdR3QtTyi/sC+jAuA2iWP
uK+zGer+652LDmH9PkGsb94HDxJPVXW+qxxE2zPByQ0d1P/RujXlClDrEBfQo6wWNWomg81TC6RB
laBJ7GTuLdR2L6UfUrd8li8DNuaGa0UYX06nxdRpXO0EIK7z+ax1IQ2aWcEusvjkVlt6AZK2I6gy
GKxPofZCe75KVhQqx2y6Y9aNZPX8mGEb+EqKUr7PM09Xg1Z6i+N8IQOsQoLvrXJuQadk4/sV0+RV
HrlrLgr7ugQ2Hek+/NR6yiDncEDjbAOTVBMp0aEcVT2sZPRnmOSoibRIWOItxjALeihM1on8aG+N
vM9//vBBxZrQaDkBjw7yhD7AdqYjrZq9ffbislcqR6eQ+3yf3mbeef2CKiC8YKQEn6cZzKleeHLb
KlZzoKGhX8cUq7U/j4OFTRmIEzbx43gRnanpoE4lxjSAewkr8VdOoO90UuaScGWRRhy2k6hQg/J9
GJlnXtWfpOJrABTWYjBpGbFWfKm/CYhoVZjhzjuMXX/38ygb3jRdoVsvzLt/fU5LF6INMe4rbTGS
MT2RKEUHx5+3Mif/hUPReriTIJcvs4LwdcqET4WNt+/WbbxU84zl9D/9y6gQJj3DdzY0RP1WM6hY
4BkXYllsv0BE76AcZlvN6RQ1S1dySaBo3QWOBlD60UkbthGHCrEbP5+BKC0JZoiKjYAlWUgD9cJF
HHT2UY3QHD600thBMd0VAcmrjQ7+lqYGFV9Ff6jzdGxVotB1tcfJc8fobj586Ggngywc0MDLTxFY
VTjRhWj4x2SANqEWOia3WpaWulQBREDj1J/qP5QWOmcv5/wokydAoG5ga8atfvRKwqkXrPkfg9uy
2mtJFqH14gzMiYZiPEd7GGIbI8xSU8eU+/VSkUzipgt6JinadKO5MmtjdfbY3hTcwn36uAcfMSeh
p/4bDW/PYpNTrkfjr9hlAVSJube/db12Mx1+HV7IhaRd6p/T32EgfsvhyWRhrV/zwuFy8OPaNWYk
xnrO5EtBFgu5rmORl54wlDWAZX3Ym+8olpqV7eyD+TvYknBSQyRZEhnuwjN5TQ8V2U/56pRcn3rD
V5TpGOfDZtWUfJjKRM5e3viwFytsNRpQ3bHgwk5vJV6ZnhyL/5ffxBE05c2XYYm3DOswC14cIqHz
ynZ0znurfQgdtMLKisQf1p1eyUBmR8+NTNFkRacxJd/acZrnnKyRxzD7HiUhLWFBd3nHNl3BVovy
bsKgKo4UGPWul8o/Q9wLQw8KuqbJwY2ufnc1JDLjHNBh5g9YXRjQmhqsHvWk4YrgtXcj0eEGUdeQ
2H6vaWiqjyNZ4dTtaJtv6pxIpSAtZcxYb2RZVCWxQK2I/HOognmfAiWcjZK6FW6KcBPpLpsB9Kn+
ysgF9oWetBbZpsezDLTlbUQ/GQHLLnOUMs213gB5bAmjhfgzVHtLDXRDUUU8vL4aF2kg04oaGebx
1/K5XCOLOkoneYDSY4BxHdDEl+ctFz5IeKvz2wHqhRZrSHs+Lt3FGF0P7rkZkvScRTrgnbefiqzC
XPiOfmLEvM2UWSU1Ao4yjFYm/44VL+lNj6q/ZEItGtH3NW6/Hz3WFh21ZxQS+qKurB2pUhYI6bcA
H52/Yt6NuPxW719gWXOY5Us4VW392CHvMikbUF2uUIMnbZGSwwJAu510DBrmVmsL10nVdREUxp45
1cNqOPkzG8SVOxsEfK8dGCgInSxohFzea4LCDIH56VmFOUKyJf4KoPaGqQywmirPYwOlAE8DDWn4
0M0ukELc+o1ukmpaIKEP055LinYxbvXLhTqA1g/YFm3F1c1XlFtDrYBgHbRbaXqvKVW2UMOeM+ge
xMP4SDYFdA6D2wudbsNkGyKRmO5Hcb1DFR5szA+yUCb2SKHDcVCdPYzFaRyOsShJO9wge8yHvMiN
yqJidSbNdEyozaAPQ6wRbHBBW089Js/wUvYE+aoQJyXWYjh0fBaFrbCt4NiV2B3GNtutOpnh0vfL
Jw5EoEkX3GabDtf/6B3PeZVy1ccngm02JJG9F78bVXigr0gk5M9mlTUvjTf4kAiJ/NwfyUcjDN6p
nGjXRVJxh0VzCas583nJoxZl6fCY0LvVCnmqjVJPUj4bNfahv8Vz2h84LNWHMRKuyyaVgGo4CC/q
aiRxjZ08rWc0YU3KRpLdwx7US3Vrguhn4ohpO3N0At8UZvnIiLF3fZrty7rD6PBKkqyJQq8t3vZ9
FzuQe5nj5nquRPOKOThdRMe7sjqrqw7ZAAgOQMOOdAaujxLy/XqrrtUB7fMEUtTeUkDriwiVxmcR
bc9y3U+j3/16tnfUc0YYaYBD4ARH7pUj0gHEfsa46uC/i4rKqLxy79nl7ItVfhKafLBae1v4UgmG
9dG8yLL2VXdAfXLS6HXFTmsI4nHcMMomMqSjmyxiVcuCXhevH1BZxYz+mGw08gtmw3mukYL52cSM
inH3SudvdFeJ8wmI/U6dKeIiS4A96ll9E3QGxUNJy/PQObbYvG6amnwti+MBFmB/qIBfMapWc0oj
yWlV3zrMMOnA/litmy74E0/6Tdpaaq4RXUxmvQ5ewnpwl9IPMkrW4zlnpSAjvZWeVcvhFb1xXsDj
9o3IbDYR5jI65QgMovHtG7tY0uUidNIAxZnyeJhQT5l/tg/L4nQA97Fz/DdTB4F9wXzPnZ+DcsKe
GDXp4LTCl/S6xHI4tl0YN3Gf4PpluBIwQMjVnD6Kgz+fYCdKfk2fY3+MEqujFzXeYMNdOCFrIKie
q641slE50ZlqrOwEbiuie1Q7G1YdUfAWVSv+fSlB9nppoQQMgzm5ghNA6REsVKu5z1+XUI3dOTUp
X7TJyZe3bNWudSZtSLtxN+QvdrZnn1+fI+OMWt/PYCbMTz7JElDmEihrkgvhokIWSObFOKZjd7e4
QbGE02ZWnlZxloVxUq3qtWZO9TKl/2cgLmQp8MDwu3nv+mfuH+3vhYAvrW7DzQonLmIycZGFA8yD
rDFsuT4BCHONCS0zrCAlHrzsUNubwiI7X/52pkx58QwCxngsbeqVbEe1e4xtGFliAmcJ99P4GROu
UjzOiJIRZtXAcgTrvX1WC6fQ6Fb5xEvtGFrInmyUnzR6Ep6kYVNXdGsp/Fweu3/GR7OhYO5trYF9
gJDuumVSbbw1rDF6dF0TslLWgHoYvvix/O87gdQ7MEj9fMTB5PP78XCxy9GRorQdo3EKnbIWA/pI
V2kjd/FrySDWzK8cf0nmGKWoBpoZYX9vIo2XVTtVDYrN1HKpVok8FRyks/LoMdRKcwFaL5qPw5if
aznR990BSIsNEO1bpis5gXzrYhqyA6U2/Tr67lxk8XhZNcJ3L4zEQc19UXvao5XlPEKZtA4uqt9m
3ijOWb+6stW4W7wiFGdg3sVYhLIUit0YUadQV0ZqfI2zNqmxDxDas/nqI7CogIJPltPZ0CDboHJW
GjE/z/ZGATVpMKymu3ycROCv05Lu3H3hN8g2v37npTYhNoHDUh15LBH7TCn3ZI8HBoNUxTNCH8H5
4o9i/hsHTJfmHxjX24RBbW22/3F2Zpa0+2LgFc8x/95BEx4QAcXWb7hyIvxgNGgrLTN/Ux23CZ+/
H6kCMxrVLxsPqNB8gCSrtXX0v2oF6cXABM7ghB1Bxp3Ijc5FgVIzePGF+3LWoSrgZTOkKdtlVG9U
pLuPX6eGW1D1vu+2dRolxP75SXLHxkxxOvsXjDWyeGiJ2hmaxdPNDeYmLC0ix4xAuQlcCJCdizTT
y3iJ70M7+450UG+p6gNBEE0mMsQ0F3XYC6wq8nsj7o4nSTxOPjL+IVW15HPErm1YDXpJDeW1l2FX
+Y/ESI3nXBI5hyXpx5t9lAcdBXay2M6WPcbplpDVtwvlR2rH04EqSizXm/2r35DNyI6S3SjIvPKy
ZGPEGO0hT9tvvRy96SZkD3uxtFDbOFHKivJReWOv5m0K2giuMJCEptgPaNkNoQDqZekxWuwNAQ5+
xekyP4OOJMauF8j2/Asso0ULWm1SqKVDD4AWEaM0lL5aqK55JQGjzzHkFL9/I4bwIBBG+HT1Ny79
fcd+2ErB5u937ssuqiSpRBZtT7+/WW2X/IG9Ny/wFwgrgEcaEztVNEFGu5USSfN3/F05HfjkfRy8
zowVbRzfihpbe15Gv27QXJDxTURVAyR5tPp8OfpNOhsKKrA/2fMAotqNXrl0Z4EnOa/kZwNemfHx
ww5RVcLEnsHXGkFXiVSjfv7WfjrfMluWPiWNZlDV9OCPXOenzTjHwcqB2TI1PyFUgQGrpPV8Ap7m
nsECjoIh/sYnmdavMJEUDktzDZRxYufOZgyyGOzVKw9aoLUrV+6BYqxEFNpF/An1Yuz0SKjNVr6Z
8Im/J+/ZgiWy2X3ZJv1bCCZ1UAHi8DhALZ9CGKukflGcurT6OYIMdRzmMGdzgAnIqduGs9HyU9hJ
0LxlzRCnZvxDUOy/Ri0E9cBnwQbT35JiXWKz0QyVIt1ydwyRarf/buFtSq4C4RSnRJDqurzJM9z2
qZvLXVtfkICEmyt0NKeBBXX9xpk285/Zte4hGD15blGnlkX7P8PoIaK/T9+qwPMKXNNz0p+5mZ9d
F4PR/N8B9gR1Ua1gZ8mC99J5KRU0tP2JKaEdOkY6vhf1M8ii3tJu4K//WsvV17AD0FJOipqAgdqP
RoBo6cPgMkoJOmpLWQ7IXgu68rkv9X7Ns9O/at0M6ch4eCZsjSvaOHUz24M/P3aBmBrviMBWbrqa
XdYNSh02/NEhZOC4qzZ4wZjF7Bi4e3G+uAcKN4zdQtXy+fBAMSebmmUY24rfAjTrF5t3A+vSqeDw
n9fimi4I8bHfvZnbO9Rizl353lEuwF3I85qnLd1Efsg1mL2eZEPXiQ5U9v6O8LbZY+NWujnQwcx+
aW0vg8qg76PeDXgd2qQjAdgx9+7VPingT1cUimSy3ml7MgBaYe024hi7QlGQZUlPpFPdpYIFPThJ
inMj6/NKOulCR4UcZ7KDruOy+380p8VmPLdWjO5u5AIcTjQ/j7h0wYmvRht/rUiPntZEx9p+zkI5
NU7o/TvAfo4z3vRjZtpxJBSuzQT872z0q5c24UxfTBagEQH7OcZF26TU+mxc5Tfj1FE+2VOZTc4e
+RKZaRL9d8JxhcRve6ntluAqRbtQHNjS3ak5CMD8d/0b1eovK607qnwsfhRdGmeRr9sFwSRQzGXh
llys8A4Y4/wXvU36GDlJlIFR3c/3szuelozleosZtgPm4oSgf6M2tqzn/I6ODMVbzl8hwjIgNbPf
PwI2LAa1KBATkRsk0U+4eDTYXhQTyCweOvAUWvwMpJqRSelDDc3toklpHzfGhqFDUfpCLwAcB6UF
qb5wgyw36QW4umQlUZgldfQ79F5uao1Lb73/L4gcMOFfDiS9ZdMwSkH5CMjgqpFOaB0KVGP0dvD6
RpS5QL++zLMnGIg/GodOIHaNYidaAxtmcqEW5KqqR0OgVU2X/IChww0GzGbwOqATn6t+wuFBDwfT
fY2VXCul7xw+lIBQPfCzLcj3ZYRwk5NEpiD80Vof9VDWorgP+xOseM9UAey84vVCKefFWgyKyBUu
EUVGCauSj01JAiJfXQfQ9herS8nFrUo7o4zbeSgsqntDseaqNYd+Ohs3m1kb36xArlJJdrKZ3YnM
xoypf9MFaLSH2F1CAI5FWHRbBPfRBQEM224ZIiw2ZU4vcvrfFh8nAzvYGstCUxF7fmhtd6K0HaQe
tGrilJ11pyWVbSS7bC+GbQyHaER6q2/3+1bjT3U5SmBz+lIMFj/KWYpz0r2KHlTItip5eBtOdzsO
D6E5Woofpdue47WLYnRLztrzNAFbWmnrI4PWtSwu7+FF1nt4zJiPiFJ2xXY1wjqCqFR1+LhbyMGT
ocePejYUB1j7WglSYUPOThgLkihGYRgv0u8OzBBiDXspYNtBYursagDE0qFa8n1gznQGG8fByohE
V4rmk0yuNnOXLnz+TYLCd96HPYMyj9S0EiOyfNpg8tGiMdmKlj58KGvmZkoZesXHsu4geHk1wzmp
Z3GsW1QRNU3JtghtUx8bzLDMaQhqiEEhE99FzNUFgfKZVXuRSBzg+GvBWmIuIyIB12wG4U0330kz
mBxUtXVchb2TUrlAJTnCx5a44w0ruoxJTFdLyKhWLIUH1bhTbN/luCGtB5UelGYT9RmHhZSLHuKK
GBM9yAQJD1jvUVVL4J1/PxrIneHxw3wMXmrnC5NVf3D6QFZjRejiLqKzhvEG867x9pxWgYD2zChy
Et2FlpJ0PyXPV40wNKEPd+2AQvZwyE8Y+cKgnywEAyy0X4xoquIgXXjn2x2eOQYj3R09TvdvA033
CcShgGxzvAcQGb1rM8uC7hOOxy6HFuNgpCS1KdOXvwOTi+DpdduAI30D++2hx5z2k1lea3Zo6aol
pOAl1GMr66IDQjdQd6FyBxC/XsjwC0RHDtB0xsDcdUtG73ca7oXwlLy412CRYVEaVTBQqMG+jkM+
K4Yj4mNqEAzrlA4ajF7XYzaxhQpOgR/vHzZcH7+De1hEWEx+8Lm3eDjvM1JBuUBk1zWkPGBQAE7Y
u3xrrQK/eLtQ+yXS69d3QgUiRKWCrOjkpRgwu5YTnhMg5jD6Far25AP6b8rZpBam9T/p2yFUrKhu
Tmenic4RjCygffeKL+0ZMOccFbNRFma5cn0wIYLJMpNtQDQKiVgBVjezTEfDLs8O5PLQQdW3OusL
Awd0+QBhAeAG0YDedqBvwvioq8fxY2g62Tl8pczwvKYK8m1huBWnudFn9K2ZMjtUt27YJaMBz6dr
fKN7LLFi+qx5vnITzJqih69yS+5A+8J159FCohhXLkoGIlGHOcMV6rLBZQArUgUzyYy49Y15qRaK
paziWIxktMDIJppUQGM1uXK9VkgRwHPIUc4aneyVHz770G3S0xYZPbYOdWchKXbELquSpCUePgEe
fwOzYdS8EZP60Z7uiM6NsB3ttMihITCaHB3kkp5Tt7qp3NGvAkN36DZvr+siQjVzXPnLCQNwcNt6
h4Lm/ounq7Zy6I6tgzDOftmVzKOEXLCm0YfuVxs43/JOzKgw2vNcRiflnxpFfbKEL3oulqBqfvQD
xVGJnNb3q4LGFhYzlzsW1waGBql3PXat1rZGHRzMI7+/hoqsEsDK5VFWNEEtEihcp3x0nFDwl7dv
k2nq81eeSAQQ/Pt3kf2FHOqMgRMNYUJfpX9Ip6H2DQpcAFNjZ20No3GKbZJdW8pOnZdTiBgCrEZt
02uTLXL3XnwuMKEjZp1a8ythZUc3g0Xf2Uw8M1g8AQ5Y5FbDwuNfTeXsG/B6g97xLlMb+wLbh+Qk
ZRBYt1dUNU/yOKOrOn2gtN5abMM9s293m2KfnMjDMZzofHMcToR1/fQQ7KLglhcd8MCjirrSQkuw
jcfaebFb87cBedFGqW/iK1ytW/SIR5KtB6DLSt9bvgmExQ7a4rV4tT5Poc+htIEFGQBLQUEh0xqm
P5fSL8udMf5WY2v4xoQD9xxr/m3uuWtQpJGVJPuXZFmi0EfANGZZAnioPZBbIeNl670oXLtXj5yj
DLIAfuwMAtmMtRIVx6sYyNm6TL9ljp2dmqPGKmZz4ZXfQXbKjDzB9LQOIVs7Corq9cfPEWh5WnUR
3XYcDeuazpWLPWtx8pWtN1c8qwJmWk8V9BBKeHo7q7c9jXFrZ35Moq1DlRJ7W0I8B5FmXy3DO0Lq
3kJY3E3aPNMa3oBEsTptFPSWzSKLUlblC7VWVkxtRmRXfVJozXrwu2ylo2MjOBBd1+2HVHgl3Sku
9szEWzpDrEPTbPMIC+xmfBjyjv74MH6/v1PfocgMUQEin9dkkRENoX/4gKMCOMQSr/zuOHPgYezf
/9mXcsJJmOGfYWdlSDUDeK6ovatkXCCJOhsXfS+PN/7CH2dLksc0wZRSRQQmo3V5K+FhRciOXKaN
LLK4X+u/4FDRyTkiJZAprGORke/ox+hgNPCzW767c3qUM47slQMSuuBYCC2ubRqHL75iVeLtfqNV
0Wi/+3XCPm8DwKH7KKFJUxLPl94Lm3MnD1Gle+K/vWBo1tUGKhXImffPuVNnh1GVyg74iHMnO+XF
acl4WSf9AI7thD7qp4YSK/AQvIMIZMTNyWgHXbZj7A2YAAzHUbOxb/SEqZdC85nqtQhZLCsCXzlo
4h2JBn1gH2rRcp0UqgGPIb1Y/Mzn6c1qhseDfdEVezN3v+DJL47T+42ndHQY9lg/bk68on+902og
dunEjfli6qWw8cC/czawsBuEALRlLkjIwCwdKFvjrGI7RWRX+UqISnbgAQAER0H2NE7d8Wv4mjOC
3EvnZJqynEwNcebleGRe7kTDAo+yWruWZ6Wf18HfidF4GUR5oWVmkt/ERCto36f7NQmm6+Y7Wo5r
dMNkbxbp05bf403gDhC2NTZryNqe+aKcIzOURMq+aEp/Wyva6OMKcPvK4teWn6ZrkZ+n04o9HjIE
MV67sfABJ1G6UG/3qou0XQxctp0CLsx6Ah3KVbvF8olyj7yiI1y31Jpc+97fZz0ce1VaNB8l9NvT
VP/waPb+5KPX7OC7pRQllfYV9W/Z+PDb6237rtrFeG2owVprQUoK9pksb4c6m7WMJP5r7vkCXI8W
lzeQcgA9EHQQe2iXw5zCXZ/0dne/sVay+uR2SZqCLWqbTmUtcuED7EbZrGWSMoe0b9wgfiokhaDb
g+65pLoJFl9su20TjmBDw4nSFCa9UiW7czqBnmHUtSIQQ9lUzSV9dLL9eLBzG2bh92On3XtCe+Q2
bTauVzbAOCX5ZQWgcVEOwOvXxQHYa63zBRjiVhjzU7sSidA+YF8TwYSnAVOsk0W5MbILQXQXDT9t
uDqb78oIJf0nYt2s5aw4NKDWtv5M77mthqyEer1dy+sIXaBGRswY/4d7RQmkB2L/aOGu0wco5VMY
Tp7MxXbr+y7iGzjz92CoEmVd3F523aJtg/vP2tPWyNO40UEbcl9s9Cw/LEOyI/lP84S+MXftVNT9
tMVLEMo2/pat9qthc6isxhW6G/BOnjPfgiRcME6sZYBG3BMX+HlwXxeLfiVJoP5MEogDGSy2hpaa
umS8ZXAvNlQy3r4codqpBu/PoaxKlDH56UpQdiqnj8skYCd7aQXCRgx9lNg3YsB6LqyxzSkafAZU
Ln9P3XH56mPpGHnYPga4oJ1DbYstIeg2B/yW7wcXlogew0mo2F74sJ/BMLqc4UtWAgQ6e5CLrptQ
ljVKqbQKCbVpl3ZZhe0f6KN0k3cLFlmuXpwhB+gdo7tZeckHsgexHkaVt0c8tH4r0SZE4qsnuoRx
lSoYuf0zb+9124QoNmjS3lAqswo8W6ze8hR5iObwqDgaLxFr3yLJGrDwqrrrryDvjeWNsPZvG+BX
8MipVDvCj1HsaqHoX0Tq1xawKifQ7WlIV0u0kYa8mzyV0yrzZqCCK4PHHNrgSFBE3JqvBscmHBUG
7Sjq2YP/elb5F3alsxPN8Qqqec+8e975xGXhb3LawsUDQhI0L58xbxXozklOeu1aegcNAEeu7ptO
cCOGAhaJBvuowVaJD83pNgX1Phns3bYaY33yhnounLJsYvgbNj8V45Tu3UbmnN3DdN2KlXM9U3Eg
2j9ujNz5rmg19Wz8a0Qsy14ozj5IG5CvxTfAu501kcEBiYLKNW9xmTO6fSGZPN3a57zAiuF6YP9W
rfiNXcyiClcQkNRx/sLH73qOFo3mMiIR3S3BCMjmEap8OrizZ3fZc95/Hl7vzEGnmSgAL5BZgYc0
/s6+q8Xo93rdd5CAINDYm4PrdIKA+6tEtnb3t10uqrpfTuc+MqS0HdMp1FSmTQ80fkxpgGF7eImi
ATgXXlWXF3CAfjF/sjhyECMLm1+QtK+GsjXK4txJxXScWFY8tv57Y7o15Yk5Q+r9aB29h5ECwMaW
gT7yO5MpQGP71Q4dhtmNuI1+Kehu8PGpEggdHFnrGruzHmc87x2Vo76N2YfltK7q1wx6DDHMxkJT
h4IaCKGAX/ivd7TEmtVjB3IfkPUGsoM1o5JbmQgIySdNQorGsLP7AG+MRUwg3KRORwHwIOshh/Sf
eC4GuSDVNKPq0ydQ6oo2wHSfEpatKtnAfgpDk0TfF1YRS7ytMOKR/2MtcORqHDOslk184Gp48h0v
KqQCqZLCJK7+CX2asoBCSOhNm/MMIk0DykyokF8QTxT3/WEf3+qXS0RfLAt08jYIM/4pzDyqRlI6
9HF3oNqSuFRhuirgQi4sy0iR0rqkBSraRBwuX4ypWZoe0q1HvKyX6BGXu45P4q2m8ukbj3BKFQ3V
i7rLsAovHcjTDJ+TgRgrSJro36ifT1WqrIjOKFUnG1iwvQowvAOTW2eIUqEtOjCIMTNMbpZTHOCo
lYsMB2a5I1Zgjled1cEVlLq2LjDQuYdXyEUgSeMV8NFlL8y0hNPo1fVlJKnJ9Sp9x62KcTJJ8gCG
uj7aLWQAXA1vCJ+BvFk9ij72b8xxKPOxe1LJ5KGiIJQULb8cModPkadgIRUofrG+PE0rUD9POmaE
vgRjPV61j0EblvSN3ZrfXtYUiD7TGDqxnku0uzGJbZcUkjruvpULuccp8N//z3sVG7JuzPc5/uXs
QlXWYuiuNs2qj2AI/FYuGUqy9LWBFocq2MU73GRHOkAcYgITZizLqWWf+y+ec+Kxwr0WcoreIRsK
2HDtMQQ6FSJzRQLwY/8RhrurOaHfFvbi9qKY3Z1SM9V9Z5H+Nb1MQioNUhq8w4IENim71pO+wAze
XDTMKYeHirqDXNQmauLrwppZsl+xnfgoIxV+fIHAK9CYDb//g718IylAuyWgoihabCFqcN+i6Kd2
GD9wa059RweDt2yz8VJoHrCiw2iOPjze16nPX8JrBGOJDA26f0c4UIfr0OLQ+e+oGfZHSUjFaxXG
rVWUjmLT79crEH45yBtCjx7KgIzpf12BWUh/ArgZLmRkrja6jzF2YO8ARrBDVntJym3JrZmvU1X+
+CdcSNL35Y66cG3M/0nkXpPfyDz6zKiQUblELmmx1Ukym0cfs7BxLWKK39tDM9P3OP/n0JQvdQvl
bJ/b0atWH6AIE+InhOoZW8dUmZqw9MLY+2Aa0e7rPg2XEKHXbLZwPD8xZFCRhI6G3JkbA0HqYRHO
1Hvge2Q+2fWs45pnsjR8zvuycCUl2Xgumszz//ZHT2hp20Lt+CzHvhEwMyrohTU7ktLwtg2VQdQC
mrGnwtolbTSlkdG7Pyzj/bx/NTwtoYwrU8/gEw+xsjPEgbjwvgTjFOQOE36SMY8cRz169WeVPgcW
RkrWObG5508V/VSuRhY89GXCLA2QsNjhTE9fPp6UztP2iXwF86GPtq9Pg/Mc+q06VQHKOmOic7lt
6zhHJZ0XrSk4V7uC2SDKAfDSG84gfpWpqPaZyOJTsIxDqOcxISXnoxOCIW5lEwf0ftrS/rK/LaMi
spkPrpsvEf1WzUrEwf/o89h6JKSiL6AWMpFJDmrX///yWybLe0ONsvK/ZnilK0tCbUafPkCaSQkc
Rsb8wjWbr92DM49n9c9jVYmLlwyeyluuKii/hr2rS83DGr7Ola+cmgVgJkx7IyxUFvkXuI4/PnQ4
1ImCGN2yNl5ugj4CJ+T9GEusjAte2qO6f8XytwKf5P8+oAgi0BrOu25t5nT5peQjF2Dlgcd4zPsH
gDKJKVBAFftyqz6FDhwXz+C/rBNRyPjpb0gX/mNvVz2n3NhGzG8fmss+LoP6vSVWUvAPFOVGWO3M
jnTqTuH7hYZCkrjuRDA4NK4R7Xfr2MRiy0AbY3WLFW7mK904WYpombny51s/gOKU1WZU2cNbfEe8
kIkELzF15x/P14Q26107u2s6JCVbTUStuXh1A9CldDiS7GxTB7yh2a/9vRfJhuJM7vShP/xsSrPO
iMjDJeqIAXEVTd+gw9virFrK71+Cmz1MX9R7euGWLU0svU/JJ99Ay0tp1yuHzn96KTxdS41RCcFK
DnHoF5eoyLesGUgi0Vnv+yIBvaXH/X1uvm39B+oqZ4QQ0/nbuZAda9kLpqpdIjHww1mqwWbGtKkI
NOmUimtVb4pEgODCluDuDXjio2ku1rZnJ8L9wY0AHY1C7dRn2dYX87DeWRdBvfEgTLMLpaWgF8Nh
JHYFzNXLoJtPPpJL+X9FC9ipFK78i17GqPpTpONOe0BULsiAJwY1ZvM2YH3yueqyQaeS5e6TxO4k
hKgq9eDs4md92dXZUjyZDXvhkSTU+N2ay59v4JLVHg2Rskxd/83SzTtbWfjybM5CV3TsOz4aqy7K
mlQ20qFmVeiDoEhjbQPBT7lFgAHeqR+X45hRKSJS2QSIGoCRTTi4OPMAPB5JT2PNY5lTAQ/hM1er
cQBJO6FgbIQyr2W2ZjC70Fr3CwjnJNXhSunXWSWu3U6qYFl90VrL/md/tXSo9qibXRADteFIZvT2
AMDZodLMqrHAbArqyEtZu4CUcIZmfR4qcDnPUo20uIqUXWlNZbc8mX/kDL+SFXxKLwHPE+jMAM49
8rnSf+63W3EYlkURvbuUKOpsUsnPYPD/3PYiC5ubLHCxSDu1n8z+23+O/LEhNvCuMGCZOtOfCyiC
6Pl4kTla6sRUSh5wo9PgC09AEG5FuX8/FucMb+ELqCAIwT+UqCdGBPPnBDZOIBYDaYXRpXyVQPmo
i4p2rBDrduZLEmFwFd4H43yjzpW8qPxIj86VvLoUpZJJ6gPXZhAUO715yaoMa3jFpREhHixv1hpz
iuGyB+w9oP0nILnxxngl0NvfqJJgC9OvKVrCSb1igl7RPyT5bR+P2SyRRd0L7/hIvL/+LC97Np2y
mu86XTy82+TgyJ1ukL3sh+oFQml4032NrnV9ey8DXE5MnOACkPbBi36y/WnksScPLgJVqorRAy5Y
yHIEeEK00Jzdiq2mCXgmh0ginlQwJs1KHI/5Ceu/L5Tlft86mMbyIaVobGx3iP/07FQ/BlBfk5H2
KbGTGVxCskHty+vsQvuaBIGLB4xPXGST4HdIIg0KIJgBV6yhM+X5rWsZpcsHe6q+C43myK/rU6u1
3FP4Ez3ozGYOMYHHnB0aBDbNojwZF4ehBq5fePTLbl4ibn3xHncY9k3FtuW6w80pa4E6hwvTvq5b
+5fnhlJn5fG1JRQY3jn4P62dJ226gAuXAA06BdYW+UuFDX4wKoSQNnyQdKK2PY/P1aixUSfDWs0h
GtoxJ7QcY1XE6q+X47fZSAXZbyDjnbAPf6wS/VFBiPi3uzFgWLwGrCi18XHKmc5xaeI1M32VK+if
bzEKid82sPbslMzdfjHvmogIQjsbawueN1S4BoWN+xjGaNy/RhXmJyzMsg0P/zfGd/nZH90H6o1m
p5+bLERr7+kAdb3IAEVWQYzvaOqQKahAVaj5lbUtwnDGmsgtszbyxa+fQOCXoRGTTKIzh/oJ9auq
S3vU+UJoaT90Wp1jTPBDnNlq37WzTIer+HLbAAuh+5Uk+oRxQzSsHpS1OIf3BwT8SBau2FLOnde+
goVldlDJ9ONS+T+0DmX83PlU5ZCRUPo6SCIBRxTyVNbA8KyYAYiwKzRVvFe8masxFvfhSr1MY5Jx
JhX14/DSENFpKO/vdoqrvCztR+pRsrJytJm11E91m/ofh/y/S8t1eYKUA6pRTh7SGXIyXg+YXHtT
J4fsKs8keN1MjiE4VPrV4pmRUOjGQIzrde7Lbgb7Nr8CpDRVqpx6koHTq+lIplu/5f+/SHaMUEn6
fQk/DGUBLH7dYuF7LrGK8p/JIN27Lrx4r8Cge8N7nDIlzkdik2wYmBo8/wPkPs3ss4Pp/AIvzLI4
6qmT4Hv9ukz7KJ0vZX+W51uympWopkEvRedhX12ucZb3F4CbXxfz1FMQCff4GSxTyG+Tie6qeC1Q
caVaEKmVtQyKDFfL1xuFGCVDcTQ6rPzyUPv1YIU/EUmdHEGaDfwrdJMrVjUtELTAL6ALCRPX3F3g
qPw00JJrLxVuSJ/9FpF7S9DJ23YKG1NsI5xKNcOyr3gR/TWIL9LgsQAyA+OWMaq7EHj5F1GXl01+
DabuK1N8bOJTxGmMpMywNFhBDueUm+59qJcHng7JpWFL/eRAYQ8VOF3++toNglrkWTcnxGPG+YfY
UNjcw7gS1VPHeuJ6G01ERMbhq/XK0SD566bBY+B1yw06pcdqwcmWEmSKBFPHd5u133p4rf8jCqUv
J27pqeeybuZ9Fb1pS/pEGjfc0EAwE4jvjb0lQ5iMrNd7KDf/GUYvnhsMiATMC+vokqJWJybwRjAz
inxaBsBV17qlUwq0v7IbqHS8UN2Yc/EzUZhm9Fej0yYvXnou29tCXaS/MEx0XTjQrOXrBQ9ot0DH
ZW3ab27KxmMDF1iXlo7qOds/WV9geESvuX9KRgCH4OiULlWaHI7qUR9vdE7Tn7mfsfucjccVrMke
8KiFhiY9almr+/PIyb7mqClI2rFF/NcI/SYk+BB9WcNo+NinE2h1lXo4/jVxewyFQLE8E0n2GDqn
bg6LWkxTWRdPXSHzw3aJZz9RKhesACCauHfyUHyQ4KlO4V+A6NDeCa3iX9oo/NomJgus3cC4bPdp
r8z0ldHA0mBM6v9iX7GNzlgseWq27dR9Hr+XnVVn4AfnK5jS/ETW34qhd6VawIicNVzVh8Gzs/Hb
Lnb+Wu69Z9Qd9pGzuh7qAayhR/P3suHTMHGXMaadR8gkFA2PbNVyNmZFm5Zu++2JCIW+KL4q1GlZ
Msyfbe5Fey6RZEMAbmBy/IAQ1qmSl2nc8imP2tSXz6EvPirpPfMA1KjTL4Y7uHacAIPhP5f8NVuA
ZkDLQ13f9eyGVBr+gqWJ1dtwyN07FryaEyhDZIZU+hxr5F57HXbf4a03eWzl9fwepZcH0Qar3ofU
zIYB8wv1dvnQN54GOvUbw/fji9khXuw+WEjLi2J/Y60/Hl4bLkti9ihaHNBTlWsiBuSEIPoHy1XP
EIrCRRwr9ldCC35C0aun2ElRssXRLKZk6IHvvaBiBk3OEutXEsngpNT30JNfqvLPvevDQ9zF39wC
SaH5srAMJficFJwJA/F8TrHQxa6aH3z2zbT/YwbwjB5AO2zG4/UWHFu38RfVtKmh6VDinV3d/Omw
jYHuGtNPnF5t5Yf5EicHf712nXXnhaz04H7O2MxRQ7lRw4AJlp6RoevqA31CvgGxYvD0d4OQlQl3
oUC5vM9r0JRRKumCL0EXAyU70VCRZsvqj4lLyVS26T/a7UcdTObLASKyK2EZ4VGPtpyN8qMjkpGI
+2mQMv61OddVG+IEyzW0B9h6GCA8o2Pa7ttqTgY2wWXfn71N/TQ7W6Rhbg/jgH73hthpMqjOX5hX
M2AlEKIx83j9LfmnHKe9OYl0l+3Gjz+K9p9G55ZpQ314pEkQFalLLPyDUST45iN49SXEkXkR8Y5b
Sd7XyC7UoQfGE7GgZMdDUsMo0Du2rXVMJNt0xjJExCR38P7RuXwocf7Xuh50KDg8ztkoG2nYxcOu
4dOpwp1XXo2PyGlKVEH6AIFL/yLGWakBD70pgP3k3uBYosH505AfkAy6ukQiYBb4izdEJAx0t29x
YuYW8dwisoMbC6bDJN3oEGD9AvMfOTxr8cvrD2niJeilAQcoPbbdZcRhAaJ/fVXwv/4iyLOOCY4k
FlMnj0GDC4dh3bTJ2LY7Oe2kf0JFoq0O95UJMMoKuEwU4qB+dsrfvO2dI8tXWbF3S5zMNnWc+ED6
37r+paqICTzwGILEtbRk0CS836soleTPDJ+QUARFURo3S64TDB7blcVppx9FBi1WHDsgI12tZaDa
9aYTV8+61nW9Krcu54eogPaprk6ctzjLnKM1GTTxSX6qAEdpwTeQiUP/dJxHssrnApLeibvCsEKp
CgUeBvUuVITjVJ05E6SU1S9IogVifE0UcmzERWxB2l1TrZynl1S0MQKNzfhdH0upS5DkjAPZitBQ
fJbs6BgaqaPVdQymr1xe3B0qEqKevumk3q82rPeirCTCKZWvP7Z1ECPJUPdUqQ7iwUVF3g14WiQT
iZU/8/Esk6XdBtk5E9qgWJXfO1xN7L2Q6IfSxT1Obi7DiZRpMHkFPUpKTKX/Uamca0Yn2H+UoLQS
ia6qT7UsfSuTCVCnhKVJFQVeYDGddWWljr/XAejRTqEOnOklaslUKn36pWXuWJy0qoPT6nH0EuDW
W188gBc7IXWf4RFjy90/h1TYyNvoAgJMmhIClbCdMSV0mqIRRCDmpPTVh2p1sIusvnlue6qK8myd
V7XfDxT4YAs3NQ22PbOpEbDOKgf1UsjPjooWGlIKCOH5Ny8KkTZFy1X22j6Iy7BtBT6vTbY652UC
DoP1zT8evidNWh9Ed91MgwpmDnDyU7bWAnWdobGokF90udRdu17dje7sahb7Ue1eo93ofCDeHSma
u7ASrVQueYvMZQlh9tzn++DKRkEHE+NY5rrjMy3AI+W5HA3G+3OezHn6LLH0lQ2r12A8byqNrrH5
PGW7A/PyCsud8LzZ6rtCprPrdGlhO15Lp+oQHqjERvh0rvFIDJsi4qJGZOfnK2jVSUFD3H5R+alM
5tEeeBdS4+XAk/cFDzISLlDIga8HOd/7XyB9wQ+KoDYHGpArQ14YqX6dgIijKHEGfYBhDlAhabjq
XTO06//zA3ZJXDGx7M/4WtipbHy7XTVmcrW9A6h/oPbFjsghsIs0r13rbgXhacTdX6M7h5XBvzbW
RMF+cheTRoe1Gz/kRPIBiqVNKnDhFbJ2l7Dzpu2LS09xseKtL4EtwB/VXefT8seV9Mw5BBn5tYu2
Nu/TlLIxRUDZSFRNMKZlSK9diBV7SYlyCGTa1pPWj1QL2DXQEdSIK+XSKOJExgaMg1XED1ObNpuR
rA5TTbBQpUWLFj854tHaOtkfl8o3K0F3Rxt/SswQW+ZJ/6QmRu2F5qphUVEWO5EeSoPWTW6PKyw9
Ad/W1KmSsLh+5afWHfvasD0g25GUfHS8vJAej2WuJ2QN2aXPPP6OUfG7g2fHouKe/H9H55BUkpCN
n75Xl1zx8CX1pVqtXjOTKzySgPwrGgBOTTVXxMFtqp8akp+cF6tjJ0pSaKEEttrXoNvOI0JLiyD0
8f9gpY7m45TrI+BkC+LAdL6pE9RZU7ZfQ3GE6yqgTjXT11sorDvD+LXxmiBCmJ3Bhya0H0MhE7Mz
gqyqM1nzsH7eY6N3UveWww2AjDUFpiGAuoKID9aWphq0QjYuwymInDjwd0NsEPMGS4MLwQlbb+y+
Tewdn00Hs/7BWfnJY3G8pmoZSTOSWhtmHj+qj/OTaP6wRyHKqpiPTOmzKrmlzS5c50YdBg0hx8tV
vQNC2fJ1iyQQ4iWXOr7A2GOUh2iNtxRYBcrLQx2avlLecE7O6fquE2Qgf37gtq8n6JFVRsHxCE8F
0AUEVjIChwTxk3XKViv4AZXGjv8lu6teAOOJp2naKeJJ6AXb3ojB1X3hD7hHL703fkprL2WPT2/w
hj5ytkmuRBQ4KztIe9nRrr6hqjUOh2tUKYV2alN7QXcK7ZRSQjV0BeBb8fTNIedDWphGCvLBaIjc
ix5qXg+rkWpXZx8dASAZeaRzYsiTU1fiHycg8fTm59X30blH67lKslgjMc8S8l7W/HSHWlKmNGHJ
V/k0rlCGPQlFDK6uji4aTZBCod5rF/FgchbP0jOWZ2+JAR/RADes0WuxzML8k/uWwLfTDXALDeoK
3cSDwvnWiEUuAdIGeE5y7VLvaJUQsNGBEOE4nYl/jyGnzyqhuhBWmhS4DJkKvGqNBOgk6PrslUB1
FLfCdQ248DtJGNcSTPQPzh+1xl6GeD8N6NulvSCE5LnYStS7UxGsoWSai7LB5QDKFKgZq8QD70Y1
2X7b78YORx3ca8MqjzZrqtcdnZTi2QAYlt/1XXUYYqpQv5faNTYAY7vIWyavwWyZZ04x2kTHSzMm
oPd3pYGrBbK9Da1kV9hmH4lMDOAQJzUpDjwpDgWSJK9DCBNFpzQOaSfMgSX7huDWZS4iQ8bDAeyF
hEYzHr8KGbrsi5dmDtfOhUfbW29sgmWuSBGntm5CJD/lwP1smHKiYlCBPin1PrNnhVaSRfFLCDqs
rcz7iAOJB80tQD2EeO7W/SQIETGzqIdzqRc0UFtdos6gvOITP65jOljvpNq2rNJllghRIJEuLKtV
ls+bNA4Dx+s77pbRbcvBEgT/sHvkE7tipAfzPYOHnx7Shcbp3jehR1o79Z7hvVBrhAXNyqE3WUsR
HiJQ+dNaDQy5F9OCy3uXQ4fCi9Ny3IEJ4MmTVRCC9xG5xsNhsHtcJouyqA2sp3AQWQ72R4lZtUnQ
9JJe+DDTJWDvZls1BdDDIfukrTQhsn0l00jVHD8g9Cj4Q/R9/7tSAel9dwhtnShjoh+LwSZP1N+g
lysdPMYOh9WRtcDUbFXiY5Kx1+NB1lVHKsRGDr4+lWJicbJQEVaB+c2PQKU4RCa8xaVfc23BQjYj
DBg+O72vQ2C6tSsbVJYfLQ5WiVLmPxlU2aBahCdW7Q8cnyQS98/aSkWiH3oQu8LmV0TkBROVWIUz
01E171VKMu9GEEUJUvd0NEaKmVzrwHRZVp/GdCzICS0nvcEUmuIYFycMOvp+xmdgC3P+2OdoK60L
6PSdGjgUomR6VU0RCzp4pXYsqKzCK45Nw6FOh1qbGN5RBar0QVR+2/3DJNFnvoCHV4sKjj/2t4pT
lc6z1BZw5HCAia9u/wucrpqQG/o7pNVvTHFIb7gaeZoNEUcUvHM0zvsndNZbWBekSRqxRvki2lRi
VbbeXj4OLaKAogTBwjbjsnFppzQL2WInffOVzFX3WM13VARcHsB848zTjiHCdaOty4HS0ZgZCieE
NvwBGECpuE8ltgn9ss3eROiJZBPp8ggDhsTzWR6C1AAEtIzj0F1tNIk0ubXKaUzFusgFMwtzUhJi
mhgQIawFxfUIIQk4gyOVEVc0WOrMqbHnPikqA00bN3Ko0/I9cYPAIv1CchZgF1SpcSNqj2hKuWnl
DZbNWVqq1B9ZvjXe5g7bfTCRfTmE/zAkakeWUcnbZ+NcKgR1oV5YVXdo14RvvoktG0OBsV1qEW3o
sft61AKeGNHBA27iz0WjwdV8xb8R2M5xdQ62qbNTeg17wU13PYO8GnBndAy14FuDF7QPpp9Ob2cm
rA6BG5sm2jM/6/SwcmGh5W1f23ZMeWjBOYg5MMFnUGljqHJYBkfUN86qW7Tnk1aqfCcu1AWenmVC
mRU3FvfckDKHCE7agE5EowqBCXhvZAjgPGmtdvEstldDvKUjqL/N/MDtZ9Opdk3aJMRz70TEcpdA
nPPeo52ESd1A1EDjBth3GrlxBE1U6fCka+V5AZOA5b/eLPuVUL0FQLsYzR9yIN9Oaisus9UfeK9D
V36NKj1veRzlRgXbCftGJ99slxu5q3bvEsqogD+5CJVErKpnzvaWmzkOZX9A+WhPSP2cy7CpyGMa
K7O6kZTrCoA/LTcBTK1Umr9pSNY7GttZc0TinWFcT7FuZ4SQwl+gRb/RC4ct/p/1iRMdv5/Yy89c
iggK4DmVLONZxTIt/jrErWzIV//ZiXy5J0SYy3/cbGkc/kMXr5+OdpPFtFxe5H0SDkgoVqZl/Q8o
gDUYKd9gJagVzWwgeJ3IqKrzQcVRsind0Pajn7g96yH75VvnSH7ypICBwfHW9sUDLtCm6H/OHKPc
jJGGqgiBRh/swsV28t2+62VLccjuVHS5Ols5aXrNKFU31IvsO8EbtoDkET8ZUTbYterSN7Rk4ME/
sAbK9w9f9XHKRjb/Sl/olFzj3t/HKMJxrtgkfcO9/KWpoBHcCXyBdoZ+KKVwKtma7rsucXFVWjUm
d2DeYLVkb8CIbjMx7QS9gCXgHuiW2SmYcXymmaqfbmrSF/rpQq9X8j6nEO4AGmxLaHbnwRfkqqHS
ZautQHTWDurMYUGpLbtyRpFYjtLowKmZZ/soKCcMFX3aR5cDwMwhTkczp+BLZzAwkTY0+7CMx2LE
o/LOUCiqZ4JMY+gZ10h2Mn1+26VNjO+2JCL7Yv42jc8ovpwkrSVhXONnY7Dp5xdn1sGFeZA1HD8O
4X05lMSCtoC3Fw/T9whsq6Vpa2KmyTjcCc73wykc+oxawC0ndl4cxY72MuZjrMA9CkVR79mA1KNL
C9EtJAmpITGRO1ewYRIKWEk6xEl8Sr4Id/udw4q2R7h97AvTipVUv+XXPNweNZa1ynXVBL5KvhgF
2G7xEabMXbP0At+x5wAUJx/WUaR6MlQTgJXtFB6DSRHzH8gWa+JhOSZjkydKv/RscPveIpYFG225
cSk6LwQEBbxl2OLy1LXJOwn2+0cKIc6itNKSF76m907eJ8FcmQy37u7JmbK+ptS2+P/qVM3KGMyF
1uIxc6LDLV0iLcIkTC+rstQzZwZLu4VtfArrsNTjvGC6CADD+v5raQjafXZtuGdVJfOgJZW13gQf
0hfsejFFbWCKiDeNdMBDLDGWqTNKhBTGB/sSdz76dwY3p0NO8vxGJ3h03wHd472/40AUBcAPsaBV
Y1x/OwroI3+xDIHT+X993vDFFbYBg+uzpsjj19w3A8eTSgqyivREGC16EFpbahS10z/OmgtRiGOD
rCRkfYLi8z958LBnVwEk/gbj2KnHEwJyeMTD+qG84B5S4sbyiAsBS16yPZIMDHarbaLY5sQHfNTs
nHm3xFrJqkj6/2PvrMuivJQGuhx5iTQbfj+q6EDk2QtVFswAvC9rRRDSwB1/DX+avO1LyQtHsCqn
oh5F/UzpRBaRPFGykHpcUYwPOxMY4Xv+xJ7i12HC0wcVfqiRkyoIoL4dIx64AIlRb0nYLANCz5J4
ndN5NMXldi5Y/nio3fCgK5zkQJAXfRNNxh03zkt4qqVwYgTy6pBGstPSUU/Q9yFHLP72NJYIuRlv
wqFcnCGkJu2YJ7haHVJ5ln6jXmCkLQ+a32PXAXuWt7hSR7aTN8RDoGxPOSXcTIR14WTUyn7aQcUL
dYgcqhYfuJTYGcPmfZvwdcmL5x5q+zz3mixk1ldfoCIfL4ck4h7U//h4ohVfexcVaAaQWx9mZ5b1
92QxLEOlasVWHAzTLPVHDmF77BDkBVCZjKuVfkljD6VNGzzzfpwZQTu2ZeiZZWkwXSB+Ya0wqqXv
rofCgkTuYnJOHAe6lv6hUAH7Q5c9YVuU/9QEQkjmSakGSxM+EIMALi5BojIB/qbBgRG8SxiNoWXa
GQTe1YakKiZRrEBlAb/nTSyGqnFh8HWNv62gdJQPtgPvaVr0g+B4P7oMPXIYvmSa7g7nmbtYJSOA
pE2hb2qrVhR2x5A77nxblc8FhSzNcd1oeY0PCRbehkcBOut2OS7AwOqLMPZOCWiOAMYAmZnUaq4W
2GMEBGDXfFkcdcIdumATFlkXKUQNVk/8SD+ZR87dziMbIb3Gt4QqpHYQ7qkTw45u2iHrVchRuPvn
bwlkjUX8oZBYgXkEZZPz5GEgn3jGuy7JJPk8sl+wMhvHZIa9Zked7QNo//S1CFdXol0f6L4eTLoR
1FcCbyQ+FCenS0dz4gVb4DMWG8DSVtimQP0ns2JbX4nNpuDsAsLjbGq+WCnZ+g11RrHEzUxm7gjl
PXNga22T6WulrudCRPknzKgK0Cn5Z98zfu7QgoUMG6IWfPlKC2JEP0xZxe7dB4Ow3S2NiGImtlnq
OSLFvXMkmfIFElVJZlCobzcNKj81UpHAvoAp3XvwcR+jI2eX9yknXv6s4UuvXTAXf+VXIXV7BYXT
E9UPqjE2CzoEVKU6sfZexacVyxuZOD5vQ/x+7zwOVDCYJ8b6zo43/z9mAV/qyz19monxw9bp1wGO
TQVYWSGRr7sZzN23mG7H4Vwzw8g0Hjpl5hu4vcUf9B4cW201wxynjbkIjDTk6sOOH2vrEap5raHX
Y4oJar8VESnGSMkxz0BMjJKtIw8wrS9BCY58Ha/Do811x9flBettMURxDvE5zDEZoPnHxpatOWLx
t+opfara5FQOz8SYPpwRwFEVsGGSg+RO6K4BBdET3lEWb92KzT+FAb3/5WnZon7bpZQq7B4ql7aE
HlLlKd2G3u4fiDlyzJ1Zorzu1uGFVfpFLlC36AE7CJA3c3nJEQDkqFvXB2nS3X/h2w7v9GWgM4+L
ymiQLoav5EV6+wd11WsSGt0H1Bduj+yi1QgH0BjSOKOYgFoGzQ/+kp75kMGe26oeqjQHUP7fdHMr
TWFcPQwvQnctaV97HwC7qavIncAaVsFZMGo/am2AOhtyV3QfSRNA78i2lRZSQ+nj8Q53StY+T5eK
gnDqOceim/3w25Fla9xbBWPqMe3zQfJUgvHQ3VEQgZhOTlKVBlI0upPT5ZburuAPDALzbFsv9aqC
P48Zslw1stNruWQfE+LYpebg1ahhKcub1bUSHAs7Q5yXiqmFpODC4O35Hofmk8pw1nTNAw8qxyy3
xJAc0K/DJVMgJ8hZhjfS60x2BmGuMKSExlM24VqqUin0gCYt2d4JIyfKRb58OJNzCPgbUDnsdWzP
M1+c2UQRcA3bnMtvl52ySE83dgzH293gBnNO12xGkXIYvesewKv7coO4S6FQGbrnrsaC2/5f4Wu+
SwQdRcGwGxKaSunvBVj2M2znbK5W5eNBcL3x1cq64Pa3+nyVJvI3E+f5EqLtJ1U+J3emNcLb8mKJ
ycr9iHZXUGPMC14pkRay25r5vvGgYDGFRnizYjsQtoYaQFiyuuVrY2TmJvME3BYZ1E3x5Hpwu6G1
mEMpHSVekPIWn8WljSPs2IvsNNFVvVwxoGjcV0C4dwBPeXJtmLmMk0FJWp6H6gmBjQiUc/uAZRGc
K9cv8BmdSo9eQ0cdBu26NfDPnV6kMEeNu1CKI5VGxxlObC4rFPSH+u6V/QG0zsPz6VChz9cq8SMg
eBUmX8R1pZS+UPp3ykKl+lP2o227aVWqMuC4zoBoSn7SDZRD+0afHZMd+e2nXyXXsiOdvRrUYMSY
amS0QgemXGdJDTRxg8a0Fdgjty8abeYawAkntHOfyVRootlueLtshRvN7MRO62BfnKUVycbS29u+
t7EHGU71IQztK8bsWuVf4JWTfktOk4+2SVPr3vKxwXFVgefomAWhx78M0sd1l2VlxztjbFIo9L4F
ny+QorQJ0P1z51vpL+dnbgWcEgLykz0fPEiDxcf6Qlgorr6gsuMuQJXJzyYeO7CeJeXuMGq+wyuD
Vmwv8ydRxHABZHZPXnc7SjeHMlXE0kpdmyYmSkE50zuxCFdZQ2xl0wilTtOFoRatV8J4uUu64A7p
xr/VmatRLIswv0od0slZ7dZlsO1yC0H7SLlc8Y+VgkiBY6lEgtlUqAesOmWBEfjElOtaFesbZhAs
tdOJ06Pscxt35YPYPoTtW7Ya06ZvhODUaHdHU59c2H5N/Z5ZNC0CJYwFsZxCNSfMjO1dKSObUuEd
AGZT6ANwFHVL254bjRzTS4ejtpgnT1Xg+cauXqqPXpRY9JzZWUJBV6g3cJxeX3z6by9mcUFsyeU3
UXa3H0aCYBMF4Zk+sx+8b7i3Y735sQg4bse+jGNUjZPe6fIsQ92ZHe9/YslO0K6eOWJ7356PEBrT
P3KxY8rTDnwUsFAe/iDQfXTWxfZkwMjpjRTu8k03rRTQByRr76TnFZs3IUd7pxGFRDgIDrNwoffm
y2UGzcjiySV50HHxJOi75Wflr44IBYm68/2qP7HN7SMPU/Sr5W3B/Z1vO3QzoQT9UIjiTCZCFt0z
lnQNPaUTa/Nmp+RvBzg+4HzI5sF2yjn+EqBnpKI5FeqfP/5pkfpRQyTYQb9/KGrPpAqr9WrdQXZ7
6cWzprIR/hT9kSxHal/FMi1x5ABpqJID/Q4uBdK4iXcRhacv0nmPMoi0qR2N5riMSpTo7FLr3B68
BvF1MvpUEB9FPQKd1XQ9X+Sdq34RTLijytSe21qd2f+lU7ss6/BJLZi2h3tNcv+CApKeApCywacz
0vrOIyv72ZO0Hb/TNCMzJL0sskQfVVRkcqU+2hpa9kgskyEAJTOfSw7RA2H9cUiRVBWHSxHF9sdr
41v5JtAzWG1kaaQokjz8S0OssgHhEX3M6y8v7FfxWanOytp+5dXk45Yl+HXG3E3V/fL7PpiM1SLo
iwvnklqy7YHjkXuycw/gxB+cpgcHn+WR1TZTmzXn7Cl7fQCNPs0E1Abz+sex68omdZx0TB6cmwU9
kDITgb4iRHvtNyiuFWQjreYfKjTFmnfCEzVAO9k765CLr5Xc/ssqlOsbqsyGKCktuhTyAQib/2ED
xK8XwFYaK/Rdp8tp4dO92mbLTy0hzuZ9oFrd8inqhfiKei/uMxyp3O2VjbdhlUwEL1NpQRBWyqXl
kfBLuHqkuv0oTs0AbBJNF4d91m6wm0It2EX6yk/WSEiGfR9vYj+3DPtX7q+mlCMfJRn+m9re0TtZ
j9nPddvJpPokfl3tC9sVWged9Yqg9CZ0Jsin5HgvWeg0j3ZE9xDfHVvxmYh52jD4t9NqL3lvOX3U
Z2xPpE0KFNqKdLXREaBRc0mRLY0IWjlWL+ljhGBroayB2K/x6oUMRyRfakXOwv2uJLdEBpHnFBHy
Bt52XM+zXRTem9ivPsAHgByWIWtw8gdrXRqjjZ6y4tRvFR1dNLKMb2gx/QgxrrdwHF5b74/4Y+3k
d6wYchbUgbf1EoTMgt9AR30RPe+NHLfMa1yMNt541Xq2jqiWHEm7GiYKd42WHd1QeJJ+gQFqimU8
rDSXyiy4C3m8gOxCK0JQBjk0tiM1ZGERawCLGnA6uSyq/yVGpuc+vS/g0niGf/BK1Lqhh9616evX
PHQ1gWqQMLPl7zn+qdDr8mBAao0Hf6aQT0JpFck2+soYNJ8uLYAtEOZdkSbuXuRtRxm8YLwo0U97
pSt3reoBigCtHoBiFJhYVOU7y2CdoxlNURgjSZ4AgYCjzATjCWzkQ8R19VN7QCrCMcBjPnHW2Tgd
q4jRiygCSmN/303DHttTdgm0uHe2RP6jAS14mKP9tJDfMMnU3WyLmjD9CPhbsn5WqCYO3C7UI3bF
rgBl+XQAzd+2z/0KTM/0ZZ/JAQ1AkEHqCScHiq18D1Ty4oEmgoCwTqRfqCkQZPfDBgT7klAZP4/E
+T5b37giXSBplQmJNmKHlDrwVQl/dyee8TUINDr38kF3r8ksroa1gQ/DSu33QWfJOlhAOkDqGTqz
gkWvwBV7WzIXrDopQIKps99TkKZ0IFNbKSRC5OIDMmUzbi+ar95yjqPJ+SKk0tV54Gw63MxYL9DG
if6H+OFJK8Wx+ULVOx4vvZ7gtQ3jQ9UTicd8w6SlTWhojoZHHppPQAK9KhM9/yYbe8gAh+6E4JTU
IZ/uEMutmpZHeTJ4DeFnRVOofkcQ7KEqbVZ5T6KxjosBG8NMsk69hLIie5gTmCgsdcFwQjw62S2x
Ti7NLh0TpXGcxAEH+MgXJFqJ40v2Roi5xrXiK7GJZ+aWaw6YZ77Dth6fdpNhCksAX6ECnJB1cV9A
SVXgrdjCFxiH1QGcw1TwmAXNyYXwzd3LtTp3WTGOfE6cGwx3oucaJMAdXH9FZAUhrYwzAS4vnsmP
sWA/D2Juq1qr3nMl2ZtWQxB516p/IS6mk/WQCouZK0laaTEh8Ik3mg1Eh7L867aQkP/s++gv+4AN
q4hL5SZ3xgL6O+6lPiOclJXRBMRczDepp+ZRxx4MRrOwMc8lFklIicPYnZRtA0CJAC2ZSBsj02BV
7tOHNe5wuQ6Ip9iu97moSDWfWXVHiejP/vdYxHX2GULUp8kyqPFhTxgjqNzpGrIdRsxU8yQOMBZP
295uwKdkxuaTNYIXsqNHXxPRx37CRP70G+p227yKWTUoeIXgFoPCiN7Uh4dNEuq455leNcZwf/M+
hr/K6oqXh+hu41PVQS2KpbNTVx7oxMxw6bsB12dJm0AVQm7tNMOa9+9Kb9mfQC76C2LeW6iB6yUY
uYtEQKDo8rXYtHo2FI++5o4fyRubcgLTLL4qne+RU+6xdd9Eg00yg29SQX/8KiYcrLJ1yszOeeNU
6xp5B3VsyOzkqrO+1XY1N0ShfzlzOleToLayBKTAWC6TajAoAZ/HTdjXzDnlEsnxBV3JYWB/8sO4
zT+IHKCM6LgB3JZ4e5E28IjHRw/n8ZyJsHx7UvxJ8o9oIP/TvH/oDwBamLwbTtFlY4NtMEKJ3Wzn
WhtnNi609vudN9upTZD/FBTRgRK3rXFoQ7FncRRQUAlB9ElNS51IRLLHDAGHg/noD445G7DZo+DG
qzImhYfQg3TwU4wgSi0g8HRjf1WT/0GCNficWy1c5xY9bF2MhzKET0d5zhhxKlz5eKalAm57U7Mt
zx+OmCqdegpINxvX4NY+y+L5GCeUoW9EvPo2qZhVQIB8DelWpKIKJ+kRPPwtlLj+L7d5SadOpHlt
HK/LdDpYGKZhD0+ioWqXeaefes6DMTXvyVNwX8mDNVjHWHvfLvnzOnmIED/0uZXNkoaGHbC6h73m
l1LRo4NIn0Zf80f8VhyeyoWn7ug2S1ncydyPzWT8sfrb+5z6eNKABucuj4qIlvkXKsiYalN+qoOb
iUo3Ir1DHuQhKAtu44yYZ3VhDXvk+EjhZ4c85oVpOqIEgrVwFKR+54tVoKjWlVgJD8vwutfhdBVf
x/YaruSc6D5u1AcC4x+TJQkf0FqmXLSNPOcAxxmXkx3nf8oyAhKMP1hUau9pSeMzKQe62O84MNc+
k+kY30MKlocAJbCpyAuQFv2C+MT75KwPAEOMvpyc5s6gUj9S/ESzvahvN4MzlwEs777S0t67lSTE
lX9GmvyooCiXDPjvEki6WaW7XZAYS6U3aFmuQUIx50eX87XcVlGu+dHQG2kdvBZLOtw9WH9HI6JU
ZZq6lc+BUd7fpFsyZHwH7mS7uLe3PiqM6EAyoivuTfn4D/qDn4seh4EmpZJF5GlDiptYNpx9IRho
15u8fP50IejoiW5j2eZtZGUPZto3SfzG3vi1CrZBYRXR5nVG6mqgtk5NkXF3mUSkyT3A5E7SK1FV
CaWK/XsFzYlWGsqeavEBBUA0m4VXDseEN6oTrj/WYmWg+fo8Fu9gd6kTIXC1+8lQJBgduQzr53FS
FQ6ouZ7pxaYlI69dIGA//slt6Pc8F+3dwseG/p7af6+y7CfNpTTSlfsqm441Mc+ibIso+nLIZHWd
0/hJjVQCcLosUEmnboNBQraTQR+BRpqvBjUGdR6DeDfdLBM5abo5hhPcU2HwxcvsCx9z71wxWA6w
Hma8sMOQmyD6EQJVkuQVwu5gZCN5LzIhOaAH2Wk1GzHnFbZaDTWS2nf4mKmB+aX9VUb2NdiDD8UU
t0xnBQXFZ3l2JeT6GZILTNy17nEbt5mR4YJu18TEf8lBdV6u2mjsZQn4vGUg5Nnr5UQ4EbjlCGK4
sZ0uz0iB8S3kJ2EreEWeEt6u9lMFNI3Aa1liDlH/0yY1mlP9oOxwCPFxPAFWKg8UJ3lITLSSkF1x
SSzjbV7ObAiY+7whl9De6C29oVJK1yhLGY3PJEE7gF3rX+aMZ70SAmeIVBwxM0YToKVdOYGfZYRW
5WcqFm91ohf6ysE6u6ljNyBPe5f1LWPpBWFrrMs2NjKe2kKRfdp6uFw3Fb3cNWceRsCqHMJdrMQY
8fJ2Fcm/MOrPzCgpPqEm/twqQgEeqbB/wid+xQ9SH6wxrXtMgQEQxbzTGn07V63VkHR3Ol9OlX06
4OOlp06kWAE7KeklCKZrcsFHWlCMFUToiedAstfozfJ/mryd9sfqZYtF2m7uMm8jXVbfGc5ND5A2
1KzfHkrCQ5k0W/l3FgbxMFAO+38poFLL/3oT5DMtok7lO6NGgn+f7lz5UeGc8UZFwMu9E8VH4xgg
4bCDjrvnKbS5EB89H9Ml3uSUI3J7g6V51Sictfo28e0KHyQsW0ULt0qlvvdG7Z0owh5HSky4L3/w
ZBcTxo7fUJMzpOBA/f5+jYOgoARxBXm8jaGfMKHUCQJLTfKU4htlaH00SBEwvU4YMvBho5CN5TaR
f0b927M+ORfE4nThZbt9Q0PYtBQMPaE0GKrR58wmtEQ14qcGFXS3zqo2ctcIbn9lCUQ+XJ9+6ZU1
cUGf2ryu/ukcmGfWhUmR2VFxg/O0zwHhTBgN5Bniilrn4kyYmDdrcS1+uLOCUzMFMnu63HY906oU
TzIj6F3R+chbpEo7i8eKwMHfpQ+pWZkaD/FtPLStXL8ltLt//ZKtPyuqoNhotTMkMbrcLHCqZdnX
/HBChA9NhnrfFdMyH28INzEswD+10EoN8j6tNYzq4vbJta7CMuF6fZVtUody32U1PihoxAZTcIpo
/eq51g7lxixzYC0U/M5K+YRJfg+tWo5Pl6dAABfZaiwj+SXxLe8Nha6OIMtoTlyheOcCjebgdOCk
39UY+ZOz7k9beySgLgHL9YHjKh801AsTzXNm5exln4yqIPtFnzNJ+coqtJux3nknr5TKYWIIJMV5
6QL5TEMDWtl0WoClSqRSiki3IktZGHcdFuW39m+6xEZswtRnhQoFMH18+I78gUFzK2na99dPSKHt
AKiUfO0P0gnX6TE7X6binPeBeZ/+2S20fMTaKwTk2kjTn/Sc1DAMZfgLS8bsTg8n0tMHgrVG+WOG
miMsEnSO3ULUoV1Llo2O2QUfPub2NBLsoPPGlnYopYedjah3pOQuanf7zzcq2ZWGp+iWNNJlDOvY
Nyg8wzY6XmTgQDiOvIvTMd02tU/DYKOpSomk541yeDmc3EYpAWdkBOLaxv59Lq8CoJHJIlaPXC5p
hrYvWnU0NLWHMY5s795Rl2aGMoQEYjd7yyQaAYDyNzNXSJKaSKnOHBwxBnyU1+aznD2DC4JSmBsv
FU+JFk4sOQdt12b02MEpp35GT9Z9oHmvxe27WXeR78I5M297/CsNCIZbvQ1LmVgiwyPTeOU8kC30
tFoPQIUbFWdsNLTF3v+gKntrDb5vEZZZX6JnmcjfWXvRr/sayrsU0ml/u5LI1hDC6m8jP0+AmeJz
3loWE5vheXKWMYE9jGGbvK24g5/ArYZlaq/cHlYCHnFchyaEj+KwANRq6PiA26EkmOUlNc5s8LS0
m2QDbdWxG01CBoP6h2my3u5zb7ZtCzHNmqAM25XwADb+hljYjns0B1j1hWzNt64jT1NNwmLcUx4t
rr4Mgg4wjwvrnnOmZ5d+x0GNdJytqUaht7/Q9QdMuz7pg69GK7JqtbsmFEZVoIOMoIrZVPS1knNJ
flK4JNHWFAH6L+Y33Xpwosq9Gl9SGHqDbBZzZ5RspXcxgY2oZAU16MxwY2GidRK2RQQtVETpQdGB
yZnj+JkO3B+ndeVvuW1UKp6Ew1VU1jlv0NZAOf/KIVJ32WVCx38rMHZ/+RuP9Tt0JDX9+scyeZe0
wgW5pZGunNwtmiOZRupuFfEtWfxfFjBk4vSbZuLbzEN7V9hXsvdL5yNGHFxtUBnPg0QLroe959Ke
jQGBKtr9N5wTcJOJz/VQDwOl9ANfeYNTsKqqXbJYdA/KTgSN26Ja7fKvbNcUU7Aae344j97+sFHx
wnVLmXKAFyz1TD5Luo+FJftUd2brcwENyttX8J73bQKvG86bz+lzFHUyd4vJU4+wRnxpm45/WsN3
uJtR3dNPDtdRjZlSlTdZelcsSO6r0LBY1ANf+W3WM3wp7ZTEO7m+l8lkoy1n243UIdrfhSCsJLVV
YhcwIV836FXhp0n0VWUDJWCVD49L0F4z/g2XVpm5GodtxI9AkWPqXBwiMMLSygZxYudprdxw7wTH
xeCssvaFPBIBxHOddBJtAUVxym2HdmEE28M72Pvw+XC6B9Xh9CHp6ZVPmoOeNO0vzFLdksM1ydpL
qExk9lq2tM28dWfeTyGqZDx56etJIhgBslTnwmgCenG/P+zsKUop+kKITDxnlS2cwuG8tKNTf6Ax
PxPzRDVllvch9o4Lh0b8cT1pbLw4/wYFyF040hr8MyDn8PgCB2Dnw1F0dmPKevk8gaos9OjT1ZMM
H60fBfQQVXm7Hgq7b9DTkVn1RJvRz0XVoyIkJ9EdTs2QgmS+OPonKnKh8mnE3z9IQmsjuopmiFTg
BoPYOjjL08kZJdMlXlhs1SilOrx9aVFe6mRLH8fSBZCLBcjFAMKBgX++SioYJkSg62NkEj8Zx6Bm
Q9pd9opRFBirCRSDzkwEmEBrdyn6RvhrLU8hvEysY2TPmgIwRNSrU0ZpXAvWmwZgBorj5HCgRLP8
i4mY7Bbfh5TwWbZvFX+HcbFd37CydrjtLx6kLhWTHY2sQKIMUil5QW5wLTF3eeD3nWda/puhxlPT
fvF/olg1HQGUi18zH0+8U/kslsWuBQ6qy2kxXWkjhLjp71wmCHP7kUDszXiWEP8JAcKjvCJAxMMN
YdQ0j5gEQKv2HuQjAyBvvrBtdAsFl44HsoMhNTK4IjcnV4qX0tWHWDQuBuaftCtWKo1j8AiXo3ys
sFSjSPdRis6pUKTCBhsnMrUDP93V50K3qe5cQ2AD92Mb1JP7IhIMtdjX7lrZVdxr0LEI2pOmc+ml
1rzQ4+cB/MhLPPGZBAY8iLq3v8uIECZVgOJP/g9yc52d/LLlG8YvVVu/CspWMXOuFX83Vto9PpPu
XZWkxgUHoh4K03TnLIE6p9RyXSBBP91vRTcAFjOYbeYMMK861bV2F/p6wc/OafRkxJhBuxoR0KUV
3JqGK+6w3aL4DKzjIBFuvG8OXUlhrcbnJZPenyphcfGY0eFsN5VyCb0jdYZK2wG2RFzS7vBr4y+S
nNgjxFtCj2ZeFxrjNmkgTJP2IkTfdxf3A1oUASXJMG+X/I7VvtYbrzI8q56OKWfjXfjYgVOMn2Bh
ABFbX0Mh4xXaQMowXIXZBwrvXmoJZmvLdj9r1pI6btapWeJXF8T1Qz88RoUDSW59XCxVRMeHnggm
owpnb8rYExZvyk1NCuFePYqA615/EbLlzx8T1sRkVBGnYAhmuW+2fAchQ4lVCMDMObL1+djQM9s1
lalE4Ta5ARWgPZLsozxwUS2VEH70aBdp2+m6Dk8PehqeHt1tVYjTc3+tVVtXXsFBqvUp9Rfg8/74
vbceTHtk6Rnvf6oPl0gRPc8D447vNDxdwNc2VrUE5MFBPpHdIR+Bedc4EmVb7oMemutYq4Bd5NgB
6IIGyHS7nf3WUyD5jyXbMWReQW31KHXk4U/h6PyMftdLVWYp9qqppWARZYNe9wGp96RlOLro73BD
VPBp6hADI3/DlklT38zU0N4Y5IDCPH9O6OTtaTIo7zirIWLdAZqxUSrkr8JlALBEycSsvORh7/X9
JM6+kJZTc/ySlsxqWKK69YflTwreTvrx/BbJYuguc/CP0mROauQqEdLN7BiuyHDTMF41PtKDjGbE
gQtDxSsJzQcH35jHcMfL2UhAgtgM9PtR28ynZdWDZbk2H7U6zTPe+kviYXnW5EICXl8yg6SKaIhx
T0mdIdEmGHTj6pdm0yku++F0+7BtinIx4CYuxlLr0UmojiBKfEGlK74dANshC7yEynqrbLTSzVnp
wtKO9gOv3ugG75AYfE+imJH1dfzXEegPthiMom64ppQ72Vx0+lUMRsvZrFErBnbS/roz8OJTMAav
+bKMr/g51BZBvdggsLNk4CDmtss7y4fBn4wLYHyy0upZw9Xn8Dw/ktqAkDLBw9+3cPAvq9XL9saE
/UEFMKEx3PixGwh2Une25jas+Fejom/dU4oqkbzbUevShYtLlk89ivFRga1Ef/da66qTuEYRetSW
tDhTzhOUyxT3V6jkUArxJWCeZGx/r1F9QPW7XtWxNSwi7p2SuBkkw3jtAGEEJR8ANSNKxgjesr51
7wNAbZIaH1zCj3G10ix1z2CBNd5YCPOs5UIaNdsOEMikQYa/o5xRJtW7ZOW6Gws0h9S2ryxZ6UEn
VAikY9AAFNDDvD2HvLGptdLLQDWiTQX8eoWbmIoa1ITyVzr/VtzeHjbVz5V4Hei/tkj11hoEsj70
XDDg+xsUumY4hRVwURZjCrZZ+bQfPnpeFPuR/1mROoo0iFqo2V2/UUFtkQdxxseZCpBkt05uq0HR
DftjhNz+vtdFZa6pg4fAd9D2NlyN+891MvBTbBmfqP9QBy4hpuFGy5RSOEPcpOEzdxO72JvjBIKO
ILGPG8TVtHFjcL+4U5taa8BlyMqHUacSn3LX0ka74uioi56Kuz/UR81lnNT3405KQMxVlCN3NGaS
w9/0cE6KBYCzoKIpLj+6pyNJ6v8mCXzIeLy81IsGgtLLO0BcaK5pA1EVEcP+XDKokxDkkNLck2o+
F7Xvd/MPbKhd2oZ2MgGfvd/vXcBgGMSkUNezO5RHbCZLvcVD/Vq9vTqu9kGYC7WF/cHORoc8G3dj
bkRf1Ma8iFkpK6vgRIbfWpNxT1hBKFN+CIZ3dK+ChWfRVDqlIQLe1HQbqby/x8GF9HD9+1YHmMrG
iurDyxg+ohhY8czZqSSvJKA5YqqJ6YagRfULsSaPDAE1fMvxB4gG5kitm82gaQzJMq5DXIGg25BZ
R9bQoidyHrlvvVlIw2hPCL5zkD2LOHED4uwS/rt6PrA7SScuax526aAXjwQZQ7hsDAoN6xFyP2Rq
8/ESiEFUddnQSEUKvAVLRXIONPqglJcfHuzYxuN3j7Xb3I8+X8a7+1VvJXDM6cMBJyjZAP4872E9
RrIhAH97eyJ4ODT0IEMU5mC3BlnUiw9CVuIsDZvvpv63/dzl2ud0IQMDAxtndVlNVt4NqJfokCX5
1udoUKm3b2i1Z/WMnDLJ3rji2YcYfapcOHE4DAD1r1tU4oZwg2rfMIl1mMgS1GWT0wzQpHQjRnBM
KHv/HekgFZBWW0go2TfxTYZ5Wydq+nme4R7LqLqQ0PiwRke3BAWlxvPE+9Zp4KJ4uq1bA3e3cEZh
5hTepsfzcv8MYCAE2SrThYiu7ejXIjeF3FFRvl72X+atDegm3WPIqP9EpFzyLKlucqlkQWh4mDw6
qk2fBU1BWJe8WAQtq+OHN9Kq3wHWokQ8RuLECFrldLMVIYniHn9GZ5YnpJybR8R4my35K9hc4x9Q
Ql9/JoMG2s8nc0Z+UK6fAK3O8KV6pAvN84+iIoR01k4T+7fP2BXOMAONXJckL9Z4048UBKNAe/y2
x0s/2EUAZSBWl6iY3tzCrjMWSoHhTu9zpfHclTPd5JTHJ5iDGq+t8hhUo4kXLRrhJsG750p3AlEC
HOkRkOV0G9f/0xHer65BNvxUqmFsFOUAXqlYIaN+6PBCxrDU5+ut4kRDLLkE498kL7lYOjGj4lbd
eanO+me5BQ8Oif7ljcsGejCad/t4JKe/Ek+PkPeA1CY7nEMzKULjvB6gPHgj3FXu5zsT0haR4fTL
PfLEDrEeYwenRF8f1xq3QToH0+bP2pwIfuYDMtnOQHaKICxWtHDZm6VFlMWbpwDxXDgQvYuQgttZ
Z9rmAg+RTI3wuC6TXWjlV6WthPf2Kwz03p9pijQVDyxh6PBSuL4lnJI+ztxLd27zOS9juSxdKydc
YWTexWtX2iFhfG+MSLBWJTgXiI2f3inH3LTR05LdIq0zCspktxzC7mfiBodRTKnJ+nKa1q9eKfPt
1KLktOfnGhdA7TMQvjdjvQ9yYCzA9nliKRuA7A/xGo+qUfF/71kvvhLBz7yTOD0kZW4JZjtcMEDy
Gg4opaKYl7yL4cv9Njxi2X5wBpu9MHGhCc6AodSsNkShY1eOQc8s03sAh8LbRlx/EVW66uLNWBVY
0iFVOTRIr25zlgp806Oc0RR+lry6ivGPlCMJbVf9y61/82eJwVX6leYlvk/6hvoL6tZ9UiT/hCfR
j+uLCncaoKI6HU8GKDGXHCuqvq43YTaJjq6VyJNqFMmP2x0PHQEd63G/blbKdZ8EhVi5hF+PKDdN
yIwsk4R8QSawIsTDuf8/6k4VMC1es4JoXtvnRKTTtCmITJmqU9Lw/cjB77qzk07YviuV5Z8QLZh5
EWM5iEve/uiRbrIUXbyyEVe8ygEijKpFFJggjlgV7b0SRVy+0Ml/gd1nGYUZTWj5RB64M+4A2gCI
dZZiz2wUcV7Xn/VwJ4hinuN8myBBV8D1kMotX64PCUq/ROnW+OJJGajsMf+Mtha53zeGhsgODNAf
k0iKUxCcVTpBBrvlFQovUkicCUq+5j7/LMxnglFBPRqlmb1sN5wQL55ajwmLmUJGjP2tbadbhvmu
LgZoEIyY0JFiL20+6lCjA7wOgI7ye3RJUuAZvEzPlrIKaR33npvpspe/W94Uu5hFD1mgoaft1nHT
lzsm8u4kXWdKsjgHGkXqbWGe4u8Ek4WRA2hloLhKEqu7lrbwW98d9v0641G9ZZ8d3EVRZSbeJlhH
rXXnNhPDOMAoyyWcXid7m8D7Cbc8Hst4hozGhDbS0sM2b1bCjO9FUVbKCbiPtwny5T/kk3GySDwJ
Z+xM20VlM1hGXN7jB/D9F/07QQvKunmBc7SvQUHFQw5AKduEcN3DllAKpSOCh3tyt0Au14AaKT6C
pPZ5D35AsL/Sm7nBJZ11uGUk2ip4CxCTJpJI6NwTJODmIvf0eAgLmsXT4yyLzAFrXHcbmMDpF4rX
dfYg6QcL6IrPAxn9vPcnuvT5+FmxNiISiwyve2zrxh4W9pPRPqICEXY3u2dDDi1QYBgTN/z73qs0
lIfAnTlyF5uX0jxDMYjmAcWurTxluMyqB91JObjxJpKxBOJuFB5KW7SGyh5cj3PjsK6gCRoLrk2b
A1m+UFVtnYlW5rh0210ds/99bKtWsa+XNL2o1lFuJft8yiSDidmzP3u0U5qFg7tp+uy8UHeG2+WM
RB+lvIIgMY7xZGs5BCu0kb2gytbpqo2VTKWW5Ip1OD0cSYRTFdgYTg2Tu2vn1GOipyifYTzii5Tq
QIjmRzc1FDhpv0Op3yvFLWuXIIyiQU1aXBJluj328yg0rn9iWgqgMmycInKR2lJwuEsDXkehS5Wn
dx8EVBN7V0EnOorbNub2+IscQ4B0y7sMkAZAwubwDc0lTnj1QXX9oldEt0Xi6x+PaP0v68Vg1IIz
YGlx5G9xLjVw0B20DjabbPCHXxumSAS/mpj4wGW1iE/jhHKts+VndG3dQlPVo/p62+8Zauj51IAj
h3RB7r7bCVqxTmg7mZHq/eI3UvPCRUlme4Y00yGc8gbG5daKaonygIuvmVNDcGyqnClOP61oa9c/
IZAfUOOihzOYGYhm0rLapFMuezj6RovXQpMQlDu0M8RmVURmiXK/WZ4/Z+bhx1iYQbpsBFyvbiDK
/ET+Uc8tRVMfVq8ncz+GBltCUoxQQr20l879cbAL8sifqOdTlVDCxf64G8dcl2PH9osFfO0S/9DJ
rai7EUdntU52JT6w9esEXn8cARGL7cGdbEp6Cv0kTEP7b9XcVyBIF/20AjfdS/SEtkiale40Qh2j
thWZIBG/hVe6xEbwrB3m54oJmri8SPaH1PPpbqgdYa8D/j7DlXOzqEjdmLWkgA57dadKjgJ5knXx
OtwoBTvT3c0mLtgqjz+OV4Kmp7TQLF95YOye/CnCxSqYQX7zd6dMVl3rZtJGvK5pnc5lTfBce8SO
SyOKgYfFCO5Y09PLjYHwGEn9sm+zeNr9iwF832nvAScwZrPfDQXljStcRNpC1t8pK0YoN2D29V0E
EHPZ1e5Xs61gj58K26ubZh8mHtM4uHK+pOqBbLVQyHEd+odwo5nVdynNFi1XlmXMFvL+NvioaAyI
6jqGnRxC69JQexytr+xMhreM7CNxlZfYawZdNHZeklcP48kXRfcDqAEEl7Qv3y7kZISL7O5vSIZX
aSf9X7nM8NB/fzd3ZF792iHDkH4JtchWPi9m1TVGWZW1dDO4kjwm6Uzr2lcRKJ+yyEX8gHFPE3RE
vNspcBF+IZplWqktjT5amvVBAd6OOKF5/XSfr37zXwzqGpz54TpBA5eEd+rQ8JnHHuDtS1zFyqxt
2PqYIvZysi0GGHLEFN8TcBToo78e4QJoL1TbFuWFPjeGvZpP4iZh/tlqR2UEpWJtfoKArcVwiicH
fx3pCO855W/LI6jo4Zas8nmew0mHzWxWBYrEqjX/Gpcjt42jaXYk9zSMJo6K/bbovFGZUjICpN6U
Q0LbuBRnBsnP5OZz4IonkkdW48YM9LCRwkXmLgAWAq3D5A0f5FpOhk7qn4ShsF1w7kf9ZfeNCrnj
RL9r6QMSxUiBfA6jn6mPAQDlUD6ZWgl6+M9ph2rhCwsgomMBJPk3vCy32pxd8halnY/RL2DdCSed
agKl2fzNE6EBQAPRWiRAqmpoxN4amS6EhrNL9KDUA6PRzBKx9MCLgxvjSC6rBoASEnxvqGS+rr+d
eIOaIYpekmhWxhXo1fuAZhFQOuw8ZeF2z75tUKXmN3bnKu8h1VnBfM/OLNufzj3xan/8H0k4JzsL
gk4B4pJIVaNwktAd1KGQf1HLkGJK26jTNOSLBTVQ++pHb7qf8U3I8XXUzLlmXnMtZwRd57zfGQbB
Zw+PMc4QgU6oo/MGXfBQG5TXWSACS+80wyhxMAzH6W8fNCPHDnDCyC8KeCT/DYsqTx99pcLFm7vs
sADK6QylKu6WqyY9cinwza3LrLFcecb3DCK1cTU2ZVM8xbUSM9R9VppUcVOAYXWHFGyTQONwMNMD
7UJS+j9o6LQBWmlyo/SsGp0lKeMPqruMdeBDoOelnUdoJ4d7gnEmCUjex9qd6zHMFdKRYss8Akm5
B9iHQcggLNaaItbjgoZ+OP4xxa/BdxLbCVTKQQv6wj/aYV9Qjr5E0FVTrtsLf7GM2vuCglEetgHB
qL9m3JqZ9iykfDKlVTMNax8z2zWWLRZIitH8aIFbsmGwKzEGaRlE8WZGJs64j3yNwcTFNfWI6+F4
TCa3c7sj9Gr8zD+XYl+pc4Uj5NcimoYC0Mc8y2AQC6rSTOsvWJ0E+sqK8n6cxekM0YWw+gNi3wOc
K4ch58MGcVGppun+XWwKbmY1lktiwni+fGgdM4rdPYiWqnG3sQmmtpyZu/4+7k9YY7pEY6To241z
57ep+m/fRLVbfgJCXDNNGYm2JRXiobDHEX4ZZYmJOC/VifeAjMNGvCeLE6YfMDgkGv0+lfEWPVW1
9VeUFZol9ZH2W8cL+NHlKKefJrjg6uPExbmux4J1ZgOuE4FwxDBci2PBRjvwTg247jKbzUyTzIau
k7JKLXJKwzgFDEoczc5NUvUcVG48Bzc2BDx0FhJyce49nyFUGF8xO6sls8cWSc3wj9Ke1uberNno
WHxyPu78xuyG2DWNZnFZuyBJzDqmJw2NVvEsFTJ0/C+CT1DXPiZuBBmXP2yMkgpue8VQaqGp29+o
jTPWk+zb3FCMBlRWvYBRlJGesWH5U+L6Id24WpwYkYMdvBZ1a+iAF/FvZl61gOLg274Zup7uPxLO
Dy6pit1Mi0MaClFcE6ydvy/PJQ30OQLDEHRteHtPtLp0/AFRmNHqLNaJkrOEeeDz9XSimtqI59ip
A4Wtm0ePNotoF/HWISFVCM+lcXDYY5cZp4dIGjWsrafnOaTcwKUCNPkIgx1/m43H250A7P6dJ3+a
5clGMBI8WAgPLvGzVCDW1MHhtuljhQ2HxLjC55hca4PA+Uy7T2AZItVWBMU9dyADCjQQmfxFZUQz
Pj2FoKA+Y5RvPBAotKqoEC01tdywVcXfpQRn+F+TZDClXwLJY0y+6k7YqZCiDWsNYrcPe/bceZeB
Hb9FE0rXGlYbH4hTCiYcJLUO3tf/0/Iyx0inzwUOsu+u3B3ogzLYWpBKkmIkUqc4dptxWMFfNLpD
3sdihchUYe+gQiWbrLqkgcjGpekX5a8x6TuHgn9C7Uax3V79iXG8tQU+d0/q8IMM6vJo0lqwcko/
4eqNE4IQLsECSbNnFMMDnkN4+/7fA5sv0RHTXkOQ7nk00yY6PKCr5EKL8Wnyly7O8RgtAaIWUA5Q
Aesx6ttryzzyLv3kSYS4dLtnkaOCTHY1qDecSWtPetOkjXhhdjRhC3yV9JD+klU5QtEwZABTDptu
W9k11nLBQXTWRlJPeDdYvpf50chKzqaDMXx9nOpqfvp9u+Qr3DY16xH97XlVK9YTDIToeerZBE/C
AX1d+t2MOLci9wg3AF2oM3udN/8JOZDzOHgtOUuvNct//GMGixVKye6bBh2pF7KfXJH5zacH1LFZ
u8Zo3qCTNhJjSYSTQzbn5h27wM5vu8//+IAqtmCgqOzbnoq3LV8e5qwIRwMy2CJGVZkD4Ye85zlx
MaFmd8GbHkJHXsFNjnZKMovHAjo+16pqaQqHSnFj+yXZj4eMfrknt06j1zU+YonLhyw5NnbljcW0
0xhzALDUpDWIWaiB7zKI8j6VZkumkn2BDnidnhzjSINPqznA7Py87jdWLh44TDAwBk+AidVhi0Rj
734tPHY+ApXluy34GTo+0vo4to0mJvwENh4wNmIZa42P8hfpHVxBQEvgTW8yUArte8lVftvBnXg8
ZieMY14TuNcbFoGE+LhfKBICHVOmPePkO9i0s8Ca3DiN/v3I/sNYbMmQ7QrbJLR5zjURtoqQMEJa
RThuot7XNTK0n3/vbL7sE7kYL6uV9ZUphCmABtGWdVeWkYbo709yAJllQCmzNdq/CoJEZYkzsRbv
tPt6qiKssV+ju57XSQP02rraebK465REmqiqFVblHpXntGPYcbs791PJa8Y6ZVH5kgNXHpl8VpVd
w41k5NPUDLHLmN4ULpm5sAu61ixqQWItxw6P0AvkXRdo2hzjqvYLnwRCQZGJdqCiQvpWPpeicPHe
Qsh2xDfam6MoEsP6+0fKU/TYFJH+8XpyZfLN/yU2sQv1//J9iQ372PIQxD8Q8IUNxDyfZZXaq7pq
NEw9u/dYQYoqdKIz44QoGmwxR3KKfb4H+SVu+J74RGvaliJZFg85c1tb2y5umw8QbOULPnvL5ouC
jj72D+aWZI1ngY2iqYyopW/WTpvqDVu3xwpywjOOfG7/eBci8vh+ZoNcPFhII5YGTh61Cco4QR7z
gCtW/Q2hOMnOmDI0hXttMUi/BLN4mxEEQnDK6gq1Fi1wqyzsKcVx0EokuRf2eZ6U5k8RTzSXVK2H
94S6rhtRzd6ezZDoyvZ1nc8ggs9slJbQIm5hRJJ/mxIcJzP3GFRwjHCynIGiFE4eixkihrQWDtbI
+iZ1COQb+mCbzr1Kzh/vihm5YHUCqE6qdg3TQBr7r3SdLBhBHsJqNMzx8e+9smiVroRWupESzxUq
qkTY7dPUP8Y3Uqsl27Hg8NeqoVJReCBOexhTack14Skt8jaRZ9b8KbAoPuIbSrhGZkAowLA5FBeh
l+AbdKwVXadr3KDc+3aKfRTYmq/MtYksnks/5aaIaHXZYFzlfG3hJTIxWp/iug66VFTz9qqcZv/V
/YR1zP8p5lYtQX5hBur3ln+Hu/MIgfRR1KVwu3ooEomBUIXhGXTvXltwtOQVUvIG+M1FFrZskRes
Znzu3i74QGXTuHbpCl4rD+VsU384SOOJpee9pzOvoeJl3gejQcJF1shxkglKUMNsuTYoe4FN72aO
D7p4SHOmtYUOtZbx+fk4AdF3/GDofg3+cCWzUWs8mvnejBc6CiR+N7uXnGcFTKv48pkVFHd7+tt6
ShXw2PS9V04RL5wG5ewhzl+sGi0lyp+Dgamlz15MCGLbDbQSADnrl9e+PXT6NkACZf8J5wjsEBCp
R1+BUyH0fCSqHZ+dROF6bUBmKzUkFEQeCAa/rhGdMybxh6Rp1xw3p+hGUySgYUrtH9IXbHLWhCg+
kKhyxk2o8W8JEBBnd0D4mZ/iq/9LoE1fDIBZpCD+tXiiHFZoeYjwREAIkFsjRlnRJAaXYNV++8iL
9A9yjiV7kKVLqGmTJZZgjKMvwhVLtP/E+uyc9yXz+PAF2KTwlmmCZX7oprztRzdjby7xYjwv6r5s
Vs6O95gr4Gd3GaudAgvWstvpszcY9q8tVhkdbDDf9fDcbiA3KhyqQrMIKj2GluWyf3QCvdPLZeWt
aWaYzXrmImidiCrE1D2nKj4XMS5FWnzPy2YFl4t17XKDGzo38nLk1sbZUDsKevrgpqFRQa1gYUrZ
p515m8xhebtwijA6dsdnsgksyzURF26tqa3dMC1Nr2Ev4/YPuGhrxtpT4ZioSilvsSU+JM4ePdt4
zNgsKLZpWi1eSpxyr2Ua2EZWwgvhBqjzFhlU4iESawsnwpK0Tug+WYaEmfuBQUYejzuRuTeloM61
oCbaOl2J01L4DYN/QUSji1e33CUpMS+ZjjYAErWedlSyczaP3gjjyrS+2orPqtYdA+7ztItLjuN1
3mnXjYyibSVsF7sHu6mv8EQ4KsmAvvnIrXdMqN+0CeNp1nAFid4RvIr4VoISY9G+InD93nbuet7n
CDWGQlqjxcmCa9zhRR4wVvA4dNlt4yfw1XfLWuEoLbD/s1gXb9Qf7qj9886eWQa5WPd/oJHinjzu
gOcAcCcP0r3gTD2Gq9WAYzaF5k2dMMWP6CHV89kZWIc8NuuId1v1THECesWOea+alBaHeRxs1SNc
YiAIL2RXKEfdi+yZOezcLky8ZUHdihdCFJojqThxsBM+2ZggoESNqXnTvunUe88+oblIBCA4mbGL
U19h3D/VUactewF1HKkKv7wBziq00BnJEZGgcL9ye/WMTIFkG+LkWpyTIlq8JVYrXVJLj+j94u2v
KrEk3z5nfRPAV7OGy6bHdQbfaVfDldVp/XutWCXpaJzHYZnOcqZOYu5gmQEtHxWjyrP7obOmJ82v
6ONQJJLYBHGDWtrAUPjzM8N5XV8IiW1HEJM3GK8QHdfoDtUflEYxrF0YKLYTVCEEgeV0QPC/6zWz
2QsAZvWV84A9lVFA2oRq83pgCXHlmRqIhcwRHj52LhBnAUHD/j+Q4OfnWc+K6hfDlZJ1XRahME9r
zTPa9iQY59HQGg90iLFcO0KlqNy2nOnTZTq2wc/H/XUcpf0+8CVZgl4a+SYCjks6jIBKn207RTRf
M4Pck+t7xUE0h8aczpsIVCj+7zKeQD++0l5IKchRsHd7GbEPVCPN+Gwk++bnl3o9eELM2s/luQEL
AzNt0QIdC51Xel5zIWfaXms8oE3Q+EGa2lW3oQ2jMHOGO2R6iOitZxsmioc2QmVw7T4tPJu7+icS
tU0vHwahO6o+cUrcYEV9ULnDFwheD3q6RgDt/S4pV8nm//oS8D66dXpTQ4oQ+utk3vi+DweFud/C
XXaht5SO0jbSv5kLsRQEzKB4EmHI1DKpgxDxLlWbFmTQtK6/yxCaw2EDgpdbQB0/zVLc1YayBIy7
bhIAXXjolypiGL3QYp8jFJkq+NKd3hgloPXjFFZrE0LT7p11rY+1kgagpGNhx1buTOez/4/ORBm7
QUz+RtYocInNsG6xHrQSPaHxUOKDUGcojW1slXL4p6Xj9P7KRk7TlpJcbBFNXGnarmOXJ2mtzrXt
cRW7s5SA1j0w2AGBcpK7gOnK/6o2mfSQo/ehOnKQDTnpIVQ1NXWhJ35mivoOFsZMHjv3MdeN+DAW
iMn6RjHOy+/QziDF5oarOUFs8fP56IBKiiB7mvC8oW2VipJ7fHN3kxlUlYIg/C7TgeOuQVzlg0y3
vr7K0ic0pBNs7ZuDbXkgyP6J//kX7UQf41qTLP/oS2ALh2Cdh8gtNafcchFW2/UNl5QdHRU96nNa
/IEimk4bvGAJ0q/+FHpeqUAEz6YgUn8om32UagUubXq03yJd6d0k3XSb2jTciUdDl8px32jaocvq
5i3eZDgCVFfEMm/9f/v0NQh6wo7W64BgGiDkCEPk/G+inHwWRRw7QxNv9Irto6PlljbpGGooGEY7
HViiL4waw61MTCS60CIZ2q6//HhlNjttqMZgt3O+O1OND0cvNOXM+e8KQrpQ6ZlE/YG8IicGQSyx
xLvGNFNbf+PAIzwg9pDGmT3qCIM+DbhIH+YiStyeTe2qRgpmDyMjb08sLpvonFoyU30Btus15Qb4
5iU3qCd6hAGimNnpSqKx5GUR9Htr8ZI+X4bIBh+c2m1gdyYXz1p5tUWvUUEUOSN1p0KH+nhzKEqv
tnMAsuxCjchXwweXhMmsKFUh5gnZ3ZkRcSViImM3Fd3nEy/yFxpjxztdtv2KgEl+bPwHbT0ihgUN
X7G9pa7pWKgFJhq44eArSASiEy2ylnlEwEW4Z20fyKyart4ynW5XA77+dOlchCBFMJCGYBHh6ki/
B8q1HoJAZAhORE6tdBbfpKX2VeP/h9b4gNyWzTuWgVZDL5koDJF5NrJdAtakaCRzJ+B08gXT3wsK
vBxmbEOXEM0plDMKlbN0e4Hmv6NfxgAlDwDgdhJtGzQWmRkbp2d7aQesZRzagQW6RKBTY1rm3ux5
p6pDT5+7HQEscUVlq81dCk6ICjjiTougEYEPa/dEq7wn1ORhjQQlVdPwf08W3dbP1XS93VK1U2eV
EaI1Xe3NjHsmj+cKPY18sSnQRU7dSUXvKiBx3R0RgyPwmVQxO81rVSkH2BM1r9skMaqrjy5G8OHB
jnEArfd6DJ681XZwlBY4mYqpKl5+w4KwI15TXdyANXwn8xvsdTxCJSwz9IOKsX8Cwhp2aVRWUvW5
zJmPTwOTPV516G8ow/JB4ctFOJgI/q9mn7KxP0uM4jCvIlR6Z83a0Q6xG5NdYa6hket9IS92WBrT
WN2qSdDVsQh8h8h+KSaShJpS7yIJH5JiNtwoh61KAGHo5ziZk/6tny3aAXgsAximkMqxouV6nYu8
w6CYPdMhrIkDe/YpWr3+AwqAzfj5sx1QkWhvhexzPkUlO0kpwvukViWjvtnAHId8C7WtINdBzpNH
RpH2B1hpZvR0ClbiTmFivuvKv2BHY1FTgVebvh64LAcrQ/IsbEK2azr/MjFsIHPQroxg/EhrV8CB
n6lmRKe14bH3l2ptcuYkvcGqhb9CiVOeID+NMlaLpryfzsxD8ZJ/YnEz27IxkNnLew0FUI+j6pMD
He9L58BYK8s/LFOyoGm/pRY4oYik/3E8X9lGlXKVY5+YK8jAr1KLS0OLLOoMaw4i8T3T0WQ/2u4z
oE64o1ahWLsHUGYnz3Fhv6O9+OVsipAY37Sw365xzH8NjbWlORIahnwxe6iQNw1mHQHiyFbTfCOO
b7DTJTfByNhC9Z2TwiWfjgSim8PW3h1l8e0lFMQqfwQBuPOE/PeDc0nwgjL/KJuRxsBZdf8aHrDd
3TaclCqWPmfwaEfiKkm+2767NkN/dA9lfxoryqJSIAzjCDLCIxK40SV4xRi/ev0hZ0dWPqayOHHp
JmMW/HNYq0IGTnTKGvYhciUthkcqWQ7qt2ABbomKQ7QcE5ShFAtKwrAbEUVqdx2qhDAaqtmOAOiz
heMjr1g/1hvOntY6driDJtTwrfoxCEhygs3LVbBIQQoXeF002qQiaxgfuHv50YvmjmTYn+eX/wu3
bPy9JOmIeXtZcSA6MXk9IKalhRtHw5hNzpVYig2uTYuacgBaOO4ethrcqu/1JazXJL82KTCwoH8P
r77mdWRXiC80YWcIZpkD7VPzCY0HPybnyMiRQDEPTVwJceKyGBl/iOiKf6P0RMIWpcwafWOtDOv7
tj+URgI4QUf+BfeTCg40HwdNBk92ACP1vnUItEz9uUf0srvEOjR3Yb9Z4YttB4sl1CoVgA+8Gsi/
kZKvD55zynwqRxsypOImBxxkE34xWDJM2md8Irnze65AYtlqQX/mIbggsISvdoS1WDPq5usf6XgC
zFfEQu3+8j5Il/T4vKxLlgWHvt0aKgiA3fH/LiXaBaUINvfqIQ/+1EgDBUfgcNSvwCChKOtwWrhl
WlmEndd7oS8oUvDtpY/re0kpfP3vSV+6+xsardO8XnbbgUMBD/nhxABJaF+m6HHioVOGM+p+hf1c
erjL4Rba7iat27VEdj7CAbhzAhlXeXlWjiUArNMP+hl1RSonM65W8Fg8Oxp4SwlVRzBNlvzcmTs2
n5eVe/YOUYrGTcmPYrk8YbhWjUuivyD64qVsOtQhJW5PbpywkjexsBIkXCZ8UoeDnrMtSrc/aIUt
2gdwoVbPn1m+f1yjrerRZgVOOLGEFg9kibfkDBoBRcniJUIiCTOvcxTeG2OMfiaOdhRAh/zDfgZg
5QTX9S94rr9yTGZNlDuAFkEosj9sGVCac8d0u+/SYcOGb9OtrX2zCxqZ4c0GaSnTuH7WMDzx9DhU
7r4Ht7wciHBGebUgYLAeGs8CEs5gw7o/tWFa5GDVa5bEJgn58w8JnPye1e6eoBsimAqvG15im3hc
PH0NG4Rianv2VCXyG+to5x4BJy+LbJCcxFIdZx9pnwdeLGXWxtkyx+kkAs9S+ASztD93m09RPQlE
DfZSau4Za+w6bTVa+w1JZXjuBpNIkvuhqulbjKuOp2AoMaSlR/PTpokIzbPWQdbNP8jOtPEFuwYS
p24RP5am04chQc8M5gG/FD1FXoytskO8fxsGxL9LpXjKjDuwytePRf9ZWYqvumDQXb79NxGsc9V6
ZEsld3LHVIXHKU9oYvHldCumsfCWRNEX7DHQbzy7XLrR7+fxyX/O7EIW6CnnpYjqxL6vCJIOy8VK
DcOM7O8uYWmdSRqBcCTQoTluD6h6hDeqA+R2FuEoneR9buGJgPpubcni+hHFOwL5KzRNKtCgh0vl
1X9ioF6v1KwBCKhawxZs55v59ZSTwLrjhRmLyuy9Dn5E5mpr5PK9BCNp1zJBfZ5AgkEzGp7fVvf/
BfoXRhPIdqtj6vcHp20NDSm3nI1JkRiSkW306NfqWUqaVJRWERsyZJrfSAJ5Xc19D/fk2Yqkh/9N
gGKMoLmf884fQ8ch8EJI1IPEOB8thg4ecgkYz1jOQje2daRhpe4nNS+4bdzQeatFRupwj7iZYFHn
/aMmsES1mmCv9jr6gfaaRlKaZIKERBsxSDVVLJdbmUHNpqFcxgDaUt35Lw5h/WNCeu7MvVgeeSrw
QAMT08yMVOs8NtQ1bGq6FX4Spv1bvtv0al/CNKT3aFobu6fqaRGO/uWkJDJvkQUF8eUeZa5tDlXD
CGQe3rnnhurqAyOaqP/MWwGT5yB9EBfLeKWWetZdYXiDGQqncnljLTorqB74MFw55XLYb2HUQ/WU
ENuvhnZtonQDzSTauTH8VMvZ2T78wt9z/mGYEoLzEfd3RfeN4Iieho0XpMxBKPOn/8758sw+i/0m
UIrugQwPOyNJIxiC+srfN33f0M2GeaZWSn6qD+8X/MO1PaXur+xp+cQrvj3NrjWErFqG0sWTHl/G
Fy7dtYU3b5clI8aV9RLJEYJg84yAoH9604MLCGwqlXtdWgd2aepOnwriaFsv9My/DJn02zdxbCHT
vTFMcMDUAL5PqLMVm32OleDzNmVck0vFjTnqoOjxbhXN6cTpw6XO5EDrPU/DcZ7tyn7l6LAuLE52
n6CJUqV8KmUBayHCLnX3VfZRY8DQdXaVRI7N+OVskAnS66uTA8VUOxbkUADuvEwYHDn5co2IFNRR
UIx4GdPPgSBi5UFJKV8voNxlY3eSXdUq98hh2lbKG3C84rrAjHVGFPv43DAwdeoM1m3fq6+4OMXl
+iedKScVIEGtsh46lgQjcO0j/yniK6N96JSvn1CObIeFsWUwS4c9+3YbmmD8ATM6/OSVUmaseKHt
jnrn9CbqoH6zXQnjGizfhrSSiuHl41Y80BR2gX9qTmiOpLgsk0JSsyrjvqHI9RdNqXf39zAg/TcO
isMiG+FEq0dGzC++loBGOaTziHDorOa/Om5RkY+qjL/z25NjPctsNaoDhLhbnZOewqOPclU8XDCc
6Gq9nH2Z18L9rSYOFa7v50FlWfl8bi+09JZbb0APcMKjs9tEJZsBBhKq0vS1R2QS82GyhztXLQXU
WCriComoCe+MFbDsn3WL/tiagP6hVC9JSloAn+NimneXVo2RX3k1lQRmwKQ/+INO7ODRjINfWfcI
kqSAuJSFcXf2AjSPia4VhXU1EMFbBduoC/7pkFLoT/derlNrmoRLX0iy4ZABcsKSF1MxC4SXaZ0i
jfxk/avwSvGDlbqVySVHUuJcU/0CYPMD79m2PNwkiCtYOBiQ1Lu9Zin9mqF/BfikQTgFhDYY7PgW
EYvHicEScaJZjxAmrwJqrRRDI91athon6HVYQvKfkwNTSmSfUNdOAu8qI266sm7Tmn9QcZrWecrt
ZuvKi9HFbs5jid3tDYftswV9ABrFufFlVMYSt3dHqUYV6Y+RF8vZYq8mXQ9t42/MfKHnsXGW0QiA
T6e+/1qHhpWcvSNnKGeQuk0pjy6JsHi4aUaM44ttvwR406OrEtIsjJuLY//i9kJBVoJP2ctCp9yM
VkAMwnBaFsjdrBeK0XtcLgXcz/WilRGGAZZyfBYw50gSS4OVcH6tZc0BxhHhKp/puc+CXBJMlwFW
4sKFSP7wQXUPhi8EQW15PuluiOlblHxCcqOGMUDv8BWJvEwremYM8SyuLqPrvr6UPVes7LDaCKmc
QLOdycvRK/wMpwfkX5b9yJ/gRgrI2mXW0cT9Rox87ClrQL6qa4JIhUbtX1Zc0nXDDBunSWl36bGV
ljTSySpWRBs3hbzJuqb9kUMoJ/jaDic403cMQzbfV1v7N4OJl+QAxai16VZDR6pK2v2tnV+XrLfC
b/GZkYzS9cYj69dz/Orc574flEcu8YWhSz3tZSfKnj7bLk314RQLWwHVIitl8GORDf+v7r5UcIXt
XCtKG6E+yiU0cRtADPg3sMA3MAT9hxHfLI4BmIWH+avKaThwPfv/WXiNe6bNMJjkwxFoHAPa+AU8
GqP4axqRUUdrHYv+guysInM9ZvC/sHKDVZac0EmS8lqiwF3+AnkHqgHeqoBAA4vPzivAxRnUGmqi
RSnDp26NgUiyR0lBQ1Xp2qg7dqo1jNamMqd7MVwc5pQEvipGE8AkprnuBdytEmXuoXSVGPtevgw9
SrkBhK7p9xRkmzhtxefxOXRnANJ1cxxb7naeZAyQzJf7J3aYFwod8FXtgXqkHosroDzKVnyYhRii
RX8weFDqhGbwAidJTxTnlNI3MBxQHCg5VwwrDuzy2n/o0UMW0zpURdBtlpOk6aVFkKfIA0yW9SUS
pki5bj8EbE2PvX+GW0JfkgO4+2wUWMo/QzOt8rLVSQD8aD3fGs7HJQYq+eI7j3zhRScp5gUtA/+A
F9tyzduEe/SM+tD17CY41V4HquV4NAmGzRhxHvfkwSGhXo0ZWq0gh76jtUShFY4HipWBAQbmXiGc
S8eyaaSHH2k8i86R8GToicM6FSYUTpK9LS7nzUNoKZQrjzbgxBjwY4JD6CYWybmUId8h/+/PRlNr
pwwAMijQjbk6jAqywKWY9R0Wun6WXli9989I+xmXf9EqQLwCccv2NYCA/vHWuf7XUYrpwnZP2VEn
Q67q2fyJk3gKJCPbYQuquZOY3yWwFejyA14gMMyIgA264w2C3Z9amPvqxPQUUwPKWzOQL1/Kfp6U
PDaAZSN9dIbBf0MXhHX80P83Oxsn016qD1c7m7WZvx4Vp9x6yqiaFitJ1wJPvak8+mbL/idiqSPb
gLmhEbcZOMgFTKw9W/SSbCOqwcXZ0gpE0v1yJFqMs/QeHowtAo3x0mNTcRTKxOn+zmpQO0IT647Z
zuESWf4uKF8/a5wRL3UEj2QUBvVUIvVO8cSbcMQjWvpXXMti6QjqrVi992bL5JcmkOfiwmskCWJq
IyEzJ60lSe0+7HFMERqjYKHloYz+fZSzJ7imLDdKOLvIo4Y2sdGXYsVNnvfBG5FwBYrwD2ysVv9M
kQtcI4Ar3jQ2CeK1gSPBp/2symnGZdPQhsG32eHmspoenWhhOr6DMZpykyphtkfeE6DxtUZpWhRc
5SRETHoNeimstXOFPK421EFwSeI43vuq8j+X/OC7WIpwbQ2khzbSQiTfCd0GoBue3JLFRLj+HZij
nF+eCCMEMAgnXI/xDdOt4xykkE6pmEeg7HFRScXfS802x9rP3bJ8xfthclUb394BnlyttguWAeaK
nCfIiTWBX5JlGWvzz4mQ+TyTBTlg128DJryUxn07ibHvoojiQdXyvAtp1WQKdYB5W/KRh8nPh103
Ws+Ns5+s/8PxeTyzg6XPqtHky1mH5P51CfWH2t+xIp4rTRmT/wIM0y3hDv5OS4WcQX3n/iZ5ogPi
EWBm0bVlGzaggeVh2b6IDU7nqtPds1e7gEWAIUnT0z55T4Jc6/YYupZ6swW0SF51B/x2bYFbuWMi
17JBRy3JJpPjNTIi2Xf2v32dsVU4av3nMnylx1JVUDW3UURYjmkCSu6fhpdWzqnNfBpROJKCHNLy
hE5ZIiYosXNx4AXiR35sDTfJei5cxtYA1S808EEOcHK9/jupTsGa8gRiJoA/zPdUyGuZ4eHlNIqT
Z3eI11LKkebc7IOMgdsejj6AxMdBZllHCGoddas8JrT4AdOx39QXyvt3/vEJGFeUmAEcZJm11fpw
jqYT0XnBri4bqrqMtntWEQ2qAlXppjn7ByBB46djczuLMuKJ99zZ126PxpTREbbcLfXLCN62uDMs
FQfE1RaDo5tDJFinr+64ixoqn84DZcw3dan/YWWxrKX7eDa3M1LEXdfe1QaqMGFBc9fCRuC5x6h5
VK4vlVUOug/zXVCPxJXVAK1uFp0yAW5/jgFA2Lsa6UnflDMIIq1QnD7JRZrHvl6+aANOUL22AF3u
mSPx//RzFJcfbt9UmMZfFkL58VgjVshcjRCL+IEPiL5yABYjlbD7EARXES2fPOyegZCJ278j5zmI
5srVFEmVodhqXJE9KbJNDCyW2sdE5xY8N/sVbkCt0xwy1frLau+7HfcLXrsy1LnO60fntIDMklJB
Ne7MPUoyJ2EuX0nSfF8HFdlp9IxH3ALwmtrAZLHB/ejhw5gJZHoTvwJhsIT/kM7NudndXnxv0u8m
ldhDJcNsygrkazti3cC8kDVN/13MXSoYVODQXCI6q7q96owRFoy2HoCrfHVPsvaqymBsFekmy8YQ
G87VM52zPqUUtiC+Rc5gm/xYfryNBrX4/PlIE4ZruycxD61wO3iW2Rcr7UwX1cj1PDjvnoXmBUP/
Bys9skdiBLozNOrs4fmrVaPHvhYyykJ9fLOE4mX+0nJ47gr8Go2+QC6m2Pb1CUWKVObrKPD1SROw
wIDvMvVSdr+kZ2KlRwCPPy7bQol8cfUSSgr7ODMt6d0RLU1XETms3oCOiAY9JTj2MinShwbREBQx
y6hC1IrEKK0vbVeV93z95KIeRx99gKOEPIGhoMebIV5lPrDqO8YDRIflx1qKIIptgWCvqxY6cvjI
IdMXWtsgnVacqX2OsZlmt1dPDIBlMHqq7pCSVMF7yRZqZQDJiVf+sBsDy/gQOoXBTf+1Ik8+sViX
CzVFKopK1LgcgOGc6hihCweZFRhwBrRipkSRTn/mCKfGYYF462mQxKHijLRHF5e9WnMOlPI6EeMz
oNU1KLHBK/Rpc+3AVsex333lVuIK0qmc2lPKRaNlEbRyjqWKHve15fNT2WZmI27UOdVYJyr/xebo
MhGwvn7RN4uk9YV0lDtzcud3itWke3M9GIOn9T1qs2YogOxkGIG9WAAPXjTkhwn+HJhn6ZTyyAYz
HI2WMs+cWxsd3qVBIq0u9kfWEQ1jN68WkPCq3XLXmV9mi0yQOHj402IWnHKy7vQrweqKog9FwXNI
Q3aVdccEeiGhqwNJWw7OAhY8VO4MGioRNah+5dQ1s3t+Pp15ksJKm5rU9cx04U/KpedFFP1UFqW1
O/Hi7N3eU1BQ8LHaAvTIY+eQKZ4iG0Sl1iac9hXHxsxiQKiBUDo+tTCIHScj1jYhvTWjqjtIXVk2
/2K/sFkFj2TtS6xvR48YCZS9oSYMkXVG3Nb0FU0Xre1AEchHelJN+Mo1dkRYU5xdv9Ot6lCsdKB+
iVyUp2rbwg2VfaSNlJpDQ1Myn86wOr9/CIXFhb/cn9VKEdRDot4lNAC8f7rAI653V8eegwBMKFDZ
iaArAfpj8hCL46xHpj3gEYLPHMzIuN5O9ulRECEsAyD1ktFGQtHMSm/YWaX0AQL9nnrkQEdZSm9e
xC+4iMgj9G7ROCGeyjvYR8XfNfnR88lh2jjWs11XtAbkcmkBqNjGC3DN4TyhMsJIZ8kqUAlq+oSn
ix6iiByZ5EHXeBrgGYmGNa0CnqbctHiuy01CnZG49y0wXiNlU30k4R0Cw8c7xDoM9J5gRVyJdmPF
1epeYvAHdflzEoquNkOrcInLcxXk54XQAvqPQckMJrc85XJafk2bT0G0zOm1AKCjoQ0pKGUhJOac
w70Ocqafxn9VRBaOcEhR8fsjvhotLWN3dzykL26h8OWVIEwVHL+UdFd1DUBlpYTCWx1hwPo6OfuB
6xeBMWy8cHy5ETGbJ/GWOZMaia5AlpJWub7J6OcJBD+XrHTOnQjhD7oTRvLU8/WCrIpJUjQYm2Zp
jJMEiQAwvWni4ivcr1xFhb47T15ZN/Gl6NKR+QuJ/986Hz6ZO1MaNqyvleqdspQfoDKs5VrVCq69
vp7KHtD+9Gw0aoSOBMyTZQppFE8R/sSbrYPgF7CkTTlZJwlRIORagC+rtXSs9EGqctPGn4Jvc71s
wZiBzh62DqJ4z3RQYRt7qd8rhgvjV91mYswjSebNQiOHKacnsotIQ3ZUvQQlOw95v+aZ8LmglZax
QXWSB8gcNkIkGS01oFgbP4l3We8EYsx/215JRuwwHGJg0LUa2SOqRGmzelXrA9a3sEVUt3TMVV91
4Eg34dXYGjlfAReoGVlioq4bInylM7DoKCfNLNH91RCq/7IZqla2qnrSCjo+VZWWOgF0NqTYJqCu
DMRBltxyyg0gqvhFgqriXkQZROrC/iY/R+MHfDchKJptCubBKdJN3YTE2pOZdK7AJUCJA8W4fOzB
cj0V8/FtD92X61cqyL21dDIEyW8GkuAGGby65U1sYQzgCP0BFzHNKH57PGP75vetGIV6EVAgN211
FieLIg7G4RVM+I3BGJFmDJmp+abe6t9TjjZQuhbmbsPfu79dbH4pBQ4iU5xn8cdDPJI4a44fG/GO
aYBYpiHRgV9ETLmGS3+Hi88/jM0bvvSjAgEVJImFWAXB07D6nggruT7b1VDbiA7wW6lfPPcb8aE2
uIbQvSX6brMPp9sYfE2yjzz8LntHFY/7t6jEd07f172grLcTwukTmFleA7tUJnqImcpoIKPIihwi
7pRWbdMNkpJYHUFU9aKmuyqSJtF6hiURTcILcQBh6ZZMMPtfTpfiBNRvNJMmTOilqvr5hmciG+Y1
n9xyD9Pugy6oPLam3ikjSbp1vOPwdhJf2DT+q3q41ee6Q+/1B0oZszs8QqNTCHG7b9MSixz9Rhy9
XYpmUnC4bNi9BCCJiWWwhaOH4gsRvahKnJuThOk6f5x4N6TvIUHPvEA2veORUD1zH//bAXGGk8mO
4SR8SvIf4XQu4d74IOlGJAUEpIYY++2arxKKIWXtiulGqLuFnIbbAH8ylRMvuhphVQMFUTgeNNmq
exSSQXeEH2XjuAWKwlvHBIuuIq3cnlbwXS2GgXkjFpu3zQzGdiigc8NmSxM9eD/TiJaBdLioZlAa
sPtWLggssY+PSCH2sL4i1nh6xI4NeXzwofK9g9oRS4+MIJOEsU6UAVhXycV5QWBWUyNZpoe58Fp1
EIAt5b0OMLCZJrfYIgdi8rLAdG3MammQDE9bgIo5tOw9vQBIAqwceedpuEUTa7bThjLsups/5Ylz
AVDKxDgrKZJWG4m2ugbbftpAyjP84lYX3s3l4i0xCVmWv9VlXpfEAep2YPUDNPjkoILv98fwV5yJ
QEPEPv7g+DjrPQfLOkKlhnbtRd/idk6V5nKlzYT5qiLUk96hAjLpm74/mbsLdAMSrfAsIx2fyrmz
Fx4yPaC0oO8CUW3r0EVetsKpRxFyM7l13q0I13IY6c6p/2KioZLuk5hzWyjg3VHzqIqUqb0TsOMF
hZ+oq+F9zj1mCxPy6ZJMK1hCpp+D7GVJO2hoIDzfTAOLIsRVYUR8Qn9NlkecP0BTe97Ahh0vF0+e
K5dZytIJOaxuWcYPyadBWoFwfM/qZtUW9errl8vPN19AEMESY2YH+GfwwVwNgKTn09cY/kaCATAc
DK1hbQ5TrfuzuBsmOqfV41tvximD1X3CNEJbCkPwplfhxycLRNMPm2w3jtfWShe0McyMVNbC9bkY
x0MNhiw/BGXBPoIhczYwAgEBvK6UEHZsiqvNOosp3EHCgKS2X2sT51RQcvIH/Uc/SpyJX57nS8Fb
c+nxPleDoLnuYaf3j9Ro1fCONT8o7XHlrcWDZMQXMNwzYlC/cIciw+B48X0gJ7XzKmuKxK1AGwya
FOl19pGtmAiHBtOj8LwDw37WdzIpLF0b1jTdvpkK4GbzgiXMt+CNNbvQsRllpRgaj8PRuPGEn+rx
2aKGrbT1gdf0/wkR2QRSjGigCU+AbO1oFf+nm/fKv8P2zYwND5Hyt+sgUpBukuVsxo4AhGKSlAAc
U5lkvu34NRr5bYfrFAJE2ib56xCM0zW7CJrMvm/yPSL/5oMExjwZKJUu0KF27qD4fHPnb8nlz48L
tpMeNf95tKKQLeeQXQYWLMd9uSnPX4y4aqhWMIOQtekuN5G1fM4cjLUhrWSyutTGPY1Y5H0XcUqw
shcX0Tjf2I7EVhTxLS7WF3xe/2TOx03SBykNyf6kpFRxr+KzorvzxVyB5FBeZBchyPnECZS1SacA
yCDn/TYvlnJT/2gBDfkLKRdmIIE4DttG8KUB3aeJzqEXCBUpN8HUnWVY2TRB/LUBzFHVzlsUE1hJ
ejUjO+40Pq9JAA9rOO8hWQPf+atORWUheXTxGzYboNfpRwp4YCCv+QrgZ62Tb+1ZimC5S05q/NfR
F2Kn24on3/4XB4GnV4ra/JB5HRsPUP6dDi4deICwAD7pkqupmH/5S7hPNOh9V2nJQ0MQDGdlrReE
/fpZ8v1yot253VB8uL95/s8u8Dy0D31l7vm78DNyRj2AEL/rThScum6wRXY73+56CCE+ZCDjLo0g
4V/JXKYc60iRdXixy4G8uez7P6Z8lE2QVqVRvs/1FE5mbyFwCElqaj+Mn12oLlTuzyc8uFm1LgxI
VtRQl9/Hoho/PGLZhLnTnCmv2YtEGhQsSvmgZeClFRqMCObOeUPQ/+JSniaeD/ylfeGfFHn6OIPy
A5wTUGnoHIiZq2c+/hugjk3HAkOTzRraINYHO82npVyp1BIJRGT92Us6/oPay5WkaRYOh2JVBA1n
akI1MsoWq4Ci8T3nJNnqbpqZlTqfiU4yBVrC7lm17wGDQeYaAMgpRcUJnTBlGjFVjzue0pO2/SdZ
Lb5S3uhcaEMz1QCQ1k44aVVhjvTubqVTd+scwXXcqLo3siTsQlAk4GmgbHIeoeLRDDVTxvvdoTxW
g7sCFNOOjR0EI0OWDQjSJZklaoJDbjOIT83CB28UI0+iLBtZK4o+qThcN0ocf+6/wPAY7x3l5tGX
rVTfXlduHUCRrMPCc+bPYR3mQqjkPr4XGkzjut+CQmjtYc1taff1onkoUhvFPX6x3BNzHuVsRaUR
lqX0BrkQtqZKI1gabkTOeSvERwYBzlDQKKVB2x16wTJeqmUOviHXsqJss/OW49z2EL8WS9LYryOZ
54ygjySJE1qFwdbtGfp0pQRUAWzQ64FbYTfVu4KeMaVg9z/SHLeJV2l329m8SOZE3NBVmy0m4xAS
UTFRhP2wQ9YA7GmqisUv7TaDq4WXSdk6yk1whcCcUH29ar8HFMWnTfphw9nFDCnU3TB7JZPZ51T4
pVJoKEKPLtZmlaLJHpqvRL1zHvDnO9CdC2rz30o52u5YDcSxuNmW2Gw9ThA2pR1tFM/yeI28ftvv
NRGns/NBaFhC+Qx4C800Fy3HOeG6o0uu6UD31+ji4ZCH95FxYBv4/0WYGMoJMtyNud+j/0w9qJAi
z/okzB1YCivUrC3hiSNiQ0p0GxASx0SGlHuRCD27g7Mb+EklVHv8tclj0c/ORvtKN8ZFC9vqhC6p
YLZ18EnH+CNy89U3FTvtJ18YJBKdjSCd7Pf0iRets+y56mzozpX9GM+aRdZUQplU9GOjySb72ojc
ko7IbEB1cyAfm1iJv4HQOYlzNZYLbDgiX8LrIwSZHUeoWXDnnnL3zN5vnQpEcXafv4r6cZzDfmGI
/IWnn5MqeBmJF2AybvwQ8XauDW0Q+2uI/lSLg/UwbWvf/kLFA2/HlwXNFXCshkUMfN58SE3CF9X6
Eh3bnBTDsGw0PT+h1+yWsInogNxzVRD5X+GlaenPbSzZF0nfxl7ikDN+/vJEeAQD4ISAMNZmcBe3
r/Po3bncBGSzylmYkZZzd4Yjq0VBz4yXLOepsxbhpkElUyuhh1Y09arsV8KHbCeeuH6QYXnngG3v
LGZuW+Fnvnswbuu90XUjZGre/3g9oqwRhg6mhGyCAY+ON5zVpnYesHyAwwMqA+YJjDKTrFOBob1I
wDpit6OhgC+sCK1wM790VAXGHnBovf6VtA+qlM89qYDXD7uM4qrNsMvZRjJVV4lM/VZHfqkmnRdo
8FUtbV1qGkkbPbH6CaspcndZX7cRAa3nE9OHm7dXyYl8kTC0yfh0et3QHxRNDT2e5scPepHB6LFg
hz2Vzpt3TerNc+HJGUlA8OBaly0n689ZoOd7ReklpkL+T00fPIj+p6MT5i6ZaZC7HEU36LxBgTao
dO39ts+ubQOP83MKv8baJ1UudYN4iu5C5jCNjsdH1auSYHWoW1f1NYn2OLO7A5GvY8HpuTRSqAYV
ZW0Lb9jKvWrs/+mIOZQR7K0ESldmjyNcvVRTeQxpmXHMBNWMJb+KSqkdwK/490D60CehjXSesjpF
eavVQD2WpY6ZmcyDD0WbqTrtT21SaIJC2Tk3DfhYN9c86udXf4qyiZcdcLBBRb+fpPzjkejeU7s0
SVS+pJ0EXHkOgrfX0z9gQftGQZz604643YSwvI3h3hAYZuFpB1nJqUebzwUfe7wYuEUBCRBepvvN
mzVCclRSt9QZ/9SgN7ED+HXGAqIVm7cOppBTn4bXtqTTizwbOfRfh3ST5YzakZAomlUnNsjQQ3TB
c0erMToIb6xaeBs/X39rQF1s618L8KXTQ7T+N7NiCbArmuPIn5GPYXOhEnCQ5HeZdd17stxe+w0U
D6wHb/ajwqnns5C/3uWyIxp3YkQWrSy4CK1qZyX0NUHmVc/sX+L1yvtZBDMECDgGYOYIGBsZsp0F
q3QiBnABluCA/5aCb9Xdu5Gq9zfbI0gdZyMODfDDwtSYUWVwef+Plwbez232zXswXz2FTyFzQ6GH
rwjEa4rBtdOlAzeL4ofvUrjWiJo4wLQUr2feJP6hMCAoZvWKgc+Z0vHEB849FqHDGjaMUKXgeR8B
mVT5u8E1ZLRCr+24/obrJ0gveJWduy/sc1WYRTuFTERjmcVrSe/AQrMx/a1bEX3XXvjdI5BswIAT
UTmKCq3uqso/rf+c01B9GtdZgiSZR/d4rkgqCLF+c1ncmf6+RhYAqdbUgU9Yb3g1I6J2oMyodQfA
VT8ZvHIRbDat0yBJF72Ud3hY+FxlzdDeHC+uuHpQWYVdd3piyBcQ9W0Q5r1ozxnF2YLYTnnIPTzT
iQtMjdmW4gcGAvPshcHVqdlWKRbbvDFk9To4Fipu+YGpyXnj5pQ/wV4wXOLuQnpNdH/ifwmFM5hE
Zy/qbR/Ae3jgMYSk81U2oUvv0Lgds7AltTvpH9tAMQwl28KvdIsWkcPOka/9IacNHQTLGYtNs87I
+gJv2K2pQ+XZf8RGKp3O7gjo7TUIdol5TbJObUtWpIvKDrDyQvzTc1goT+YQ6btgV6MGfEkajJvT
sACt++1RFX1WCOMAHXMV11wFCmEw0Zq8A2rYARCMW1cwHQGhxAN+QqXp960+COsw9qPCddZdwgoE
qq3HYVs/d7ci1hESJccHXV3lHqvCy6SdGxs/vgJfpwS5i7Z78Ehlppuz3H4LXLUfTf2YIG5mS6r9
+eLgiKrJoXYAnz1hRUD2uAMJYhumk2iB/6dZ3J8AADt/Y4gk0Yfb25iZ5Gj8jyN1zCd2XbcGE/ZA
8+wucHG9StBQ6ThMbVoR1wt+bhGW0mS9eV81cBvaygt8plJVJVFlLEdDm1MEOF7x4qtVwT8C+tCc
9Ur3g/80CYlU/3mOmft65/89MG3ZH5Cb0zC5+br13mhDMHcV6bgf2BI8Ck6RLBoopyR9vjPl4l8B
lW2i/odeXwsPBQc0MEtUZfeMmPq0NQUYXBuUDgUaOIPEo2bjgUk9OvGGaLgBX3W5LvlvhFwMqxvx
wzfFDAPwIf2DTssxrY3nBtLTSY40abLKUlJ30kVqtbo16voqSw/00pd7O7CSH6StRUIel9MJjmPY
bi6D4Hl5UD0Wth0tVIqXp2q5qHUgev+5dKxrW8N9bme3se4GRk2C0XIOIh8Wm9XAuF3OHCNmEC3F
YsId6xH6ysKzuKPqmKi0n9OTIqstr0hDYWYw03ec6hxqLe3dCyDsdj/2oPZOOH6+OKtSr6G9eAZh
Au+1K316O/vIBVfUqEBIO4BuEI8iFst4U59xzniv7N8z7+KHBO1A/mp6jhoOcvsYH1zhM1vnHbBU
pg5gGGYt6AWqZm3x+Q/nezK778GxTtwSxuFG31R5MP/7G1W7hgh7cx1XGqvOI06bzWmoE3UB3+e6
4SD6obAvOOPw5IYAQf4Az2uIGSIkZkfBzXzCGysk2airM0pvkhBRRpmwWsZowv2Sh1ncY6ZlKRNE
7mTYqmF1Fbd/L41bwXN40/cGA+BqXzVGDKk3sROTdr5IFEsvXPRq1/zOk0cP+dHsDqtf3usHwSpn
6WmpGI657gT7N7tGUlKiLuwwacWlELjrght0ziUcX7r/l4SUOKuz+bjWiHIraXk2l3j56ZAbmZf+
lEBR41HG4jgCIW0Pq7NzU9gocBNMbcRYDwhSRo+Iihg5e2M588Yl+blbRWiZH3oR25oqFgYknpFj
NrCAj7zvgYnodKj6oQSZj1mUPAf8Y0k32buGW36XWdHA3BGAiqFm0oFy/DR+2BTYheRnpWJd5Lob
EalFtrzj5qkhhAVS+aN6QegV7XUutOCRz1eAObQGyDaa6OSkgdwROd/vMuOVh+Ee7NJ4gcZiVfWR
J8gDoEa2UakIUlyTy9T4i3Th+S2s2JLi6KoMN5GBLCMd8+BfgyiskXKDJ6E9nzIeY8QjTfDPiXBq
1dxJmRPiOa+ciNviDDRTptlzTeiyQReTkHfKMihL/25P5FTEMTGGG0d0uhwLPhMZpMGgJL5aE2hf
25XXYpyaIxyWVijb50sr4m/ddnJn09ckB126vtMzz7pPMNhiZAV1YxR9NBcY2Qw/nL12m4t49niw
2trXrTOe2cuvkXKzNTS6Qbg5r7ddzzpPx7e9nNASzCD5NQ2HNUId+Fayt3bvJ74XBFk4uso8DkeB
VqvtJ3GVSaT/AJn9RPREif2LcCUMWd2uL02CNhR0bLKQ3bWMqcZYm3O95hwjvy2zAAMqSfftxnwE
R/3KCjXWZzeLYZ6G1gQRfXZUc9eSN5oxa6McW3C3NHrJDNxxb2+db0j95Ra5f7DuyWEG90YxXdVV
u5bVe2OlEVpgAIfu8FnZfA4BcogP6Iq3itUl9FrDi5KKNZKobmolJVoxPlXalyQxv6ZovnZQu0gF
GEoUazCbkSs/We5nN3dGJL72b/7pmA/xnu5zQSkiwDc9reM1iej3bsyAqoSjsdhJldUvAn/Hb6HK
p/rToPm18tgqc89zhNszs1WNJF18RLOpMB3kaaytx8gBjeivVRqM9xLivn9YJWPnp1/Jg+1tF3hc
gTIvUoprEZP6vO5JqMciNNhMI/9ppSjcZ8m6bKVA4nxiH5WtE9aBsLpGYR5iFiltwtItGmo557bT
VeI5uJKVs6wLDEAUlAAgjqtU8JMdsiz0XJW8DdZJRd0F5FXLfR87a6xustuS8f7TYXAjgdtCPXiT
guO7HoVq98iXTzWP5sXjy6BKXyY/6SmtOvk5FwumvRfbo6s0F4urf20+ODGlVIqeLGvxzxQpCNsz
adLt198YRvkHE5ZdIqEYZiAyNBqVKE4gQfuJBS8h0EjDHWakj2w3broJtMeJ6uQuMmn4kEdsZaoo
/UOkKewBQ3yP9njSYsdjul6d06PF6vGtkcXLh87ebkoSO8RbDt9VSr4j+pfwnFIxWB5kzqWTJ66Q
Gy6iUar0zqNaQ3vHD4LxU5Hkn4AALAeNc2vxjNxpogMr4nbV3+q+77BTP3p5KRamVPykHNJSUM/Q
fpGx2XKzDsdoJngXh9Ymb9eKf5bX441vsi4zScBhk60bFJyV3G8pCGKSYaCftO1T3LPSji9Yyho+
0ZqSQXmKSM6ST0+HOdp00+e28df8xlp80bSCUQ8uqOQt31ln/NPXaYI0/h6rBLwP+MJ2p1tSLclT
XSqapqeGrLYVPC2tmGJ4DkP+3qWKejiI30N6Draw82czxqt+IFQtD0XuwVlZIlDY1lg6fqFVBxo6
xkFiWe3qcmVAedgXjvWeyqauc3krd1yGD9gtJJQoUJ1U7VlfCnt4SE5C34JtlVSnKJRBObPXcKek
EKlaXi5r9/JA90I25XkUJqPJcXil38pN2GDTyqtTvDTW83vUloWck6Yl5b2ZEvvjAMr8/YhgJoM1
UqQr4/SKkqNYZ2kQS1StyJNJ5+kHsGz9/xiwN2sor54VFqNO5eKw7NTAmqIPhLMU2trnGWOqV86G
BL5uX3EVgrwJkjDiLpBIiQDXC23K+LMYrOpg0fm0XIbkekt/4EgvWk/CEneQdUxFvsvVrhsQXIEW
WP9GKc4Ij/s0WvyOqN3Fsa3JIRTWmVi8+r/sATM/dZ5HZRH5LoiHfqrdsT4YvGibNRxqaTBZ6dC9
Og8kogfSSzUcwKo+JZDS+wQOrzumhtCQg2pJwUOHp+G6CGJ4ysjLTjl3RYRbH2kQZmA1p260nNCL
ZxzBUGDpTHWTyV17MV06/4BJj/C/RlXM2T8nQAFXeCCFweWx2GA6ndwqvzVtewjDbyEgZqg5/sce
scMFp5RftlnpBEba+FAwZYTIa0oCZHy2WBrASwZef8/+KFqp1x8MaPuAMiXBc91xuXSKWVkgMO0Z
HdoFdW1UfA3EouF8tqEdnvYaNHKiku6iVu0HSmCeTjMStQaqcEs/t6lhI4q7z3FuzwS41WAfjMKw
VTO3ft4AELvyzdalsUW07XlQjJfN7KcjSD0Pmf6WqW1v+9y9WhCRcTXxTzzDSe+gnzuQO/Q6pRXB
jVwd7WTX+ecxz7HIwGj3VKedbWqHgxgA9Hca30zyWIzlIWMNpOPH0QKHpxa/eKhhRwocNZoICI3q
dtz/XcHWxjWRS+Vxp3FIDNd9aLYzs3cnybMYe8BRpOZ3aX/HrGQ5Kcd1x9iGXRNJzGeL2n+D104P
OqzhNyLyb3jUZjl+Bs+MmJBmVbES9qzx2wjCuWE1j20bOT4DQZKYG6pBzpANVEBVgZQZbGV3Mlhh
xh2RQZVGbsCbmVHenyOIqbuxIp82rXdSh6OcUZO5m47Ee+U0wOvRy2SdvBa1jf80TxPXTOT6EABz
dN1kJY5v6CTIR/w8Y4kWiU+b8aAmKmpTNzLQ2ICvRnRHKCYTe4k+OTLVZl2ZnLOMATIKifWou68B
gOsszzk/YB/WrAbPCzcfPkG51F1obigeqPYn9RpTzUJdGsbcVFwpk2PfjAgTwnGVbMiqNqYKj5nV
wbTgypPvXgwJ9M3YvFJIzKAaj+uMNb3EqBh0pbfV4Mqf2SdzJpl1SXXzZ5r9BJy0+HkGeTDsKjYP
Ff+uQBH81JAEHzE7aaQXnJMUMycTxMAQTzi1L+UcyGWBB6oVeLRM4w2Fn/jag94sDJi0u+3ECGAy
8FKZ99pfFJFXs70Qby4bahIrDomKOgICXHWF1VbVs313Eqi9CehpBzw0pM7ZHsnI+pZWfzdUjtQA
RJJbb5QPvAhwwK1EymQEFZjp0YqlPg/ONNysWSL42Zmm1DakozJ13khR8kRqJRHWvvUdhpsS3r+X
sfgbBTSGy/G44Ssi/PgcSqg6lYKW3XEZPoJze0RnGTmgX2O1vkLyQ4T8tAzMbh8wBO9GjsOBiSF9
5aq7P0qbkGuwQdjSoMVp9FLVuAvzjFuwgQqpdor5QNOkEonJCTPQw41PONLxnh3DbKpuSLyBw3tx
HsEcF23PP4cpWQqSWqcZzBN6/TclLoG5h/t/JB6z+KOtbXdX/tbLyTOxORVWf25NgoJTfGathCMm
Ft0knm9U0j8VVS1XmzDzty/jfgjwhKPMPBPxnFUs0VYVnzo1CxCDeXJSxrT3Mv8dkWO94oj+ocML
B2uQtZnK+VaX76oCQ5aAOki9lT3f6A5eowWSfxwwY6Ep+CLHF4CchI+IjavVBVGlMFsTZtGFWz/3
2jn5GSxelFWRJtalwQDrHBrSKFmDbXzns66w497jBqw4n1IpXSLGJIoeAwWD3vQWSAafKmPhyhgT
qTh6ZNG7xZHHLp1rK2iQreszr38b4DWz3+kM+2gGg7D1X4t7GZCq7516ti9dUSuOPJj2eQ3S85Rx
GU7ijMG7IUDwrOFYq8xSlXV+sYfSVgo8Jgzq5LB/cXhrxiAM6+s14HTKAKziUqXf66EtMB5fSeU8
PgDw27P+kEpDSRFdqLr5KlqjnUIm8JMoBl2ecvr7dk6mCaDKHDSh7g2uz66xmjBTSIFaefENoZ1/
uUse2INTWmRX6jmaT44LtIoenF1s8o0LqU0icDUknAqs9hrFJ52VsMKZQ8sPSzJEg4iGwMh6Lfdb
KFyC80xL070zKkNROISU6H9XlfCTb4XRGD2L7Rb2gL2ZkwkY57+oC0PyyfVSqVbupQkXKDZJA6gT
btPJnjRnk3vydtwbkex8IPz2BrGqN3jRjC8qScrvOCHcote7SZTxkucT1vdcCOJbc41zcwa/bUI8
Am7ufMmLyNTsQ9IqiV7h61OBXHnv7+R0esoQumUf6PRKvd4RzCnnOwx7WsPZSnU7LcG3JDvesxXn
HMTAIS44pTfz+gJ5m677iFH8OjU3eJGhSyKHj5MGeBJ5dx/jvKbXmjypIY/l9bDlRwxnqIP4N6E2
NRYekIxtoPl3CJHAX691CARJPUuXvGu5111P7+qmsmZzZ5fBhi+z0PVWuONyXbuPV7oQ5eYMkDpQ
wpyC7E+HelINiHrnWU8FY3vhmmOWJoguDJ+cDPSD21vVg/jPQpVmkIb43/MsilM4Q2MtY7hjOk0B
0ziwolnuJGr87mrjGavMIw2vzwKfbW5NMGxMcnCQKOC88jkLORzYb44rANDb99D1uwQPbufEWrkN
e7UW5elUIzLpnerdIS2cS26Pu/XEfTYJHL3KSdf1O2tCqcOuVZSQtsH3TGp1Rety7VzQogmBaotl
awamikAkiFuw7tw/8wOR7uIHft30zL2uqqI63IIgCblT/v+Rwz4RoS8QF6Ip72ACRbepd1zG3j+d
7KofU0HoJ+0pyLb1WuevcE1bfH3YSGUjGt5UoraU4KziWcS8XhC4RhAgfhnJh+81GqHDiA4FHWyi
itkREch330Ql78290FlSLWiVNTLhWPZRoG5HHzq6me4/+WvsU20P+E93GkN8NY8lMvO5PjTlSa2V
WuheTrEL8CiuLah2k0n8QZnuOB4SOHVdLu0HTEjowi9vhsFyTx6TVCWATK5qy8O2LC6PXI3x4O4i
lVB8ocnSxh6lLo3yMAfXgM/z5mpF+hRF3OJLTWeWSdwh44OkK+iy/u3PxyM6x394/g80IYQGDYJ0
6lqaRiixxEHUIBCz48uT3xnfM4rUs0qHv82A9Gdn6UEh/krLmjYnLkIhjmnR5Ji8j3fYWDqClLY4
2JRH5odzmCxBSinlfi1zmZW251xowI7NuHEw+dBRhImiW7UqIh9o27ewAcqbYZoz6yO1t7jfcNZ9
X9WQRUay30U4ImDYnXDNrKUjcps4rXBub3kssveSQpoiWhJ2llIXGCOnhuQSIaXodUINTCqaVAZb
txW3wIMXRhBxdAUkFOFx2w49h45/RT1ztwY8n16a+jw5D9h9QjyHLsTR7hvDz0Ae7ufxUnBIvJ2O
LnwxWVXrGBMqv2KS4PYje2uTWnWWubRK63ZxbJxN/POTV6UfKBPYdTRqID/T78pPydN59OCm8yEY
43sirzwn0CuqkvHtPlJcN6jqcghI5obR1aZA6KUOc8z99kPqDqUJWlpToe7zJizQWh2vdI3ocGR/
H1rF0lp/wtjZQhPeZD5lgzz13H/eQ/cq4BVettoPqURFXoLwxg+hTWeMANsO1noJrBgWBFsEWPOh
ehU/8Hz1dIJQGUwTvj2gPq5roXEG+UMJd8wOR8Lm4D2NTDMJtIWiiaWGlS2ZsagzBis5t20BK9Q8
TGz/O9G79EiHuLYe4FikPUSija0geqMFsMz4AXwiU+enn1R+/XkVmT9Yduc6gpN9eZE3lbDoVwVs
mqoq8BdJVFBHpV4hWu1wgzReNVekSLVrTAyl08KMCdwMf3Z4FCiBb7mB+6iiSsr/xxOV82i/6VxA
USS+PGzcXto+Eq7kxdzTbDNDXLb0y8kP5/ZMtTwi5hnHhFDGdOu71m7hj0Ig3RqKPZiCjBqL0a8Q
fUSHAeJramal0gZ1CviJ8+lXWJycu9mISQGgT7LeozM3w6vgChnElsnb8iRJGC+OHpAq346hG6Vy
e4hoiELVKXKz30EePSraT8Kf0tnKZpaXdFZ1ex2g3hxcoxkx0NiBpApi8rpPFljFU9hixDZ+72Xj
/PdzGWfiXfcRoFmUvwaeyGM6AMb+QmJDzEccg9M6G8Ggx3hK/9X382VFXQkgKju6J51ZOJBuSMt8
bH967JywuI2vJmeKMkwCgGTGTiU8uzUs78gmmyuyBTiNnwK3T6kJTYl8wyPdPEA6wLF0/uNYHvF2
UAS9vHaSsdJq0iyzs0T2oiHGP8XFrcK3mkC2GXJ4mbaEtPDa0/WHDTed30vlWQFpAFK6toGaKy9w
4lag5u5PN0ct9mqXKFDbtkzSJKM9cOeieJwTVZDP6IdeJwQXTPLwQg4OL9tJhOER6y7/Jlx/VW5/
097AAHuuG4k6VLvgXhFWkrE9lc2hm/KsJifjWnyWJgDsnA51JlUJGQOZtK+27v95RA+Bvi5JaALc
W0+RjTyDCiV1wsZKOnMaQJbJUPVcwfVCvRb8FfaDSxaBrsFGO5nuiKyACp2f0pHqNP/gmEAdIneO
n3A72HhB7EKY+4rvpxFi3Q71m3yiyDK2wSUcc0wKMfrnuNIoaCtWoML0RfXz6xXfnRO9a0V4KYoJ
eiVntyLVACHbTDsuvpy0/lDgwWel2Y8EEXH8bxyE/ADf5Rk4f1jtlnNJ8RINQqihfO5H8Ul2Mfuj
0Hj/6DZdvAbiFeFfWyRtjP/GvzU47FoJD6Uxn9zkNdAjFgtASey04MKUDyFY9LB7aGZode/v5S1I
GjTUVnrKYqsdEBLpVT6DLrIz548txFfv4/1bZJ+/6d8omJ5/3TyVkbtPNDYB524GhkAsGO7Uy1Ci
vPbg+oO/aFvDwsYZmuEqAFfD3tmXq7QhNo7m5EeLa8DUs9zVy+JH+RI9qCziAtRUcJhtw/kGM8DL
xoX6mzCHd49vo23ev2yESaJTqM5CtuLmDilhYYCXvtByko8kBNYYy9GSbZDCREDe2H08xZgSqrRL
rO5pBxsFoYELLb/bmEp4vzatY2FmZWX1W2SfrFsMcRcsbXHMjZqI96PUch87H+VvM9Ve172XsDuE
Qah8D31d7i/Km5+6F53W9Yk1pEek9YBaeFOUQUQgtHyt7LIKlxoTeFunaeqJMrsQLe2HDmERyrwJ
RtNILd32xjKZVpUfITeGm7QpdJkYsym0AA7XeCZ4tdTfxZCetqJukPV2lr/m+cqI3JcmExyEAsi9
WJjt6tikYuHDcd7POwCEzCxqy9cNGe4A2hzAU+Atiu5hjTRZs4wBzKQZfF51qaaCtlsYubM4rVG2
NX5BIVOXTxYwCHVXu0QPSLvvyKvvDL4pyplZ2TqEkQ88bbweRgh/5LErrCO5u1IHhqgXuyqFwOvQ
krZ+lS7LNcsa5RVsiiQ5dC8askV2DzwWM0szNjyi9Du6W2P7CWeSLMlM2zCHqtmiPqOhN/VjcU5M
ObG6Ljho0oMDZNi2P3RfO3hxa3JkmLvrZsrPuNwKtrd0FaLFDyhoF75DY+oQDUATSC5Q+cznSpTL
x4eS5puLHDHaQIFpbAu/gEzhe5IqPk3AZDbTC46pE5wTKgb32rFb8SJQFrCvErMt10cWI7YAwajg
/V8bxzmH7ZJOfiqdcORq3YF11K0si5rIdYjc5u8WyotNUCqTCHGxF7Wk+xrynCWrAlEW32IPJVw9
16VNyNNlmvFnbLqJ7Wl/CGNJEYk2VGfT37fTsm0dHvjx9fCtN5kfGse7/fSnVtMKNkGsV6lbuYBg
DMopxwgR2TSCDE9k3SPOWX6wAq8J+jTiv6XoRP2icnd3k9vv+Sd0zh1YIhOBJCUr8BpV9oIAfBup
auacVqyA9Aem6NnZHy7WslCuBQUdt9JOwVuEfSup29xe3yRVODQ1Uu/9HHHsQu23of6+73mgqVrU
7t6lLXQ77I516ptLmiQbq7ZWQXbdsY0yRqkmlSF8ibr5q1libqz4pz1k/KdJUK3WydUkbK9fqta6
Ci7AQXHUEAHNn88FftrJQmbxkadvuuJ30hTfVUwOGNpBUohZLF4uRJArUzWnqcOqEfzbNPT/fXsk
LgXbc+DScvyC0VSpT//jCexSwzQKS4IElBS+fYZKqvEn8qepMmDlSudWaPdDbPVXzw648Zi3IpzT
iM28qxfRizLYfZhBt+CUQkRlN5UbcqG9+h5w6AOfZoJTMn+Q3uq8PZx3x4Y4J8pDSqDF+GbAt0gK
QZ3dgrqpEErnGXFg8aso2X/r9+X/iIT5b/IXf8xslMuhHm/CaojP4ChHPz0UmqnffPna2V029oaN
ma5iYE2V+kh0mP8nj2b8U3Rcy+BTOPYr9l3sxAqXF93gyCQXzfQJGM5nuH+3z5n7sEwiU6NQFf5Q
pCLmIlBHMvoHtrROP7VWVQONmwP2L6RDfTtqJq+2+DKFv5tKXRkYeLLd6CCnBpX/FzZJ3YizGE9X
GwzuM8f1e6OzynUf89N/P/XunOhoEr92SOo95JKCd9LU15YXlGdLy5pxtHK7nKc2vDhiDpdD7YY9
RSu4x3K5kyOpAscpxCS2gdcm3d4uakJI8lhjh0bRanY1cdji9VETY4UZ8YqxQ+iBlToU41mGdIoP
EN5iipmv6olo0IObr6Riulfb4gLCU5x+R8BOgixec71MJoy6Tr2fGxZnNgcCM4WDizPjKUGqb7Am
no7/nbzZCkP4lMKxtP1kRkcUpaa+bN2q0MXPrUJszxJKXJhcZqQvG0Zt5cxQaiDaKK2n+Ke543Cn
5OAx7J3GVHcxBktF3Yb06eBDCkCJOGjkXgs4uObBSl7k/KJtev1Xq/OnTvQxjLPRuaHLhEVLADsp
cuwEr+kXl1mcoEmipk1LQPEi8d6Zuze0tLlo7h2ELTJqcxOLX6oE8xfajN7c0aXj0kmc4GF9cNjz
eFog4hRRBJsjXMuWmalgDKl/L+2MKB+XCvZUQYcP0tXjWjASzpdhDucm44mvtcrT4j15BReBsvuf
PZcR6UKJgME9e2HKMLa/cKikfeGEfcTWdmMo8osyr9TK0DJX5wJWqCEhWa7swppPZc+uOdTYrtZI
NIw8vPhKaZhtCOj+zp+akAqWZKZdVmc/CaPmzjPHDRshNQqDn/DKFgBKEGPAtz6cDMigXjfR0H/r
lwITvZcTgo2AqrfrLQ++Ql5Tx5BPqWQDu00u3ycs1i4jkYKbdhYatG5w4LJxQvv+vGlUcIvJ218B
ckC6hRJSRxgWYyk2jw0ocb4WOd/dUX2gK4qvVyNLLkgGptpeQ+f1zNa0iN8nTraXy+OvQ+oIZ1nI
dpz57rz9nZPl/KCSXFa4De0ncbdiMYzeiRNyuvGesyyGt8Rh4q6HH1xy20VSnRoJaemcnjA8pXAa
CGuCtVu6qK0+2GVRm6dEiM10WN2s3d5GwD7K/OwXsyBeD5LXz6an4PLLdDeqNlD1FqimeRZ4QpS4
YPFfbw6hkqAR3dIrcGbvC/sdvdLUVmekoBKemWKiclK7qbCqCoUPolVd9dUqXm05zZ+NK6o3BXeO
Qd0EX2V6l/QMu8OfPmaQR9DbhNpy9juB18YTGK+WtaZnY9DzmpAdoMt8iAQBRJiyg5XFjCO/AGO8
5Fh2bWJeFbWbDngGijw/pJZUwzXOmewsEX7KzWB0hrHhioN4u8QPAXIe9eHPhnJUcmlDB5WVpQiD
Gtf0ThfRUPAQWFDAgtWWgrjrWSYRIMi2TdI7Dpd1RDk4w6gzJj7kjylttBB4YtsEDhFP13Xkqsvu
bu2LUzmmDqwYcywyjzIQMkxAE4V0QruPudgPjUeDH2WDF932BYidhbHrWP43YaFju6Fdvvn21P78
7Thm2PkP2z3tcEdnZKMtwkfEMLj3VHYs0/LHhYBnFnpGPqSEkqI6R9g1MtCq/X3CIhQswK+fRvNW
FfiLJ+w+i38qBdhMa7Lcdtw6JBwfTBIHIIMmh5o7kZfRE8VzPnJj3I1nLEGZL/Fj5ZFGEmQXF+BX
ky720YG6TtnDva8AE0kf0U1Bqt/vQPr383FckSVEylGIv3m0IdKuF83qBFzWaY/beZi6PtVSrAX0
ehmBJA1X9oI97/e+Yv45+d1wQPcQTaBFIlM5dodg2u56rLoEz4z1UpCPPPivO8x5VpbsMgl9qoBQ
0ag8k515W/2ohmW6Usj88QBf1NiY9L/3G0oicrq7t7cUX43DuLfexEbsBvF6j3D1FBJ8mN1eRe0c
u4WPoS/jYE8eBeG7RWb700HmehfCD6XeGRgawb5/5kOPUky35Jh0H5661ubZBvhWLK8W0LTkLAA5
SLj/TiOjCEMvoO9aeYvGppqD3VmZserM3Mdk7kT/hpdaG2GQLg1WNgzvlvazq8N4W4qNSCXn59H8
Cr4h1cviuZ5utqd7I9tokVsxOeK4Q1X6K1XnpkI13kvxyVM+i1gCP/gmQ/9rddbW0iloO2hGCgxj
AZhovy+T8xFLDyKjRhxh9keYYcsss4HmLvjVIpjle0HJW6JMbSH7umyjV9AEmwfuhKxlC08l0EwF
Shlubo48JGZJVEFg63GikApFFIVc22120xQEF29HNbFuUYnth/b0VR9PLupLnzKy6f/kVAWomeAM
IRoc80xG36iI6VXVpbvsSNI88o0Y50fCx4wpj8wlVflU24y7igf9+X/VZiUAz1+dfZZiK68GLlXp
4SCksg8fF3qfUIveSswIUHhaAV422gZWsfvBB3K42a+X+9174sf24ZRBM+rE8huEoBUTYsSHtsdw
brbjJLM/XXB+Md+hYoruTj5JuY4NvJx4XmY8XGOzq23E5dMNiQiDyKxa2PdmuXTCxnl5gVaCNxBL
av6hc0GMUiT2XlngPLnknFE51q8cv3BZEPTnrFSjUW7qskCpflLU/Pc5j9omtZNLlObd7PT8AdiF
oxeHTH9W9Wk4S0RMcF/FKtbJ4p6zcGbiyV0gNR5MWGLYsj9ZVsaHv8GFevc85Pn11RymVM4ggzBe
skgdvz+8eogHnxOpLirUFhP/ooq3e7qcDHT9iaMSAuMQQvVbDtqHG/04x0JdxhjbcrDcsrubTGi0
hl6MMwzubQCxk5b6mrKV3rzLA8UVLcBUt+lPVhecHVP775pQPSMnjQId6x+phzNHXjkqFESUdZ8c
MPhNdzHXejF/DJM4DlNfqOcy+QM2UGRdjORrKeGBtxOixfA/OjSAlAFrIzikftQiVRmE6OOltYfS
C+5pQJu3vKaALVq86PYBxBhAjyCBahNV/grirarWPFWR7xiuzSDpcZrOlMpdgLDz5BGeGgrTrgI/
CX+PttfhtqZ+fiG8Mchs/8jVV+sGDwu7f4nmPM/lAyJmFYHXaGGmx6lrdW8/F47mjzGZNZ3svX+3
qPPzUyF9CBQCjSewf8zn4uvMxbpJLZxylvZepKk6R6OIlywNO9desMNqdwT/yVIEzSHohvU8CbQG
3JmuQDdIuCq5TJ1fFDFlh+VWi17VVMRyqtqqVXNJedcT19Y+ibVaY673WaEwXfQECIJcaWoLAY9+
nIoxohOerzQVE2NWABxjYDbJNv61hIPQLMaQBFpaXV9w3fHL7XCx7BuV2dUfWnXKX99Rq1G4bvhB
nyhXowqcLUSP3mpqAx8lbE2MwrOHd6nA0CmoLUlrMw4IWsCyLVafAg1tI/HT85L8f8rKXO0kjFfm
eiocZS9tkT0hvc+uQejc7yHF4pmtzthRN3MdguKlD7cQ6Z3f6kQUSV3kFiMmbQ06NtQ0AWPUdSUN
pQn3lvUhZwCxp0kw4kHKO1pBojiJrDSOOcEQb+iTdpnkv7jxQ795iibKmFOQEj5TyUa9nlrfsdJZ
tYEmipjDySkHsjmgH7s/Qom4nRSbsiGY4PeOWNwXTxFcUb/pB82kHUtpIdfEwxEZ2LwRruNkk3Yj
npco8VhmlaOuI1FY+YAvchKmimHjtwk4AHj+SlGaT9TSKBvHIPQP5MOS7JEuwJnYdPmeHXukDeQc
tdyYnCyi7NQ1z0PaO/PnIhe2aXsAqKFT4DMTII+Kw64wLcoposNYd3pwjC3w4Zf2CQ3dtHzJN+74
TiCLSLyh49o9dEAm1pe7+Y+n73IlzixzxbeClGrEwfc5U6mBXpnKVAQVOFPIQzT2ODkeFk48UPtg
7XLdvap9fy/1fPBYhLZSyhuAq9v18MkD1RMhopeRFk0lf8fmnCj56thwNcgvrUjJFE4d+/neF1+O
I1h0GfrLbiFbgWPLxBDLAl4Uk9Xc+YV6+LNatPUaYKvoNLhYaRwiXbhIOpna5Y1yLqfAuLADV7Pl
1UklKbXELqIjNN7zjcT5ttKR0OEvQzJJ5k5RF4zSmyaQaS+33Pg1Lfx4JMKCW57iY/xHPIuERc05
yxunPVI4AUmeMCGLkxcu0YyStY/d23awOAPF6QQHiNhXU8pfEL1c5ytXVK59B3YAlmat+ViHXBfv
h9PFGgWLGxykAcQpZ1gxFOCXX/K2pQ5epdoeqUROCbpqqeNImlvXf2Ecz1d7VuUrvxLtbY3dyvv8
1mtOJtwLFxfEnE080Jlhq0NfIwVBIcLgUfN5i4qmtQ8zoDOtGT6TJaRZ0Wkj2Hulaj6Mj+TpwFWl
AC3lrCKDZP9F28iuTzil5EjsaRUigg8UVkgNg0pDIQiIL6XpUYDAVvuq07sjYFuHO1TfFuFPpwjO
vcQ1BQvKjPxH2aCiIiJ5HjMUnkOwWuNcS2efJs5YnYoUDQQUgkHnf7PSIFjUIvVe4UUdxSpsV3X4
q1F61k2nO+ZqwabEoSzkHU7XaJEnDZQWcIhwVXaP6Sc1HKtGyq7UCbiLO1v2IgJnpvBper0nwr+1
BU4U6A5rDMlmQwnEKMIiAVFmR+CyegMmyXR3z1JrzgA14Fk/w86rAwJLj1G67+oVPcKltp8Ri01r
4gLCL+F9+kzk3VH52UUak0zV3yAMkbBlP6Q1eG6ULiREtJEj2u3vekF+9IMvAlsPLUxdk4JWxx7c
gK29izTcQbUUMUkfhz31aFLvMgIdX36EagrV6Wb5tcur/rKo+w3bqvbd9v/MZHSVb1b89EB2d3Hw
nOueiBUKOic3oO/yTEa41Dm66S3djIDamKvaoAv0Kzz2Covp7U1zJoYfUF5s2pxUOVP8LytY8M5V
gmH+JSvDtePU7APaW28lxX2suzEQVgpizCCF1nnD/pQ+r5ngMHmA1ulZErakW4cYAQNQtAC74aL1
UMf3nPHecuwi6GusDpHJQU8QOfzkMtNAhZfdD45k+uHBQIObadx4E1H94763jjx+EPkgRfdSV6M3
z/2gU5IAyBXUV8E2UuOyY6atHUJVf/X4t++wctBRFrGkzG2FFdLG+AXEKKVPyzPODkVqtnH7T94G
kjKe26g9pyOja28/HsHWLHYSzV93iGnmQ7sW00yxvQuNTczr6xNcBRhoLOBDTCriimpgTmnuwo9T
+fZXIt6V/Tgqju59EybrbIH4aFdHOHHMy4H5uwJLjggjnIhIUTmuYBtBThcxByyO66/j+nF1j6mF
cjEIJPw3XH6AIz7JrDmHVZawuXZnDpzt0jdPhkwuGKtXMISVobGSmNDqMi0NMKaF5S49aYZauS6z
/Zdikf3PiS99YDeU3ccH6CYfd3U0kO+uHWDwY6k0D+McLPE1vvh3wW1I8T/IO+HEIgb9pvDyedVA
59RbLKlb1Mpm6U0TvuR0+YwalY7KQhOTefonUBwEW2b4cjuzxgkKp25w0/eFAz5jnLwnTGSzbHtz
sFUECTK6ypW6ao1f6zlQe1jEba1+CXHJOnkWnKQml/rNVuZp2P86teyCJD0+w04aIT2GUjAu5OAt
YmKeJhulkoHTP1cJQqw7tHfVTExIvKRHQgMjAz9ozt1mUd0CkpOJPqd9fUYhYuDbrv148W18hEFb
Yn1/COZf4eEZ4btZfnPQCdfHrshB2DZ5isYtJkHTxgv0JAiclgq6qdTGhs5g9aLjrJjlDxA/Tj0Y
NZxfIIsymOEZDjVHxEUA8GI+qchIdsz8kdFl/yUdzWywi65wNycz1gMx59UF25HPWcMj0HRhEIxg
fnUplAqk/hV440mJOiKlz4UEVLuJFJq+AT35CyBv1sA/4Q4kh3jOg2rUEj1mx0+EiC2nqDCU1xEP
y0/QeMrmpo8Stf8B8//dlU2m1ZI8yDbjJ0Q4johizC71o8XUenHUnPJrEgn1MRqPWTzcbzEbGsEi
lu6+IJQEVzbqAFWlmq9t8G4M7XtvTL1sb/Lp8FwRH38kS4lcgq7b5T3GuLOvzYS/yNGOR8DINDTW
/F31QHCZ9VbW/GYkYIuDjZF2dBqroYfMoQcKHqNP3d/X7icrAjKNerqni5/YuvYF6b7ycFzkTjSc
u6yqgT0m6K7ieVm7UDzKdna0yICp7n6X4nSkhTc/mGV+odVejPxU8efq5T3wWRfUfP1nVaTl3D6D
ufIQanou3SfFfSApal6OjFN+e11n+TYQCT7MJrIsJgKJjfu0epDjyeLDde6XoQ5yeutOf+Ohb0RL
59HhEMgp74aX/Ad8DCxcpJqis1WEPymMkDxWWDx4O/trNmYdaSpdchqP0QsyZ50CLsyKJdbo+3zr
WCi5l10m2w0b//E4bCB0Uv8L1j4XPVwn/swrnu/LNMrlL7X1z1glMdmCoZtUU223rUUreNMYsF6T
t7cdBxZ/Ax3VXJvZ9tqzfvSZGPPQL0mlcRBeIjL4Az+KRxh1fKh3WMRSwbUllSb8yPx3UMYcAFFh
SU02hdOkBrV+ODJjq2gDXqB8cMgxnWBjteNy0f1H4mL6s4kV/Oz4JG2pxSuuwDlZZgEp+eMg5ykg
jLuSDqwb6fAS+5e6Ght/WbDh+6ya5Hq+COZZEa42eA87ebTdyu5J3Qo4/GTCLDM9L5eB9mYCtxzY
zdC3y6jWGh0UhVKlfuC2iJggS3xA9pyDJ9qI02Ul+U/x8wrY7xt4ZAbsxb68pFnqH7AlnNBiSzTh
rkBc6FVpBhjabHsGQF0s3bbC34wXEbq61Ns4D/zjfMfk7T4Tr2MIOjiGgddqYtr76McWTUoskthN
Jt+dh/NV+1Bczk0okssBb25qffKTTjei/rOj5OwC6s1TCUvOmhn0gcHMHVeQWmWxgdJgU32eKpWW
oMxvMncvdQitRCH2x0+tjvdiPfyuvFx1sgHR7VZQOE8tjj9p2Qp4tjsEWBYQQ0GFYeTCeuhG7/Oo
41b+ipCVl7aioKUzACq5VH6t49BdFsuWJCykOUdGn/vPZqA3TcO4L5Q3PDB/biY5bN2L8xhhGjfd
ewFBPw1L9yaTomKRNagrhr13Hd1PUJZ1OTJFB6prYqfy3vLD/RiikgNiuHInv0CoZbp1jdZ1UrG5
qTgK3gGqahS6HtjCHlJFq/CEqkjsf4xCWQIhf/iFHybfkWhqcW+nEEz/6FHTMrxoHjhfEO9rTW2p
9QK5KaWeX5/LFKet8NM4FPn9aMayt2D5bQiBNyS37fFCW98Bf87X3dEtAr4WQQ3jnUr/x7KJQzpj
oh5fnJkeHN277En2vWQnvgWDPur+21v4Jan1C5mRqN116vPcUvmpFhdJgfH9YCIfYGzCk8O8Ws7c
z/y4x0usS/cryc98BYhtUeyKqD8L88YwGUmVtbK5KZhcWkRnBeBkm9ZZLiaVfv3ipVAvzDnN6UMs
rG+xK9WbDTd1K9JtpZMYw6bW7rBZk8zLhBEPeVBkaqDscFUtF1JVswnvMXmovOnkj6X/TOHrMIv+
DZ0x6N/NRaUA8ndJcMqn68LnX8ukJTJP7cZxk412zqWhmwFnkY0hfP0Hng9B70F1I2EWI3iKwK0f
f+YHwK8VdUj5ZdTJKapTy4L90mAeDvMrDheAAEW8RD49+COMuL2Gj3K329zwQmaTcxa7xC51N9KJ
ER1emWEVG3bvIOk3q0YAJryzId5qR4XHoonnzwRNuur8oQ70yp0qhYyxsVJxWbNBJNnQSMy6XsWw
P60DRFXl8qFdMHcj8TUlVRImFErDS+GuIZjI18ZggFrkKauo7cgBozi97GHHnGCPR9DXYdwbsc19
MzRoKi9XQ29+YzmmbINq/gemsJyjL2Er4Saabjxhd4RV4CXZqZ30R3RB19umPOZEBmVOtqvMnuFX
VGf5JOyIaIz4dPBjAv2bLDovyPk2q5xc0IWLlNq3jfvVyrR0YVVbLAbtJXmVJckFaKca/+uWwF/d
0NPE5TuT3uYlr8zQYmZYTLrpLMSJZzZgnjETWlVXh99eI6dyg1th4y4uh9KLv8891SFtf4mUlpo9
mcYUBH3R7KQ0PkGMrBaUuJO7b4L32tE5Z3Hwzuhq1AEeUmOHhWOqLk3b8YjDM6U71XA4g4FWm9PH
vYRdKEgddmBowUKZdxU5xNCoLdQYaSLWNMixkqsHjuIOR4cctzOMYe7WqODQ2DtNihRrRSmKL+Pq
BsWppVVgCRfl1n7NSfi9q7wG04EEekpyR/U/xHq2iRTrmIa1CPM7UhB/kzyrDnBN71t24xOh4Io4
ebTokPuajdaYJOwFwhh25d/MYw8y8wZtYbv9Fyeuw8NHnEA/hysgSrVPCHktCKIWihFB/xwCLKcM
QrHEtji3xtsjh/UrJ897QJlWDs8H5huhtfVtHx5DmJLr/OBgqCWA8+nVkRDNJbMw7vjZKw5Rxuyu
GI6IZpQIICcIOf0HtsIr2343bIUkXvVFfT2fgxRIQUMmDPWcTlXJKly5Ndj5136QrKijDnBkAEQs
1s9Z1alF6FyXNXefsrYcv/x+q+0EVrv8N0GhdgMEu2dPa9BhwvzhiXlNnunHCbejj5Vh3cjGP/q+
7y/eS+mYfrxhXo94hLeFMgGP0eQwWttw9yaBGqdhH67tfaY/oga8S3KOVNmnxE7dr0Y6C+L4MySw
NPMs+TVT36mQ662XjRRwnJivOmNbCi/ItfqVxJnCK4UtGXDsx32l5+YZSAMFSGEopRadFOxhHLhe
DpwluukKqJR5yOX1+2w+qsdSs+nTSyc/OjEy+dk+s1pmNSv/vRPXBX7XznbXCAooE/bqK3Y29Av7
ifyxKetAH3db3yqEqNomQBzbz+f15NuKpzxvGn195fyXnj2f+VKVniTiwABGV3Q4nR2jpRmDymSY
7+ByTQtPDfJewzOn226YgbTeHtdtrRoMaEj93l8srtSekImJuNjRsXo8/AsH9tQnRY8nsbXAxv+i
r40z+PhG0UnmxMHXgt99ZhV518MMTcKiXpsr8GBz/PbOSGscdUJ4nRBnGOBsFBj8j9An/dP49CB2
tzDXxzAG2kNx0SgQuRs2+kc2Kiev0XTm82lq9KeDzVgJNuZ7+zeRM/CuVS8G5yTtIdB9GnnjI0nP
JPwylhTZ4cVK7MOqo3+r7htBdSQCMm3KhzV7zpScVUeFoClH2WCf954KxuYe5AaDlNV+0/RkYxof
Hss04tMyloGNS7hOgSjaKxMQGkl/SaKhkfNBnzqfpn2OfCnDk4/BkyyGznvmSORXxC4Gln8Aa4JD
a61UeKUMI7gX6nWKKy0w9BdCuXGfrNXZQcFUETPlNAKKMeflpeO5T5G7F16LWQ9ZyRVR1ZKGiG+T
yvzKLmZ+hofJGTgzX8ZO8uP/ToC2DqBfdKiSXHf7eCjz6/YQIVk50PGiaSKrM3O3OKHXze6Zu5G4
7KTJskV2ZQOg+AJ07STFDqwb3EKZSJLhnXp7TvQjlV7LnDcPqdoSSMYsx492mEbC2VDmxA5mQT8I
wJWnl/wMDADub6AFjcVQq6xa7SsDaCpBYZDet1qH2/DPe1mJE7WEsI1pzXsYw8vrR0VQhWeWLz+l
ExKdikX/QKzLdhjxfy0GOTUj5Oisqmp7MG+2CB300oAYFWWpMCSSAumLRxYfMSxa7nPLh0mTSkps
YVecuQG9zkhdFHfAIVuOdSEasiX1PIbRpb61/uV6XnZ2YwIPZDG16Tgcc2VT2m4vj8ZZoARFRNhW
BxGtPsYS5W02scADUlRXE32Io+c61ozVNs6iapLQjWQE00R+G7IZyXzMO2tmay9nhrLnIxujRWYU
+7ewgkGOI8HlFeMC62lYTur7xY8G/XaWiYaGdTJwZ4TH2ZkSsBwBKxzAi1y0rePC6BsMEAzln+XR
yOhywi83mHCrqItLdZT1DWEaBbVHEINe630t7z59w7mKhngdSpDzT4zRKpVg8CV6/tWyXuH7DgIP
5rClAkLMu0TiWCM1SGrp1hE9h8LZRxENz7LBR0KnSAIuclqtgYtFnIZGM2h96qzztpz14FpNf6rU
zPAg7hc9jfeBfPGJ/0u9bwE7SgFjOKsaOIAl0IGZgxjRzBjgBpnWU0XbY2TQuQjyrge7PKBcVSlY
8enNZPZZi9/gHLGnh/5/1E8RRZ60HCD7fGk3YMZOAsgXRD2krtJC8AZHwjj3b9FQh//jYLGNRn4h
PvhtdVQgoIHwqbVbxdZps6+CHlPj7nOpGrfU87LaKVBTJQdkpO0Izch+4CzSC6etsx2VM4tWM+tK
CTZ/xy6Xvw7yZBD3InDrHU27bJRUrdzfDrHcrIK2wFGBuJ2IZV6l769feixhjBP4kUkdXEiXK8+l
4qETBvVtyqRfjVPlb4lTIeNFLiUJUyz/MM6A+2jVRDnf54ND5yfknp4lrD/DVCd1CFmlrS5Frnv7
1XOM14PGhrY2lSCx2s9RrC6dF5NhuulkR9qBKcsp+4yt5s+0KHdPROkCSdbARfP10wp52IvH2jpJ
Ky6/U9sNP8zBqDEZRhUH60/7kChOjM8LuW1FdDx69ubITnEUAVM2TgBgCDxK+Pz3kJn1zA6H0KTR
qP/jA1ZTM4444w/yzxmlr6t0EBF4j4gmi50EO+j2WHGHsKlsPHwgk66pQxF4B7fh3z7mun4zxV1k
VwLmqodcfhifDw1cgUrCn3WVGIXm+u1Z0PksJNdvIX2vykOl3qr7hXyfazda5HvpJPvSmGUGhg2Y
PzFQ7RyXYj14ldceeaZKyJNzgRImwdZCF9hGjZ9SB0l7ePK2r/7nbLkNNkwYa4FJAn/DbrWxhELT
XZRL+ANQ7meJf9VGzCrRQZqyVHj76T4ji9Vt2x4wsOd7SNOzaHY64NYwkQllEc6pg370AdkpwTUx
Thy2VjIXQMwbpW75DVq7QPSrPeQBQ3dgLMGrr9mQ8t3cee1v/fNee98aE+fjRfyXj9cBhSwrdmBy
Fmx2hTKr0g2x+ujqU2eWX6+npPemDpnwcuUtaHJ9ZwODY5e+CySl/rFo+7dCA9L5gK4XDeuiNPQu
0C9vANgarnRcUB2M2W3g72/6sjguILgwgaHxcAZsU4I8P13dxhfuT97LdXl904T12lt2pxuY8Get
qRZKK7CfTW9G4EchX0Lw8m5UHfJ7YHpuv9PlL1Y59mPHpuDYjxsWfQa4znbeVdNNyMBatloON5C2
DV6mvCFcWhpBEn0/nPt4Q921S2pTBspYIX8bz0MSoZDUCyn88qvAxMtHWqSFiX5K5ijevaCz0/Mw
EA90KjEd4xlpMuwUyIRgWI/C/wBos/hP2xngh6xQPUfvBhCwZLvvIvGplaPu59yxDkY7HZ0tIsML
J+SSKjs39TJUchOnDnbVQCtll3+EZ6U3ap4aSiN4ZQ6bezLtBDLXJodUBZDfH2OdHkReSBn6vcfN
hznREQdXjhRGqYNos7fLDflfgj4xI/JB0FcYqTdCB6LGmy8v5bxM//dJB2ZtKVM4NHn3uy6hsRG2
L1ARH0AbnL7Zzq9Q1kmOjdp+BNjlESZY5PpABsQ88+6Xjrx+rpq1GGiSvQir+qDmr9G8MFUuUafr
GWTS6DJpDCRcGnuVyt7bVinqGIu4PvmNs5yHwZbzo5oxEQLCmK6MfTNPaKxoPOPCjMlO3cuk2CME
YpIQrTcEjF54rWyFuEh2uUQgBI+l8ww+Cl8AIPRfSCnezpdS1TeY+74zjp6vYjfpwYci0ffjLl//
8U6ICToHbkKoCtJTRPxoz6Nt5dvG52Vcl62XEQfMubp3PP8Vy4Hx7/g/X1aPg7Dwx9sQCuunk+iH
BV1/wvrXn4B6/ccCRTSWJF7ZiqDTeUNyJrVs9Xszk5uMT94diGZyrABckLMyJbHJ+9ailwgOhhdY
V9ZlnTHqdrU//emxVPhFP0N262+AXFAt9a6cZavdFvhKJYRI+4ZszfiJmdI6s7NVJyK9+73L7d3a
i3hE/0WpURjhWvhJwKRA+ffr9fo8H8i6ybQN7/zmLueAD9ToFIVJoE9qs8W5y6Aw1qdXsOWN4VvH
Tevhry9+J/eOXN+t2dJby4WcWxjPwe7T/r8weo8pudUQBYOSRGYX+8s7Brno60W2TwvTz6UqpRHj
qSnz9Grn5icWn09Bbh2mcKuA/b6wq73LxgX8OyDg4hrlBfC8GhEybZ4brCAlCQxdUCN/sc2J3jJe
+yZUITWs1B3Y/hwP1wOIAlRyXXGtgGJZZ65g8X1Id3Qa+qS5kW8lmPjdlWvIb03yajlFFx3v/S32
aKjE8hJ40L3J4mnpw9+BXVdJTXuPg7JF1KTf9hcfylJ8pwVh+WyRGlhDJ96jEK9toFEBF2ZweBXF
N43p897m5Q7Ff9AJGew9arTrQXNrEbk4roi/u/EQxK1zXUhxahsonOI9Ukr83AbbC1R2tfY2/EiY
YwnmQyg44g2f9GNlXf0GMK15in+zgPQ8ZaKbz5hwxQN/E7BjXTdLUEloDTqaxxQLV2kRz66FObHv
BRb0zsTidYPovwv0XP2kEZifxYTrPUEmgHKKZx7xb1bAhqHSKcqauzZs4+rdiLW7WvjZrCTtMwj4
qX5jLLSIDPdzTpcdtN/55tcWUjD4X99dJRqVnPM2T0pcj4KIm+ZrzJj8rUrQLXJuQ399cHt1soN1
IMwa3sds/by6ZgjPqqhYl5kZhReO/WZn08KMn8uaWZuF1FOVFaEyRsigNTYARsnhbyEtGHQtdnaE
7JnMe+W1e2cvvIr9nekuEx7h0eb2Go0TTwTKE5VEjeyVBTgwJ9leIEqd1il5XuqHUSpd6StxHcBu
qw8O4nqv3GU0U4RejgaCwjLgR378DQk607PtYvnUs5Ik88ETOTmlOuH9Vzw/gUuXVBftcx0OcBbG
tC9KWkyINOqXc81IciWwsKruLhyU4REwIIe2pZ1C3HGy++jZmAcP6bAHrapw/bVJg+QfpFG1Q+Qy
/PZQIIjUfhWIoYNnNotDYrzpAgsNdaU0Yelif4JbJu3o/Q2dI4jK/tt4XoRrhUjST1BYIfYghgLr
6GOq6xvY83hngeiG/Zqm3l7WRr78Cz4WfJT6qgUIqHEL3ekY6xVG6fc5arX6E2MMY8gj4LmSaNxo
CHOCQVMwapwc1E7Rgc6FTq0Nlsp0xTD993AN13WW2N1LEOxAgrsK70yvC+lnABJhwzniTUWFIzOY
AWzBsIRZhT7BkAEufz5kcsfl1+IX/X0Nr7qRQZ4BVxm7cbChDhrx0bZOolpbdjqkGs39mpW0uJig
mrvPin8/vZ0MAnvPFdZiDz83MkCEJJJPdciuFQk6YeqT0YnSz347Yg11d1izMGC7twoh/LWIOEUI
sg25X19pTgfDVXEpneIYh4fjVqPCKkWVVxNxAZRIN+A9tKPPYsbBtCj1kwRq8lpW1Hl8ibsdqwF2
j0JU3yhXJbU9lVSeowChSBG6SPSJoscYwhXkItkIC7x5xCuRyRaYcKC02NgFFbJZW0WUlnw70eK5
HouPO1WCbMIWhy/s711nJvahJFUrpwG/SPzvq1l90bvNBTiy79FagAFcrUDkiSUMuk33g8K6eodS
OgPoQRemQKECc383L3/1imiIYvd68Lz7zAWdGsuNOK+9pDX+SmCTfx+Iz4am7LbVUi5D5rJ8DxHY
1jCtZVTDO4TEUmGRn8a5V/OQigAM82iDo7OQOurui6nbgE/8JO5qaUreG3HngfbkLh4KmHqXEnz/
oe3f1kg1bHElHE0c9WwL68zsMVIFOSr0EeHCYzaBYi/UMXr1mw/ol6PZAPUIvX7naOzgMts2J7cH
3O6kOU4u773Eoe3D/sUbjFnzxImcKUyEVN+J7UBp2Nq1cA//SsLfXCJCtwYpTnGJp+8sgJABMrAl
7S0DIyxKBLtZsxQBZuTZO/sVLegnvAAUH6HXEt9m/+CdjrjD1mV7xNF2BW9BcIWXfVZAMlB4L4gd
n7ZZigDpSWAbtF34ZCwlv52X10bk0NG+s1Re/MvM5D9twdIpScoOeA4idLG97dwzr39Uxya51a6z
LNBh3gXC3wfQCaIODFhouNM4nSIqGUYNJSg0f5ZX3WM4m8FAuSnzU2u8mny3VTBP6ZZb4OKyea0m
NR3lnn0/NkLOTz7xsAttFkB1Vd+aQjoyZ69HsT+OI6be64bMGG6gVG3tgjPjZo/DscRye6XnQX3K
6yHJan1niuMzs5G4usy888tSgi3KJigdGtRB0FGKuZMo1cks5xUQDPZBeDIktb0cAd15Cs4TSH1B
L4mUSwPr9zfhE8cAXB3pTQetMQFToj68KWqh14XzAfXxv4EC2cuSXQgqOhefeg6BEC7SG/bWEk+w
+UGcbGLhSS3HaTj4oqvHwiUle6wfBxMBc4XUpfZKgvAg8JbQFWQw7UZUgPLKif2V2qVIKE6lqoER
2+j2Nbn0+C9XG9/ALtjcdfVET8SFX4Ol8z8xs2qh7RHcqOUnG7r8AEV7sYLaDokYBP7hnQB4VNd7
8RU1kizGOfgytz+gWD1bRtxTHbL53u7qAUNJc45KymFqGN4ddjxHUn4HViRTUGkj90PXekkCFdPw
82ghCT6PI1vgQFhC8P8MhPNmJLX7nXO9ZGyt3v36f8c/EBQonFt5zK9NlDLQQtFiTe7CVVdbS7yg
r5N1rcKwhRd11p7XoLoqajt9ilev4ZqlIJcToFeeaEAzzia5YIWA3XwtRsZZSzA6ggrwXF7a/g9v
xFzLs2xkD+Mi84INi1Y6Fi3QXUiOH8DG1V7NhlWB5GWNbwku/4bDLVdmrU7ZW9XmX6RGAhwZNDLX
faVkrtxp/8y8LwEqbDjUNyVQZUbi+fy9q2uR8YUBk5ca+sqjcWQbtKQ46hUexaF+MUazpdYhdP32
ef6PBg2Ui707bVUMOqMbXeh4v9jBzAaLdiQakQyXJZTPfFsoNak/c/KUb7aQh9YQGWb3XL77paOg
0XznWO+waNKONNq2dSbSmkGFXbAqFNOsAcWNmPeaH8D6PmC2hjnJZ4CGU8ahLuBoL9qT42vqAh5Y
E3MrK6CJh9mzHos/v4lnSqeijXPm5yBRcW+Y/q1b/gsgZx//jFZU06mFrsWoZazQYpWT3XlGL+VT
ObpzoMbPpvME1K4Kbhsh8MyZIneCDj6q5m/rueRCOC3/pUf1Qw41utaXSzZr6adDACn9KSxa78mz
l+zovRbfCz9FJsLrDvCiWkcuCjjQ3zv8X/DTLs8181wu2ygLvUQK1sFjFvTDOOdNO9ovog5z/d8b
TQSIgFn6ybEvjT6xa1W56jqKkZcH2QEQwrrSHxsRFDPcJC6oxVKsmJO2y7yB5fMIWObChqYpMth0
5Kb0tGeDZ00jyCnwbaaRmuO+8wpZGCl89vwe1cj2xudb++LJchL8oXlitzuGmbxQqWp3R9WMPh2W
oZUBFD60JA0ufl8hjniFwCiEBZf839s3RP91dZGoMeZ4tbSEHhGiysP7HCs2jFwG7+GfiHkHBHQx
FzIYOxafPuVlNYY87wUXVhy16+9e+q/2EaqZ8ZlJsVxnuhaJcZnfHUMrLGfFSK59ZONHb3o4vjBD
S1PY9RhJ9jqKfLBTWSMk0/SzFxtXP07vjgGLnUyCs9N/P/AQVDcLLoncabuN4EKqJKy6jCH4ORoD
cUUA8cs7VkqLCWSQYy/Nlway1iCIHoZaI6CCBGU/VEn7djtNGpcqy/49NBhtxXU7E41BCqc8izWP
LMV399iRQRtcGNb1jBIqTivIcCfP3Ax12/+MCzdCkWl8vm1H6IrCZyuv321P2V2IS8SjXMHUZMgx
KzE9RQRhLPXXC4LMHqR9e+BSeiFFvMeZ2lfDIS4X8IQ5JSt2GKjilacGojzcUXiCiBJIBXe+2ryE
ktJraoTpKzSd3G9xeW55pd78H7DGtC0u6KnFbCyCMCwSa83/xyhatQQZQP2/ptozfv2CtyKo/gYE
gSfoGSIbugdy0jrxccoW8qyKJsZLoCNq4El1GgXFjMvZfQCJkSxhz8LjR38Jxg2cHoQ+dTF6IwVr
OaB0l15s3irMiHTZWZpLZNGYN27hgvYJ2vImY0mZ4QVJUgKbgWb+5laGZfRSKqukwu8x8vni4NGf
7x1XEDKwasObzomthzoLh9bNYhZjO53Bi4N/jNO7PI4SPS150npKzMHFEfZwfE18O+PePpMoBcmB
DCSh7OI70TSKgvio3OthSD7L8MuCADemcRgbXLFBRvZleHS+Hif+KHQteQ0clrTN0hfRtgVw2dS8
lrohXkLjrYGQS+u/hMFVp73FDmKpbgJby4UXGbuzBe2y5Y9SyWgcpn+Ewsv9ZE7A7ouLCnMAp1Yb
qyAMQTEj85Rihq3OO54YBLwqAUVjY1UOcli/AWrK9Xqk/iuw+RGQvnDtJULOlnXHxkiI+5IZ/uoK
m0lA1luYMGOkmk+fUCyele66/3cEFzcYAwnCLaTiPo0gxRUlPO9AaNvikH6gkJfVh6+Jg/FiWlHp
BkYzWZWzvj/7GQA2nuHsqcT61jZEGMq0Lmt7u+sI5Gbus6TTPT8hYYAB4JyDSbdOhybYcnCI4+Wq
QJ+izF0/6wTDA1KY7glU9VZVNeaT2P2jbym8WJRGwoqIhRBxLhTJ+XTxOwlMU8mo+SioUP2eUMRK
bCnAZzm2sxZIKTQcs5/dJjbKibOtRkfKEqHbuEWVUcbJEwPeolkEK1hu+7SOO0cVDEzqk5YGZxun
onMHBDrLiaG9z5qZa/48yyMFTGt7HuBW09wUJz2Tf19bxO0YJRNQPiloxRV1leZ+pdnYRBKaU4Cp
Rd2qqGX9kED6rjc/4lmWraTkn+2vZKok3FmpK/8weonXoHcscaTiKHml+mk9fBHuoVqItWH1LymC
W3LBCvL6CYqch3nVEXFA2WQ5Sf05DerBIGsVUizjOo1aIOmqS/Y77iL/woTnWrcqhAnmKY/Rpi7V
GG30NTzWlfqMxgSG+lZ5VkD08tFupKUJDC2q2pd2XU5KittiH3Smg2Fc/sW6zPlBHC/ggh7vP49N
R2NIvZYmxPXy/N2WhOIr6HROY9Bp0xkY8nSdHR6GHSQtZrgQwhvBq7zU3EivPvbl0E1pu7XCdC57
cP7yV80WA0/W/Gb48+33CFmnIrDInumRrBuOzg/94SjuDA0eEvIoE2bXsbfMxjfdf00wjidY+jgf
6TrHH/4Aa2rEraIgfsKR8vrVYbL01MVvD0p5rg7J6EmTsszAWCVktCF6YiZMU4zja7QFuwKjjQcd
/tGSUtHyC+vaw1dOvLSokAGmsY+HWxdzlE0V1OJ+TaeAgwk1cKp3wngJnjQNeEnB39fyFRyWqpv/
i3kYM9udqfvCJ7kruf2TrppZPUxSY9Zc4+e18KkeHLQLrZb5+oA1loWxwx3G5AaC002kiGBd9euZ
92xHL+HQD/oz72kSLiC2PIJFvgYuiymemWscu2SCywJNJEAAXR0tIkYMC6Nx+ITlWX+UxW9dbUh2
M7qoEtkuJRvPCT7ImxZV75dIqvZk98CVhPj4kZ9r81fBd/6ffHbvRKDU2sKkMxMRS5uUCSIZO8vb
9n/92KAF5Q8MQ5QyxaTQKa6IPQ5WWAFygxWK4OCaxH1c6vOkjOT3IWCydK/vd4W/J65CgumOo5qb
xgBwMaljpnLH4mql+wu/avYmGJQh5/vT3kka+KLS9hlWGCS8JlnRVXsZ8OFdSwu5CH2E4ajFm7L+
drEYeMZU1hP1s7Gt7MF1/SxbBh0hk2RbNwnEpfUBSvL0ena3BsO6HLVssYGpLXzANhzBa1+OeT/V
jA+fURuvE+6rNq8N+Kb9biISm/JFooIyHG4l17FdhebXuOuI7neGouAzbLFe1BlpVSZUBRgKr0TM
7zZkZ10KEZOcjvtyyMpyR8wNl3t+qD3qI7cxGDkY7IGbSwpusG15NeY85oh7EFahRSfS7TWj2OOw
TCV5L1g2ZxaUgWn+d+LcUNP0fl2oyEJob0pPST7QtH4+tqfXaCydEGUavNCKOp1sscU8MV6rBkVg
4oYBG4u3ASCAEogwskqEsO4ZOB3jMDSMJjDKWDayWkp24UeB3zXbABEGEyE3gLokJV+xMGbgdfCj
uFJ2NaPOV34NVHVBkRI+uRNbuFUYdqkDm1kQFqOtoMZXKvEWhhIGiTgPq4wVoZbd0YhbB4d/+Nd8
j5q2jR69Hrp846lcb/6yh3plmJURnzTe9deuicKTvJr0+bENf3EMg6LlNfwhIxPc+37mFAZXsxIy
jSvWdy6PUf50ILtYpTgqaxUDjk4fc03LYU/bPUD1BAmz4fYVTQ8mnkmFBIRmi7sQZTO0XMwUEU1j
w0RbOYVfy/DxK1N+0by5QcxFhPsAwq3bcIPuE/1wdj8OhaGuV1x/G6CfcFzxLdzyVJmr28n3qVSx
bAGtz8lBRw2tdz0pOKxAdgsH+LunjG2KkrOVHJsmHhmDIHNdnadKTMk0NaxLKc0HlHxBoK6yWr3Q
YwI1UbWhHaoXEqsldeL+BRVSAzSlknSCf6S0DUzmGWB309HprqLjGhwz9gP1ahquMU556KmGikSV
pkcQxoOAierG4ujmUKKwgh3+GEoown2qLwisnHApJcekcsKoZsAlSN26KEE3YjBGPCjSmeus7NEm
3wxofyGpORs7f494HYE0XcQ20fv+4WfxxO/2+u1I1e2+m8QCD8z3Hs8XqeXSvkE2uYGu70ra4x4X
vNYlarvGkXVKLp18iZM+AISjvkUEFE/Xnyp0gORuE+NunCzQiu2NLyCO0t/kU0VgwLRQit/WWZXj
KYgRm4LWivOI7jTM/0ZjaRBA3fY6naclYJuOPLh+I5ldNp0dtwrILSAamIl+maZmn2QfIRGP1DV7
H3JgKU4jxaHpcUdtvC2HeQWpsjIGpgC39azeULnNTOcd/AAHi8+sSehcrfnBlbAEalRKIjgShgWj
UtBkBlKqrrLfz6dXV7aFWm0Xw025629w5i8BWaDK3QtT2t+MuQGQF4egsIUCc+rbNV5ZXSjDgh3z
EeUNIrRf2xc4oi1EmklHD6PrxVvAQ31e3sH7ry7CxflZBVSBKiVLbmcFo33btpGIwnuXLZM/Cxjq
a5vJTHOYHjUi0dpOBY//4JdHpFhqKGxH9/wkXAwrLvduXh8QceTtPYHztDN9BaGtQoQrM+5JAkxz
xc5Trjc2jXzPVcSDyVT2yDmSqMOBEJoF7c1RxEp9v5Eb0IE6kHYwDkg5Vm76Ns7nsDP0N0PGy4pK
cN7WZjlAHoKfu8DGl3/gPdXzZOy8mUgMxlLCqxsJ4+G1ej6gRndg9zgWz5oICAnYTo1XsK9dWAKO
jn4vmjd7/gbQqg6wFxHjFXMNim+M9bErAIa4WE15j0USD9O/rlxYszRolSm0rSjkKB+9lzqAEc85
navQ9w47U6eFPGqOSX7nagwP4BNWvDHMgU85634GKKZ0XLEun8wGWg6iQah5NEkQINEJcW7gzxJe
qYAAoOeXBT94rlCO/JKUw6LySZmgDD0pifc2Xsj1pjL5Afo1753FokWOm1q7DoIu7Jgh7dPgJ19A
mqsskGXYiUg+GefRh3PPBIL6Lt2RPxAit5IYxP+Paqv8dWHU2AiF7t1+lXTZKOIavycZKfXP2W/T
7MRiyCfEQumXTpw706Ab9t94Qx/u04PP6Jt8eAsZpvhOWW1rrZyFu2u6rMBosRPGmh0CxO3kmjhj
Ww1K5aRX0/JXznaUWCxqX0W3irgZ2Uqsdeut0SlvX2CdH1czIlSTQUMJe03bS3DmGk6Luz9AnSFo
8NbNTf5+nx3K/coYN8hKG8v9BJduDHmCiMc3N/zMGC5zj5X3fe3X5HO15zkdhvOcKItvraGTytgm
oStxxF2k9sFZQywjgG0/X0HDt4sHt2veNkiC8zg/Zswem2Zto3GrWBTEyHsb6rKBxC5hYWNi5l1t
wIBTv+qMTjVo5uyQZZ05ppIHdwqR2NmgcAUjNIrq7lDqOVBpn0o4XmOK8EQVhroQYLLJr85qacF1
wJtuGdiN9uiO2PrXDnav2p4edsSw+C0ClR+6U1i1xBKdHz8xJZhoM7odYeGVkc2WQ4UdRqR+cE2a
l6kHkBAChebgmCggfDmOth+lfEKI111fcvGmxheEg0h8K/Az3HTrSqJ3PICbHdjjEkah2YeBTfVh
EfUsR6r5ABXqgh5gL713jX54olQwcVfjfaWDxyHI8/vCCeUvgjnIN2YvpW62P3jjhRSd5IqGhORO
ODh3GkLS1qMbJ1qxV/R1PNiF5/pvRZX3v9d848Z7ejBZDV7lPwGAZad5m/WEdsBPMbarfVsAZSUY
j9j+DA1GcYgGkLuGDomuTVpLXWqx/G6igHRKnHiqOJpnvkV+WRazys93GpPzPv+iFpQowG1kU+eg
ZzlYuazbqTj3pr599+5UGNPlWwGEUpQoiYYx1ZRwABNK4HsYjXCkrXyIzLulM3fAg31SvDtK+dPp
unt5fPUDknNgmyJwNwKrEmLU1BBnXEqmwNryuOCtkCtiiZwxErfJYqLzaRnhF7D4htyB/O2XVaSN
GnH/7GznhTcXTpKApH/+jrKxZaD7eIo7XlpZZE9Zgb/zUbOpF2XoLGeOw7MWMmlZogJ6OF3Wo7PI
qVIEBojSJnxx4TrpboLgRDlKFUuuQGllXOXdnfdIs4ATDyBECY7F48nuipcXPAmaztSoLMlmtmaX
8V64MGS3zs7pI9c6Qxu7FX+eTwY09e8v4sFAYrNJRx0RgxRY5q25NnOax1b7svd0m0DapvnKVN7H
gQcGN+HJjqnQV/kmAXJ2MwVg7vnvKsbNW3n71TbrjXQgVL50Y1NH65Be3neACe4QHs0SWTkClLbv
sIixdFogghp6ZkTu5uOBUY4o4t4Ir64oGOMocwY7ln26wgXZsRHaBzEV4qj2MmAZmGk/JD6BH09W
tfToKoKb5Y0HJxD5Om7OkeYknKyfDSiHG4HD+6p9/UU4cKwrpoPGnXAzdpp5JxxItsHw1ANw3dA8
VjKui0xgUC5WfIzyUn97TEUE2WT9vWqqGd1acQHAHVn2G2BwXM0ZJifmECDxglJZ1NazfRp3DoQW
Jw7UdrTDbx6BALzHoN5Uv3FYy7hE1pYPlwq0+X2mHA0++qK1Y9WtMU2xv9hFZJLzaHIz8s9vZnOV
4t3PSlkzr3z68Mbh+M22HPimLobfjldlqA3RLNq9EjTlZFsO4AeBGWcA3mAoMIUSxUhHQb4YYw0Y
q0ja9R/MrimJcN9S16BU5TM44hIbIZaJYZ0PYO3zHZ+9eqGUzJwRrx1to0W1QYax5Y1XaoCBHLLi
noa6aY9fskU2N51+TUJ3vJrElr2dS69+EInCfoDBq9+sY0fHAMUPM3ugLUkku0CHOgl5yHtyZb8j
bkhCeRDC89vtw55v2jRFZfeyV0CacHKp4cOeoRCGVtjrXzVDb21EnHwmR6foaHSmUWrFno5EZgVK
ypekbTCqMmMkmvQf0uff2Fi0a6uFEHkVRXT+d3uhMIDMheN5zdcZ+ai36ihQ9PkAovukNeXEmKtH
YjOIe0m6eUpvvIpIDnjFeJHeIjr8db6cQV7oNkslVTmss5VWLM4+//2aSMqdp7llb5ki+DdwH5X5
VCMG1o/f0fbg/jb9Q++quNaioOHL2OCvaJuYNNX4yMTtKnNPKjEpNoDvkXE9T/3TKgmUW2rh0DPa
cvJor56iG2MNWjgT+FTWNvP1dB1sWpEuuRXY1eWdDiP0vxvZ/J4izmRJcSFFnyxfQuXgF9CzPWQ/
KH0fqeVRh4+aOe5Iw3dof0tfWkF62TaekSbhvxLvFtyMc1WxJuYPKA3ZkZAvt5JKWVYHJhGRMLr5
IwULgZgyhJ/YAYoVfnUcnh8T4idv4+JCNv8pyZ8pJzouTSGSOfi//pkacfPT2Z0E6FlL6uHFAMwm
duwqGzPrP3VL/O4UXL1D8k1dO+NyaZIAmglN1IcsbL0duTu9nP9jclrhx7UkG1uqgsuknnETD0P1
2tGQ2e4dRcMQTFXlIaobrdaB3iYWK32n57ETFFDLMH5mN0g0Ufym4tqu5xpzw/o8DxJV0IqfbhlI
sKtCCNO1VvubsHLpP74WaqmXK/cA0J7detNwriADNztXw6HDsSPgdKuAWRGMBBFxfgBeSla0Ki41
0nacSbEN0pfkk6fuIbB3QMBP4RuUfJ8+4aDprMMa4wbvSVTzTIHvsGiRcUH64bB9xYMZNcvX/z4S
panffjKWcnqJKreEG9Ky0rgKUllvX8td0xuV7G26ik7QDKpbhCZ4xis/GJh57h7YGsrmjhy1zcDI
jnqqxx6efiLdKTA7RT7NCa8/ZM/8jjji10LZFK+7jaCDuitDyBmgKA0MeZOnTLOt6D/DF8EX+TS+
HusZejQkI3F0Me+6cgpOyBvWdzz6rSmavs5lEFtCeK30LPSmZYamYVW/jWeLgOu07GIsQ0fjjLNE
v0YsRy6ibChVP3b6nvfct71VtvMOlHC6GP+J14JBD/HEjCgJFKrjfysvpUGq0iLUaBgg5vGhMz5z
q0GO9cC2vHzjgYIH1DF9JzII/C8CuGZUg8z+ML5e9bWnB9fqUk2j1nrXOHoRTKY1mXMA9ihQ8ZOK
CTFwl/LPpImvWMbhFRj97HYrVoUeblZyoGUNKEPsRvRWfpH3Yc5l98FY7jjtBodlaFEzv/pJtEIS
mEWSRskOjfIGaAumn4DmGSC24oS2rfd8IcKfhvfqgFiqxJKNpmLgoyUgppynvO4xVtIN9JbIsr53
/AYpqgAmpGoGfSx+JoMXnUQBtf8vd+OtFvP/wTTEkj2U5VC58FvJyJbhMVBX7mwJzFyK0TkMUf9x
myEO7VcG/aC68+PkvlS2sxvpt8CCF/+zCFxsR/zNhYp80FDWg+p0kpYt2VBRYW9yV+vLFm7koxWW
xNiyDXchX+wjTT3ybX2RcK5PMNB5ISTo9rMU9QY4DaAj5tCQbZP+vN8zMpBH9FI1NnXGHKXaqz5F
IVP6ISdoiRcz5cZnSBpnG14HW+x7XKGFt5Z6Ygiw1myY+bvoEXTSHOUkQkOjeLmkVk4nJqbccfkE
L7gvqywmreglaf5YcwsgqLNKnJ4BgWrSqZBLhokX/zVYXkOkXuYXU+A/sFkP24I8LxPCU+Gt3blj
fRuzOMUVAOVvayCEoCBtqgXo/UXyMhy106xZmUEBRSv21n+/jcV6qQeWx4HvVWIaMP2FmQwMEogu
hXHxanULjInBoTL+huaqCqBp1awUsKeGY8Umm/cfVuq6AigY2ArmQYGPbaTF2OYqYnw9/xN0TRCP
WwQIAI8PvXUt81hI6ycG46YlnJJMGx6VOmT17mkIIuy+ZRrfv82wqKkvoOP9OAf/yTu19EJ0JpOM
zCfyNCJdf14YlwWBeq3wUdHSGgMmnQkMkgby7XzfynjBBLGKhdgqs4wsfuyu9bRwCEhiDEWLH207
q9wPNZ4Nuy5Z9/FkzpIL5S63yMrCkWeAomEc/U6MpSmwEgGkw1ITe2tL4hmlVvpL8vj/ZSK5V/5r
CVxROim52ZGGUoFvpnH9FNtqZ9udVHdQPlvUaVqsSdo9maGe/L4MinSPIoxecufjwMZ3tI+jZ7Kp
OPGscA254JhKehsajDcHw2d120XV+cnsEsTHmrXsF5DhvCcPo0J0az12b8T2vhQ8P9VOT7qbKeUn
/fmnrraM7FK1zuSTR9z/A+OStShfWh7iin+cD8cM6/3ouTk3geVeY7O2wle6OXMRoIYa56FdzXrB
JpCW9bY99TtkMVmF7I6drlGBATE39caClwX0KgJ5pRiZ9luGcAnJUphVPQPYd0oewglifR9PqsLT
ZKJCpuZHPAN9pNGT87ELgCcKEPBZY16Wjetl0/TyT4hUg8VvqVck0rpcplESCRs+11VgyP2hXVKJ
MSczW/5IftmUm8GFOEXZhA0sDLSFZbusLFP2ZlIF6dp4Jkx6Sro/6su4Xad62oEWG7qLVYJHKON3
9+vYSv8A9XKokNPl8tDwcaHMZANa2myROptsm9Q+V7HZosM5tQwFoZ2AULK5ZL4PjVHEaZbnpbH+
bsmHDpwx6gCRqPQMBxRaVGeOsDzPU9y3CnUER1chW0eiaIZ+K/tp9epspWpy3L8STthYCvu/wdYN
SweBAaKc5z8/ZkLb+kppWrio++mdZBRcfqxX6J2fl6KBPJnoDG59Ug0E56quGRs4IxGjEAiNcv2P
4Rgz5iu4UMnYKX381+mgHSSiPnnuryZYInuRpQNBf3kpM87wQ4kiPDXLsKxFDuFCtdFL/XXHUu1w
s/Uo1i7TSh21ykiTYL0LshQWWEvBrc/Bp8Dj66J2+XdyIHYXUOZOJzTDxFsT/AdpSnMPCHRGgggv
6S1q7ZWJKfBg081rMZP4OvIzvtdwfzekYLJcc2PvHL4kbFKx2p9hDbMCmwcwptDRSGMkbe2Somex
dZpkKCusoZ/W+nK5YdKQnAD+fqCBD6v7bJ5MceVj2VTbTW0XCzVKG5ETh3+LXhG/8zcilhgJBc4V
a7MWuSTkBch0/jhWKHOQwo/WV31JFRM5Og5HD6j23yjzqNZr42Seh0EfiXc8qcc0VyU5BbNpGRHK
fQ5pDIz9zA9f7ST9tdlwDQyni89L96wBWGRaZU3oA4WYYyBZqWipCBYv0U9DXjfrz89r+MiE5+cT
MQBjUd7zeOMtSX0KuyoKDeWcNsFB4O1FPXgh7wIIqOYHSRDY/p35jq6TvUjySaQCoi5Ml55dSdLY
2ZxPgoss3Lt3hw+x5kV/b2EFJrCDNpqRJ4azwh59WFlRXUemDplAdWG8MCFDdF1xONSfcNQu3NlL
XP/gUinWbOfcLh6SoVqUGqj/DX05sbjPDiB1OnR4Ztd3e20rxTdL9dO7tsN2dBkm3rsZY4oZqLtc
liqXeLTgaXNQsiOcWHN636+WRjDAcr3dXGQR7PfDtHUJRPVqAsvJL35FnLEMR5XkaHUWzYJDHloP
X4LLf3xGy35QHGyDthfX5JT38YaskzfMMhQAjXi0tv9X1IQkuFfRoW1Zm7+ZeyhvnuLbo4GF+oQF
fG0uh0yNPOgK6dDMXGD35PY7Bpp7fjzodUxEXxnPWMO94UfU7Wl7YqGuuTLh2DClvDWiZhUVHcZP
cwDXtRR9F7sqaAjas7Vqie1wi6R8X94Wm70SA3WR7LcOYIGEcoB+9081J9aDlVn2jcms9Bb/17Dp
0Ye2Z2XGigBIVwBnASWRBfgtebaBacz0Uc24/VPEihIxorlI3/Rxt4PYgto2HMmweFlghhp61Uuz
hwG9Cxo+Gs4rzOSL32EBvK87PrHYtn5ag5pWbYgpMOa+7BFxjCHiE987l+x+6DvK0E/sQY6MP/Ld
srfnSLe13UL2l4SBem66/ZFYdoMngdAp6mtD1MMBfNxEuapFGW/nWfN9IhWaHPBsq4IHNx3X5wcW
Ijm9dNsI2ZeA43jRkcekz1vv3zlkO8dRw2W71r5++uDeihH8cS1s6z3/YjgHFaLMXf7wj8hCErqg
2UB/SNOjRXEbrN84Ovv54Iy2RELobzkwK8e5vJZ/+fwlItGVVqe25MCx3bRs35dNc5LokSs600wf
ovgAQbMurbHCSczfGLNNaynP4Tja82duMXqQ3x8bL6Aw10oNBXvBxgCI7qu6CmoF+d11foW0PQyd
CGWp5rosc0Z9xdfkC3H0ih3ibHmS/hoPTIyb072CcPB5TPFcepAwN0SVmH7ZdQxGaiS/hsOfk8C4
AbRgV8r8WjeOplZlc68rZQzm00mrDdmJEVNRQ2v6CAp6xSnPDQe+wMI8zHmFpOiRrTp4LrFxCia/
6W00Avv7QJ2s5y8haX8MmO/w0k4FIPdAM+/YnDqEDlUP2SBFCefVRQFd49ACNmuJ16CH0N8kjbDM
ZSI/LkutP8gSkzQawIzFmqMmaYivogeYdUxUpj0SeHRi6ceVNyNZPz/+Y0u6lUCuu/tvynghPnUW
IxGST6KwpuWpW4hb8pbvJ6f/RIpnucWV56Ovp2U/m1TvtI/wH30k8jqt+oc0w5ylRqGILdOzhVuG
s8JDY1nJCPW+YQHoZftzGaebdeGHOEQvPlcqjAZYuUNA5YVZKtI5EQSshQxps7uu+5fFVzR1KYW2
MDGjTkZ5bOuLpvGL6pNow1NK47FqATUMRPsLv1VU6RTLNgYPrpqz+FAyG7ygF5vqlCjrdsUxzdJS
sgq4GWF0CjT8CJWJotOwHu6QtPCAAmeSR39iJa+Vym2F5YlGg+dJP5QcGLr4tOYSgzSXa/H9zno3
7ZkfCltrcyrwH++jCTwRUGBxa3EHL9b5/Nf5wcY4J+4miwT4sRruLDpRWSQQxRy46SRMECnVa32Z
Fb9dHf8Xnk9cZlpBF3IQkqwvY6CMbm/xarl5BI6trvSBi4XW00Mkg75rLcjINZLYJqOdfFE9Y4J/
oDu+zWqWvO0I+rdpxymMpWPoDMkS5uTOsFW329xhYU4VdA8RN1f2QlaunYA8DJXfU3/NJdSEv5JU
iNwg8QWc5vmpdrobg5zsdJSvILerhcjKcuJgCnyqlYxu+9LQFM8XUVs640Plq9/lUcU0ALXR4EXa
EgK3QVVMiCUprHS8ut+dA+echrQ51oQub8wDuChYmF6eEACLpB8YvxYqEpldeT37iZgK2HDnhzKk
DiyB9HguU6ydyUlz66muUaVbBaTRPtM6JHtybDXk5nLyyE/Ourul5ns+jY3VuR4AqzsVCAHzSiDA
3v8HNffiiJFbGM8o8ByUVvTq8Tz2V7amYzT59hy44YEa2MXBdyLw2RDNK1TFirB4xvjnASFtcU1E
xrMQhBbuGhSBmLdnbWfq2nOS2SOeHjuupRwOAIHyaN+P6s2nfLZC6hJ3GVRKMwYG/LvHR6drsVDl
izrysADePll1RGcPY/Oulb7NIS3FngX26eKx3XP7HNRVOjM4ev80v0Fcz/235zk+1e52pGRLdZBv
sBa3voVGZ4AGliDA722vdEv5toUMh24eP5ANSaVGyngWE3+ulwVEkCXuvXkNOzCxAwcqAZbdaOeg
Le3R56QhFZWCOk1pfH1D6I74TAzhEWjZX4DB000iaUGctpbSU8o+wfIOS66o9iHYBzYmS6iBnvzo
UsIqGLHw6pxA+lpnJ2uTDJ1PzBo7XvFI5fgPUSmWyZrG81iLXIlh5NXu1dVEBC+DgDLtZ0WRT57T
f6YMowFzHFMkk1JMtGiUv4/dHyiNK2aVNvX4hA0Smm56JwsQOjQm5S+328iBih4CjcjUKstA2nTs
f+NELmE2qSDGb6PP2vNdaA2rr3y++dMMdVlPCiJEtuNqKlCUKwtyIBudZSSN/C3QTLKySva/RU00
H1AUW/e+Z1DFO6iZuBykUHdiemBxTQ5FukOxSajJC7mLp78szonbcnNgoji/uNqdlKC8TCVnKJAV
UHyBLbZ2hCWh8mo7UK46Ny1UE18TVCE9A2DEmWM0YLCU11h7QF2ROxiBBe3STHbj3oJQlwniaC18
crCJLt5Z9XQ+CzLO2gZHa8BI6SsMQt3wjbKYZ4XLrp63r8jv205AgrVbYH8b4fGKA1UjkZpKAOBJ
9dW4dwlxg7ip+mKyTsJYoykYEsQiSC34qgftO954V2qFSWm1qo3054ssv9wbVV0GyOzn5qMogdP2
huI3Cgcxw8hrPMwWYBR+xpTvoHx+kZ60wIGTDMlYxPbsAO3fYDPyFylFdONelXoGWRfZvcLWnp/5
DJu7qBE3T2cfEi6+MAwsdSiBdwGmHpsnlrQJGoAngolMhmNANGoSjmuBBYOESjlxZSMYVFk8Tu8z
n5gmbbIPXdqwJdlrjz3vYN2PCW5KGPbidSCP/9/muFMwYtr/DJb9nXzpFcdXR00SeJYqzkhIeRLg
h87vTfr660Bp0bRbvMKp2UD7Ya6a0hgFWTwmtS5pqfiX9abPl2Ac2u/kjB53OiNpWpiXAgM8SEqt
MO/0GegpLFDy9277hCZ4xbZMoJ071fIjLoAOb4CbLe1tTXzgADM+riAX+l1DHDOe1ZkNbZjupZk3
JitBjt9AcA40BafRxGGJLvaP0zhSZo223Kyfru2WoYAOAXAlOVN5knai5NG6O9roLeEetcGdAinp
S25lIm81toF3dNWaVbHStQAJpZ9iLwRD2EcgqmcPcbl6i7VSBL0fs5T5a/ZpO5Ko/ku7fsNi6cQb
0bi2ygtiqyw0fHUpiR5XN/M5tja+tuNoJwsBJXx6f8yXPKaU/RhQp+4eTnJl6u924WYG40TDKy2K
zuFkjWUnqTWnjMr5P2amgQcGNfgcC21+tOCjb9s+L5oV9Km4tF6Pin/I7OST8bGzCvn8J6oUqrTe
zAzcAGu6uowR60yM46rZ6CXIErS/+U+IvPnsetAQKUhHpa94gOw92APu7kfgJbOS+wGeYZajqPyc
ZHUQHtFFXYDnCekB6fT9zm2Oh+VCaDMqpG3bIgg4L409SX0hVrL28IyuI37A36EGJQodq/3/BYz9
v/lYIDJFpKC62NSEz5bzdEyz5qvvJOH3jLchCO3dTciEi9bct3ADLvPkgK0SEw7ze6ZAKZrh/vLs
KIi2tV04GVvcpdz44zfK6oVMSMWFW7aeg80NhlbSMhYDsbeOpY1HhJsMXYSdeYn3GHVQxkwsalIr
9echNO+k21wg1gSgOZ+F0r8NETW1EOwIiGdpT112JyVdKa1l77EFJVfoUJT2VdjlJs3qRW+fZD4A
8Fs4M7yhSlOHL7BBtH3ta9QuL/Tq0E2dtsNFTwB2eSFu5XlUG1rHI18NSO/cKM9SgWUXv74eMne/
tO4e/CIF8XGU9BpnuVA1xRx3k/1CG2/u6nWHfE00Z+cT722U4cMZIMtO8I//YqcaEHqDw+dShlY/
cn08EoLRM2Sx7h+/Dy9/lyZzcemwX0N5P7/MQB+I7AtXtVCfrD6Aj1/7bbp+G/J/0y+84Yrgw9Tj
RHHdf2uPRDLdz8QsdLT3PaaSb4VkGSYz3VFZ5Q27bhhC9Mi6sftB8q+9kt2Hkw20Z78JfFeJ3jGt
FNlWyiyrEfAgLJgYpJbF1fmhrevtHFHpQghC4NNtlRv+KzoZXEiP6Pk8jUvYC1RIbQON7sZVfBlj
7BmGq4f18I66wTZjvnfpZyOR1nU+VYEmV+GmDbpk0d4CbkmCTsRjhd5C3BKhU8VteRcS1NOt8hb6
+r+klKUbt6X+qila2jCbdl2wtsdX+2v4WCFFj60ADC/KzRWwXh9JLheaCmbm0XShML/SXTS5qCKD
gIZ72HpbxfkQw4ULctYM5XPEBmftwgdwyxd+PbpQVSyZR8FgJnqUhTG2AdXWI4m4gBXPQdj3VCkm
I0rgzQtt54Lp8IjTFkq3yEpSBkBEHA6mk8L65zfjL8WBN8ld0rZhBLiGgvoRuJjYEPxL45jL4bbD
X931PYI9S5i7mI+aYAzVGnCeG6L5/sykRHWtXxKZucY83ptT+FDvq+3X9K8T5CtVZrjXjlaEr1lT
JxSL7lGqB1ab4VtAvBKX1X9OJp/MoV0DMzAmABv0nlj0s+ddOfbES6RxxUa7dOLvUhtZDDUF0Xdg
S3e6lobswgdAyRIp+R++jeGin/Wl8v9X9Gnq1P4sUVyrGBoHl55P/ElCwVGjeyjwXYfmk45hD/VH
ACnrrIZCMBFoAazVfbGgwAE7y7GDi8M4YOwX6ownCkmF4VWx4Lzr2j0yAJY3UWfmhHw2SU/wMKF2
c45/eo+MsOWAZPP3cNkewTqkkrQh0cYHfSxsYxwAaB/w/PVvbHr9r4n5LTgwHaLvZ/N6JfVPIG53
aHqPd+2ahG43WEo6sqprbg1GrN1lbok8Dj5SAcHq8f+SsB76QdkBdI+I0fkm6iINFiW8w76c1g0D
kIW17NrsuxRsCBRP1QisvQYf+10ACs4VGJf7XZaWiLPfwgu/5qh1HMiPgWpN/+REr2fUhSWC7l+9
YoYNV+0zmbPnn1YB+wPpSBN75Dk1bOkfQYpi2Y+CbKuiKcQHfcTtHMnujTiaSJ9owBbYlwfBQUjY
0OW1KCQSVLSjS+G5np4FFNZc14lR5R9vrJh/5aVtLkzsmyWF5dzZ1GkEc5zx6WxtxgjQYmAjvOm0
sSiqjLg6gVjU6mnYwSXc9EL1WNdwaZfayeB7Xp5PN93OC97W40hr1SejnrD9tzJSzJW+FLehXjou
omQ+YiC2YCzhssqsWh+uDVam5cHjsoC2c1mIkbYogwrHCVVmgK3q7+L35+4n1eoZ1pfYyzhuRn63
j/m3oyFDT9OV8ZUAQlzOa+7uorjgstTGNpZkWI3IqjIcubnz2FAdgkGQ/ZoMR5wykG7kiB41JpXz
8OulRSYRHwjvvG7G/n25JzWIG4Pj+p7ywObdhjzjt5VQsgfYnyZFl7BsfPCWELZ/4BbNxrLvP6Jz
aPXMBCa73v2+KfwHjeW2setM5f1wPbFyLOCPFYzIlWVX4GMP1CvseyL4QK0EY8cIXvmEIaqH+RID
uKu9QHku1F5VbhF1l37rPB7wrRjoVaYcuGnD4Hb7sfnQ0a6pNkhOgs3XPPnmMAlzFOkvIvTBAR0h
qE8RLoRnPuin/WQqzeBsulCelxmea7D268osDwGWKmjRLvOAYR6ej7hobEpWsZUzAAaduR//+tOP
9pkEryesD/GBiIdS6+dt/Wo6rL6HjoMiFC5SGlOtFUJoDhiB9uU6ANDmXIIAs9z12VDNYBxcCLX7
maLa6KPZPFn9YHZ/oRKRF5xFCtB4Ko1NQhxVpvoi+IlTamuunCPcJM2wWE6y5kKXUpJxbdPc/+Gh
Wi1nNPaGUM3SCBk4ijqXncxmE575XyIsBQ6430y4Tl56eHZpVdkuhJ3A1d43A3HBK9DiwWvThjBL
PKpHmWww6B/fcqdkWqZIFUP/RsOsbXevuXZPvdx5RxrZznUWEneG6upFG0ckUNT17ICglhl7MB/r
tmVAIXuuh7llQIQAR8nIBGcdg2eLWbk3Q9APUXbTx8OvAS4Wl87gel6Z1jrTSxcrjlNQecVmTlSZ
1hKhmvnw1VKp/H7DC5jw/13+0+fSRZ/Oy/erQ4+U4yBmF4vbeNzi3lnceNV1pBmHadWJ0iojVWfC
6VULrifxXG2yIWciOTTM4pQsC9DULad7PbF7oPuVMUj3nrxUgltw4lLTaHaMOkC2kcFowAjCFoTj
jdf9FPK3wpQreZLdxo0AFbqGhhlEVs2ZkZtnqalFarQRAWiv/X4RnNEYGhI8FBP1+jSsJuzdtdbl
eM53MCncvu5UZBKNjKspuamcMDi0PTgAibEkQ3uGdlvBp91eG9PjIqjBgaUOORrnmtqOZuLLglRc
JJEBhKE3Kz0n39Q9QFkOiqo7vU/NA+0BNfNB3x5JDj+UzQv+xKbne2zGutjvPR2xH0YuIhIm2PGL
/3GSYZuNLxxV2wrcUmOIpn18/77KyPP8Z0FoBBrudN1Xm2NsqW/bGfct5aYBPK1Qoyl6dEztT5b4
bePQLb83zhUGdxq+KBlEWeuqR9xw8EHkawPSpIMAgUsXtxok50uCao3zBNETjC8WyHKcXFznBLhO
gADyjw2S8SjUrMPxO/FhxNZqvGsGVcdHSpqdgGEUV8Qc88W45nBKEGZk6Hxx7PtvBwJGTiPg1I2F
G4L+uT83f8lBv6eFmAdi5UZFAMELpbiEpxme8HFxQ3SFnHV5Fs5XDFvkMPDKvXfxA337RpOMzVX4
dtbeqjOwkCpzxxbAssatrS8g1xNVYaxYKDq4IrajjApbOd9RgTknVGjM+dDyLTo+9YFglu2R+3Te
hwZPXaf3oBsgwILba++6XiCwwKhRqyTYRI9o+gRK9jE1rJugRCaiYHmHH577lTDGxo56YLlodbMF
ixt+SHXi60xgpFnmNRWS+muPP/LUyDICYYqKi+Ct0qmJrISo5jduQyAb8ckQIwaWdayT+YBeSsmT
wy4fVZWvSxW/ZgiWglOOeDWdAAt/n99Y8yjY8tYtaXAZ362J6u+ffW9SBLncCrS2YDHn5lSrF3Ih
MkYx8VdGXUx/8Qc9aOXMQS9jWZPylUA+Mznxp60WmB6ZWMlt4Zr2T2zdW0rjdHVfiDUTnRVkV9nQ
qDlPBGOkRzVN8k4OoEY2CEUk/pMKGfzC4lX+zVN0ZqdMQN+WD8ewXKaC1x7+P7N7nxnrYBtipFLh
S7e2gX7eAs57eUlWSSe7Er1wKMoaOHEVmtxSIal5guEY6V+sux5hetgLl7VwMWxxj51WpSVQhy1j
yFRpsNfm7ivABafhs+0QT/x8ZbBplVY2zygobbXShSiTrKw4LK/l3SzCfPYL5H7heebK1L6FIafN
xJjC2cIKT8QP0YzA+FS9+Nxu5tlBEqsb6m6yX4xz4OHKGB+80nzafA3FgXYNxPyeh+6F5I+ZiKDs
sGSdZZAhQKETulUTm+ItTuhyZCth9SVS/A3Qu5ss9f9grD2VZzdXBVyHvaBSiFcJKq8meJOSJJdy
PjU2+iM7tU3A1mmutQnksABeea8dlKU4lIt9+cr1gRjgdqCQrC6sQBPNqtEDHFxOWQuY44+0nc60
YRdX0ZnNk0/DJvDDTzAca3yEKaGAFJqb1rYqlNCLTgt1gv26zfA3SQyHDy2YsbytK/ibTlXnjhVi
gAfCg8aHB3df52UPrMQy7uv45RRYCFTPISGca+CoyRuYaNJS9y5863isct9Sm3Y3xkYM2gmpBNkN
PP8iBrSBCMlOGT6ZuIRjDmxhZwsHgs8tCFZZqii+Xsfs4FiXbVfX9TZEkLJNIwEAkCQ3tU/GvFfS
ZYmtPBh7qAUorFItDIqs2YY860SfIeernTYggd/OWmaaDiUJxwjoiiiAxFChZVinwTT2lhk9uxX9
oMYjf9l6UsGOUwT3CkDylxEHqt+luMlyni9D35fO2KBXgBl4RM3ntqg4FM5gktNzSeQHEhaUJGum
eFzkzG/IRWEUKA6Zw4OjbNjNW/eFa3ZPKlPy5cLOXLziZezxLPHlLTVRJD//7DHrVSh2n6QvMAa3
1VLAlLvDBKctpEKyrgdWSSFxB4V9Od9Kfs6jLLnOQFYW2VgbCgI+145vnzCsnDNeVExDU7DmEBo7
C5d2jM2I08NFbO5LnEV1DoiPeToHEVxvz0bb4KA30goDNxzJJtTdzYRntycWVSoKBuSpt5Laht9+
xSglJ6QMhdCVNKQ0RwFTZJMdqHWiJGoKfYElXERUQSfqwz+Pama4O7mOxwlneIlyt54aSR9mA/dL
2AgSpGypC+YFpHVtlyT8/jkMT6qUfqLDj021b3N1+B42Mp41/4N2a4c6Hk4cfc8e0hr407Ib0gOT
N3Gj0HZAqqnkgyJ7mr4k4t8Zy/YzbKM1TCfd6BHvtpF7jZNa86zJZjdmXYc9/IjsdykOZIDN2hjY
TO0LMxVb3FieQ1pK/N+egVhMyLBZaZEa3UTD8Qn7dvPNR0aZjg/Zyk+8/pSq4pH0qyEqriphT1J+
+I4WxF7VVdAPmPX5XSqSqAGAvdWQD2MfoJKENDei6x30cErPqE9ZDEtpFI+QMLXfvuKIECNbk6mP
aOs1vtLJQLQKn8dnDEx4Rj62nOkpMWWXjwkbR8claOWikrVO8BEqH0SE1eJy2T5/IZrW8xKZnwlC
cxh/OtWufgR2GTLv1r6+KyC6E/topbXNGzxGRql0WD4xVM0R+thZ0qKlSFCPnWmf7xGoeayKIZUf
lHptF/qMveDsO08wHllvq7gPIy2pD4f1d/Jrv0DQgQYCH02Q+xHIoa0WXiX4O4tpOzLeCeCemvQ0
Aud5GPQPG47ohkKTP9HwHkIL9p0Gcl6/xyQu/6GtGtpcSjqeVDrnDzWZFlGtyuSnLsbL04+7j7xx
5/RAZKS9ZAuKKCUZRsk8AGamUzTlDipWBsDVzU3vEJ+KP3EHySqFa+G1PjIjL0ZEJz98qsUqJTbr
4+M5S5q3AKpLeuk6MiXK+oSUYrNsrBSIoTCQXHD446kIvjY/mJRVxW+6CmjSUjlKbs94FTFdzsSP
p1Jto3W0Wt3YMOI9wOu0ZKHwgad+RZMExgrD3qu/pCK2ioObmxuxMX7vntNf44tyIo3iym/a4OLg
wlUG1maZWUpHxOPvEVFSgHFzRxDJygYL7JCec0Xwj4DTkeCcaH86+ABt84BRJ/VW2AGky/xuql7u
fuD/Q/ic2iqLtuPDaEENntX2ocwv3zrcdyNVlp87py25KUsRF8YV6ajiaCRmJaeXdu1YhwByfiCt
frp/InBJUWQhYkSzsqoW3yPNu6gp8SeUVz9/um1sEfgdkXmv3Yf1lJuUJfRupN11JRQpu7ggk8vZ
mzDf2X8TOwn/Jy+AaiPS9we0bIrzCqS64X3bA/0FH84ymXnNW3JFxb25j62KHF+PJtwOtF4C5jwZ
DGFt5+PKOSekkEiRmgtJdpoGzqDxBd1EezMmbESl6koDwfae1nP6WazrViOaGP3B4D3P/JnWk7PK
SOhsFZHa/xhXcqEWpUWedpo6CQTegtBO5HsTW+OJuoaCpTUvFU13ZkARBqW6c1Exxja30XcCSGzh
0Xln/nnU94W3sz7u4QqVkigUZyJxuchGJGdq/x+oBPsWZZ3VFgQSKZtN1HM0K5iKkRmGLiqo2AYR
nulqAKSfuf0/lYpLZdC1vpD4tvNCOz7K4FTld+ScBH8ZGqdBJ/+PstKPOL1npELLxZCG8UhdCJFD
SivO/nYoxhWTA4aBoRQbJ5qYNSDQAVPBYkTMLYXApL/0OA7jif82EtkWnu//tOMdxGYJ2bZsR1/Z
nRUR1f05n6+B0vgdgPnhGCIj+wVi85yRfaxP6vjlsY9exeZwYe3g4qOjxp6R5LOGdcUAReZoB17T
revgHWDF3pULCRuteWw8ZzzHbGep76SLO5kKHrJCRog/VjymjfqXkXc2++vh+MhvEtiabG2zIozC
Ew0vJDOukSMu51rcg5dbTm7Y1Sji5M4bN1RdVdA6aMD6LHYjqQTvnmjf2xpjMuQF6CcWHVvskQwq
4+k0JWxL2AyRBJ/kPCjG0TaZ7fsz4el2dto3ThsMlV7z6GRboZWlhy0tS7dcwNdp1MhLvKJ1r1gm
yZZe1ImJjZdWX7CjCRbwK4D0fFBIoZfLQg4oBNR6v8B8DI7wAiU+9v6F4YWTGYvOYmhkA94fROFZ
kS/A6s9foPlbkHXCQ9MmsOHHgoaGvWHntkZpE3aOVIPrqmFzgfnHeiYlj7OFyO23/VmCSpC8isq/
vL4DucwY8CwRlR64Yf5oC0+XNu+xKK943be4oi/zXC+J7+UB64rMUhu9kGEe90gLJNOafjp8fsmm
JKXLLqJHwYZ6xrxqTwLTDGRM2v0Rh8p5bO9GcynXNKp5kmf5Bapx1qhbKZSU3iGsb+jqpDyzyv3A
m9/LP4z0a+oHqCJJ53oCLLOw6JSBUGpNDvh7C8IfYFNbtXsUEDJDVEyl625oSF86M3WxgCPdQ+9i
5jy8IYhcNnC28BuaYSdG+DerNLILWF7G7Usak1EJEALYcv/jDyahV3iVsi1Gc1xvRz2fdAbcxs56
djJ8Rwd2WlmsZ2U6UhPbb1EoM4kTrOXM05xlSG9/b4EL1EfUbo2g4dlyg6A8gs552+0i5i7ZvARS
o/YFf6/upxS2i6TnySKFErfuxCL6TT39Jq2TYo00q3b5m9MoB0h2C9Bg0Rxbz0gS1eMrB0SqN9D7
CMQU85kUV2e2BZtI8ptMT5wLe0+6HATxTCOiH5AWH7lR0ruEZKnAWcVhiCalseGlux+o7JcxGexZ
gU1exQwS2MNh1Oh2lnWgm65UZpuYXIB5xcJ2V1pfwr+2fMI8O0P+C+CStRJx6K23O0rsb4RFFI6d
VFNHuvr+OKsXxK/daS+PCH3mceCJ2x+isN7RSnjXqBZqUDb7bX+GtpkedL+3YnHOtyeDEol2c39d
lIKyLsjXx5k4EHnABkEopFLlAWhZFPo65cUh7UUKbvnVkeQf1CuCedIlr3soBojZYaXBJEiKr8AB
VjMlnklTT+ULRpJwlFQHMRl0aCJ8v5c3Z0Yii9gCUEfAxjxpQC0szHF/x5lzWbRSwtQx69WIwwWA
26Q4jWHXxfQDDOpohll73EUZiAInxV7odr8+nSh0SnhLXaCshYjcktOLXiCLVLEyjs2uwzX2py90
kV3eWqeiiTqWDCWV8qN749wU8PcJIjN+vg6sz6XDPb7GaRaqb+tlp6ye7TOjnxmRZLtzwjbKGftD
riaxrm0GRPFgZ5DRoKC5IotZ7XBd1LLi7XlQPBG3Mi8hFs9DN2x7hH1q1/xMSlQDFyzBp2ERzlX0
tVme3iiAYpIuu6YtQHMs7vWvrBFzLcpVXxyKBmK4Hy/5+zcIdzROZSA0QebabE+Yrkn0nhtanJ6W
u0XGhKT38Rl2Gg+PNSsFB3WgZA5hcpEUQhxMMmPF/rTm8cUJrrBXKF1Zo33YQgANUTFk9uSzqTRG
RyuTscVySfcsWeDvCLeODay/z8fABLSqMC5wH5Y3Tn/L6gPDekFG/ukPXLG2uQyb3LLHh42YnhTo
QLwb5h8OnafhqO2HktlyU9mvUpYSoQ1sNkT89Lcph7IRf8hQITiRafyL+JkikcmogI5gywuygn5n
seytuaK5jUWoMUB5bEzBbc3qRWGbHq+OfDQwtaQIIX/84ASUXmUIMMYChhnLnydhTuZYkJaovtOG
xa7gpfH1dSTrLTj826lkGdJ5NlQeJix2O+vWw4PvI4I+DWShSOA1BAbTBepdi6q0ElfI06Smssvt
JgLzkzsJ1L9isD5Id29HAUHTK1q/HdNmdG0ZDWJ9KlHFjgx7vh9d1RE91ShcWf9KSrXUJbTYpZHn
bUU8+YZEPFYQO/GLXPKKSJ1Hh/HCj38mTmPRMLDE0yvMxf2MdBBWVt7kX4Gtp4Pz9/HeEPmKP6oA
2kJRZtcJ2uh01KC/ck8L5NEeYh7n8s83s09SeUwbSOVL5RKgVzyPQ2GEJx6/RR+Zv9lw7e+AvssE
wOwv2R7X1dJ60JPTR2a5nJcRrGDMRDEktDI5OyBEEj2W5mr0lERmnDsCPQqclOzIOFJdUbHObdS3
fQbc70aEEIM2ErOqeKRO/1gqES0671jrBUsHuUPmaUXl7kIn49aKFlDdxtgzDH1bvFoU+Iu6Z8jE
ey2vnLTBGIzkj36th/Heg+VSroJFbXG/PRRJcyPjlIK8BP3ea1oxDnPA2uBaBeaO+ojEQ3Kja0ki
DseZArfjoL13AUzNFtxp2if8en2+aXO9ZOrUZoxbUnHEP2H5jS/7aF9pb4Bgxdf1IfYIzpPJ+04V
LtfYJXJwBPcMxP0dxNPaNDqaGZn+aVg1JC6zaGbHy8vLphYJtJNvAlYh+xUrEjmK6gYBJH4fZDkj
s2It9MzPaH5NLoLd+YR2yop4wSvMbdz/kZD0BHGnzro3FaeMIelnJLeXM/JcWMNPa/TPcbAfrPte
gTjVgmbCvHB6mPLADSpKMtCajznIblpdnMYQ7fJXFh0XDetyzofo3QEf+WVuVpi84tqMaEIU5zCG
VRX5Objh9UVkgrdwyjwxNv8bRORI2eS2LaPgf0JtYvqptggFMi+DmZVG1xTiqjbRIB0mW52JFnm5
MJNnArNoddEOcMvbhKa/no7IV1XIpzfBB14KN+O55kdOycokv33EoWQMJz96rraF02VM4Q5fJz8u
olaZH7Zr5sv3IyI1IooCp2+BaK8baVqQXeXjnPHK/Y3EWupjavY/wlhSU3dws23f+acqxa7LpQFX
5CpPJycCRHVUe9eEnxSEBtworl4TuEpLVoJCUOW1f50bGbXOLEqIDMWdBlCwajY41kNyaLn+YLVH
Xp4naCzAoSlpQAiPMdpyvHWyNpCmEwesG5adrxPBOuLsihU0YqZEIVqUR2zEmEr8MFRgfSmBPAjj
VfmZL/gRdL0w0cn/2VOFUGehYPTRJr3KxBfFtoOhovA5r6QjNLVufcN1BflTWqBWIGDXAXCDliI+
NeMPeRRxYYUoTDmYIQSPrIV61WjhIiWl34DTpK1tf8GudyYZDXCmbmsGAsAspNW9M9Bc+mT++G1p
cWMau4lqnDkwrhuDLfOW5x++7XQjBN07Du0ZdU79qneuxp0NuchwyGohsnMBv2VFW/OlAP4DcOIm
gootYDp7MORzgFQdNLD7FtUrfrBBFdXngibDjlpnLV4EvR/Gh7JsBmuwF2z9fz3j28P5c39o5OWP
jHlktV06Wq76hJxl3dlPL7BIoCDedMQcE3QEfVnuwOImsyDMwimPkz1wVJIwfW1jyxR/ZSxsFI/X
6YlXcgdmaUHs/5oZdKsXEbwFVZC83rYOfezsBXbu6bbW+Pcm45+BmHyHvrn6uIkpEm/35gf4NSii
gKGXS+taJZFdJacQzsfzx12RFDZgnJuF/R7SgF0YNHHskcMXVM9hpTQ2aaUBS7rGImuzXLkBEnwU
7e0w/Wu5Ix23DTRbMCCY2dHpYvyNrhv1xJwMN4VAc8soV1U06zBrmr4w5sJ148wg96HDgnOOrfWf
+215hVBCnbUbuuJiy3sPoqzTqk7ryVJ2j3qHF7xByzRsp9pyuqEx8aD1/fb57jdjICsWDDsl9hOl
8E5biuefcb0odKDq0oEFuVAmCxS50eB+yXNDktXnl5O8Fpvi4led4V0SmxH3q2E1W2dVNaE9HMKU
NRNqXHAY0MCijo8IT2/35krukEKu+p0I4dvMOyDuRWCvk1Egii7L/+8aFZwO8tX6qpB8cKr++swr
MQgE+PX4EmLfko/DST6oCN2LAgz7cU0Ikd57MCD9Q4MEcnecJHxovElkTPZMtvyCwkg6vo/TwQBe
+cPXmii2CbxspdmbEQ6ILYuJRU8se6Qve3MuDUSCrpr6QAH+QgFQD6PVww35SpvKUrPdu0yUxN/F
x1DZ/CqSABGK1XBttJxuwO00Y96k9Tin1gU0mj7HMEnGg//Ph4d2lF4jfS1mW7meajguBc5Y9Slg
GqVWr18bordfYWSBjEF8KWZvle4Y4MGPY/LO3Hnuv1PSQBkLvXoY851Av8rAOk2HxK/Wzeu6XDEJ
EOL+JXJ3bhk8dXwI0liYaw8iaFfUqHJd+f7BiGMgkkeprPA+Mi9ANbKi0BMaTUmYnPSCoH9/ALKg
uuAwxhEjaAQ+tBceVKamcCfkJgMdw3RJ5TODW4OUC5zpdIkrNjDQ8GDjUvSj3PxhT1jd7mRlJ67z
YGJNEFwZv5hzkmiNiBVzvTTD7o42F9BV43lbE+ocQigEdaddLWeLcVevrLNHd7J1ecKVX/tXnR8i
Ew1RAVDxLQ4hdqA+Ke8z/4CsUjqLesU1wKnWgN28Fwt8GH7agRut/LR04raYuEzs0sF9d45GFsy/
Dqxf/Hy4l3tFuWWM7quFFFyc64/OM2NT5bHmAW/uA3phejYCQnpYkdGP2CCWFlFRiETW2xk4WKWl
zsKYl5MS6HTjB456zVQutNWMrKS0VmE+HKwa0exyZQoylH5Y7PkS1xCq7WfbFoPEuSqzNBNRe7/h
8MeCwADE3EGN0pLLUhb+yic+vEQKEzioy3d93vHWrYHbosxv6tPnsVJtyrdXSR17A8mavlr6F9vi
w/CGTRKd9iltabf08ZtpwCgpRGCRvUV5jG7kYL6uTBAZaO4b15o3zHcmrxaFNzUPQUqdXCGPHftz
JrumrMNDz+zn8KNNK7Va+u/RDKLfD2PQPn0ccUVnzDs2gTTw5herPo+tfxb7fHst4vwE4CY3FNj/
hJ9UOf9sOeR53jTuVUcaeUczOtBDEferVbxjubH8qBwM3/t8i41PSjvj8wBUlRxJiMqiSm7rSAiC
aCeC7iha4Nmm4o6IWmf9Jb0e6t+HsVcQiGnJeyA4pLZww25QO8zS1hSbHoy8AQSQFsZrmoehBWbG
UheKk6ptA8F8I6rb7fCOlgYnrSlqvjcllcoTsFgsXLeopssBODpAmFWoVPdsNaeX4rtdDOTM6R/r
YswbRWkJLVMcQhgzKh643BDo8LxG1+NDi2nXUsfC6r/F2U/uAA+T94/UH+jvryQdM8uf15popiy0
JGnRdsmojybvsqaAfw6aeRM7ctCzCnOzHEX/fodzIVE+KR7y+6WpFvShZ7GzEG0Xk0NhCANm0bCq
qr+qNCcTYxU1UfEStKoLPhAELLuQdF+eFMNp56ol7J+Gj9nKniUDCwTiQIFaFLTTgbkboM3iYl5U
6U8FJ4A3XyesuLSxKG/ZlWM2Zwsoc2dUC3L+auC0tZIeJtpjiyket2o9ufzrwV85+CoG5Z0bTPv3
m5h8SzA2NQv5kIb8vFXKLJarh2rdGt3JaamnWFZE11x1H/PGzqDe12ezsfamQjlUrAW1uVdQYXu2
NAUQLS4MZ3sejaRLfZypq0mRxCmfXAawKklpjp3tb2zBazTBV6pt6+u0NKMSfSuW68ID+ITUzRDw
OY59Skh2LMU3RzjvI7Oh4VhjR2zS+v+5AWQzG4zKiRzoFHaKIQhQsy9D6Ccb9uLFQYnby/6+dizn
7bnI9Qom3ebDMN4CYgLP2U+qitlyVr3MXel8oSk+er0D761unSClVHnoOLGKIyFFpDgoEsEqmAhy
drHVhipp7it3T+7ERaF82nvrOmWpnOZ8k31znsAkzrP425w8RmWYKEqn4AGNb8gS4MQA4vFucCdG
cgnkfTO4+CVsaFPNubWv54jA0GNepELXjTCEKvU+8DBttZlJtCTPW+aOTdrOazRoL6ZAPEF7IweU
EH3kON2UySG2O2OHXRUAJbxeTjf8052CTfz73P9asezdY6waKPxBsK/oQdN75t0MeVJ7Yq3IWH6M
ZCfzeT7hNY9I0ebg971VOWoxdycWrDGyv161cvMHUKA/eqQ/HxmsdwqhukWDQ8joZt+gm+QaigU5
a4a2X+Tv1/R9BiVS9Y6m17l5drbem7HubZUepYF3YOqfaQsNyYiOcvlCdvtPjjhf2cNaKupTFAsq
+lDUt5KqAQ5yETOmgJzqo6jTPJNqXXtcZxCd9DEgcOy4kmntTt0D4HW8IYX0lOdN5Iccq4dxip/a
7Fho+hjTm9Jh9LsYwXPq1x4SnSjSsXChTwoGPdzwwd1A9ZetKF/ofUXprnQfL+hJafbUjcWjK4Ef
rgH4O46nVRYeknZo1Qrlvhwf5M6VQHoTdzrT8zxIi+Joo5vS3JkZwBNpYquL9TzYnuNf9n+N210j
mWQ0Bd4MbYJtrn3RW10rlQQJ+s7Yyd10+XRCOj2mxBvNn7/lO541ysmXrhlwGx1IOXpE8Q+nsYg/
0y307iht8Mm2XkvAWYoIYCao8glisBo8gqWm6w4IFxTQ1Br7yK7UJdI50AEYhL0YyWihUX+PTNk4
nyjSNuAOYTuokgGl5Wtvzc+GJGhXGbRFfo1FIge8bOUwMV9ypfBDj0Hl6Ok9/v/FPmZUGdvNTaPz
Zc+9iJ3a7YEGeXA9z4ptLvHTRf53y4oKUkr8EoQJQMgglFF33FQwWyhbPcDrvF0t/E/aFGJfSlsV
wh4AOlxNcFx6gOnzaII/e7ktHl8Y6hnMETwNYQoBagwHxzP0cyr2AFhtxG5xwVh91Z7TEaxb1A1+
9woSDJJFnDIQ/MzF/iOuFC3+8il9mW8SfGcDNW7sGNOzdNSRd14NptWk0mPHbyf1nybIclPWkuaQ
Isk/6ZvTYHEgyTiLmzIbM/bN7n8pQGZN0zOhOco9FrReegj+oPkGcaRfpGA4DuLu+RmduMQ65cgb
wgKhDpks5451ox5hCPFfXaQPs6brH8C8bHYk4fPgEjDWRV0geqkOlFN3G5zORw6EmRc0Xg4bG2qR
A09D9HloamvWdwWflRnyAFn8727dFu3QvIIvsAzDPlwWRd9wtT+UiepKTI9qd/4RIC9WRn8mzvGA
D+9xZXOhHgVa+CSn/tSvaAnasYm4McEdgK6yiX3M3pTsKMWosIFOrqyAdkir2s+o1HG+lK2QpOvD
LOg1bhduF3RDJRB0nO0mipvlo+zzBjS/hhVwkVMwqWjV4oBEaJuEUY1zf2yDiRUX7JX+PF4XDVtr
Hy0MapiWuLLfBVenpybSBIpWswhZ4qIrUFQeIYYsBuue76eQOqucFMw/ZQc374ensabjePGZFOab
iOPQ0yyBlKEwETklzbjtvXfru6qycJsA41WAx+MmpAD+muZxNpMJ/KNWFReq6klME1X9pZ3Ox3q4
rjeDi5v863cl7vVdEov0YJeJFUplS7pt5iSJ41/eTMhV6cbipSxMo4XfCKF0wEzV3JRTlqQXQLRs
0cHleIywIxyOfg5B1ZLD5I2GawHh++n6fC0BkuQfXV6diyg020ry90a8CANmlDrr1XJ62TDuiZph
BED1aRbCa5xE973qFMYj2nvOMkCH0zgNy5g0Wwg4jZH8FgtjQaOaCOMbwRgsLQ1JwOe4DPF0mBIT
q48VgrI5J/mT3I2tQtY0mbpmd5iAfEiKIu7yEY2qOUN1Kj4pmehagr+4wQevqMWsOfXExHRHjO+p
psibqx+r8qFlUYYvkgZQJwTAvvytLGD/5lwP5KuqUfylrXdcVmu5HqXyRjbdhXM10Gp6zz9S6P3T
64V0rGE3iBbFUumG5hiklZH915He08oJRUXUjIUzslUMWwyhtzKD6Op+6rx0jZK7Uqd30lBTII5d
w30MovBRBbisP1CtUHIQAVfOnEKV6tiysaEgm6Y5RYAk3NfVDrAOhJfbl5F+vXIFcsFr0iDMv5gW
gzt9dG2SK8EV86h17d6ts9H/+hnIQFV1cR1JnaZi9DIJAPplxClkG/yEXeUZmj/Ih2rxMqn0stnL
V+RhGsFwPRT02xL6jqX1Jaowc+BEDROlkc+S4iNGdcinrXNkoao03oPzG7Cc8TBCFzygKwFtPoPp
00Cpqn2C5KtF+EWOePeFlkGMb/jPKLzpmxk6efWj4DA5E+/b66UkODNvdDwgRh8r6Y8mx5j58k9Y
m24BjLFHkR5ZMyWMxv2wSybDIKZLSHzKjQNNGbiIPCuOE+yHHFXCu79YplPb0KSiGDoB3PtdPCVi
68z9HpFLZ7PU34TKkbxWY+upkWaPc5d6VPbHa1rYdeNZSGwZJ/6PBtAwwVoph8xF1LUSNB484wz8
/qZskvBzNVAIpizvN6Z6Tj+x38vOMSGpPvXog1jaUn2bY24aTOQf27aAwO6fnvML7bO5BcbitVAA
tlVQ5nek23kyyrI95a5G297gYIfP4iJhWQGHSCQQ8eTMGc+GSfyQj2MMfKcD+GAvueME17kAHkxO
ebzt6V94USUq2ZHwMUZCyeoc2lcFWJxOibPsl7BsK4zlYFiJmrNV3ZfUMPwXWaH9xGVwKloMeGkv
lVU+AGl1HCd9AJx11RuVEU6Ks/J1tkeelNRvcByLANJVOvaktIUVGswIpYMeN96cC/2pswsODUdw
JTBH4zwe2Tft+oFna0RjeEAR7g9dwMYu2VY/yiv5jVQ36i/9eSsmWDV7Rscxy5ArYuS1RBolXLjJ
NWJN9pVAMk6ptTglGr08yHPNKgqGAzeyeJlXT9KdG8jd8Vh656hyky39DO2MEMXTu/C40mMAwf3i
ejn3If599vT1V0J57rHpz1n6BDrKMj1qeQGdvLQbP8Tk23AWJUG77CO4rF8rGiGTd7b7/3X5TwnH
REjBzwtleo54eJwaZEhHRaXVtQTG6LWngob/5xDcjZe3AJXH36xb7PB0p213L7wLh9gb5mZg4Xx4
HB4g5z0pvcj37y4BjXh/KGzBMmv8jDkHtQgrPQIXaiHFYaPNiv+ZQ/h0Xx1JiweP+NObM1XUpNP2
+dQuqq4G0q2vxelE5CuOONOog+8pM1k4VpmEAO7s2acUMu1Xe3zuMRHz8aLyyKlRGodys9O8KVL+
PG0oJNXJOOCgxIoPRCcKFrCvzXtbswGjuxGjD+qWxoTamikbeGc3YjISt3Cl/Yh3xYrI/5JNt7nd
bTnhkE6OWeTNOs6yANHFb18nHN8EvGXnYipAKJA4xcRtO1rAb2RengjgPb07ctiOtUAtmQzG2jOu
hGTCIv7RA0VGSvg/U79S1E9XrJB43u+5ULwLjiQ2A418I3dZzEybq7rGhW87WrAU1ppdZehB8h2u
SrA6YRfPJlJb55Ud91Kjm1TkNx+7E9W3MkS9LuHAP/A6bYaPSjBgTfmAyjkztHtyU2vt2DVNv4pE
g9HDPZOThLJByY0xGAkwhq6hpAuo5obU98a6kRkz5zLXlPWQtQP4M1y5G0JXFoHyp0Pif5ApHdz+
oHjuOIg/WQmYcCbq6hODVyY1e1L1Hb5s4ggi5FIPBdlBWqHK+TN5EpOAvA7m3zj8a5GdbKID7ODr
nUOY7+meNHuXvQRYh4MbQrSyRDfS9R7fvFiDBdvBwTIy68ZhAhQJxAQdbUSPADfJHcFaGPG5DSK9
hN51TSJXVXttN9Z08zWm5b76zCikoSTLJX1IQ3AB/Iuz3u6MchP55Yeu+dQoWrclAdJKUqDR/Kfu
Os0zDjl9E2Ubx9m3MtYdj9YLBA25921LnLod6W6CnXgBJWJffF2grYDyq6VjnyaoiJt3a8WbYM6O
Y19SGTZNzJCZMFSvsX2+eDEEsKUR+5M4/Ahm4IVo0Hr1d5xSMR/Yqs9SRBj8fNaFhL6ML6s/PwgI
XvVPGGbGUOfJBKsn1J8fUIQRPpsGrWSZxNeDYzQCynwytSu0KueP0C9i2QTDKmeRxny8ZpFvyyIn
+B4JU3hhz3gmSxHhlaSgEUvrLmmStFkqdhJAqJ00uq46b2O6fCjhMU7Rcz5rddQmSxRnU7eQfD2D
sG8Kyn10jnDoLtxsx3K7bAEmSskI74JgSEZs5ZH0xU/KQRwnDR9fEwfA83y7A4AtZ/GX2VjwfccQ
++eDxCy1a/mjBWYc/iJI5BGUee7tS4MX59ObliuQsnvNUYpQqwRD2m+nLABsZyVjfUzI5J5GiQoc
vz5G0Os1UsrzNU/J61GknDvKV4pup+wKonc3blbg82uV03uacnstqWiGsZha1w8fa1wpJ4THNYkk
h0EClxR3YZ9gqIR8JRemT9jyBLr5yvEK7nd6UlD0vi6kT0Fqzpu5mlTIRkUrEXXxpQxkA4ndFozo
VKLauDTxOidcIL6AbTZpnasxjVyeAn5W0kWN229oKQ9XNXJdKsL4ZRiMrMTpdUshMdoIaMB+jTDX
UpETbl9LxEYXKtTlZozNZ0p7t0Lvqd/g3z4o9e9bTWx6Vb0pNoB0uDuemD9HWoCGeVv5Ao4jyJeS
Jvidh++WarhSbML9Wh2VR3XrHynpXOO3qKowDtFy5/n3wFMNP4fAZ/d4qlRcgRYnJ/rVyAacL6On
8imSww7L//AWRmzJl+T2ShmAPWNn11fU+2g3wZHh6dbC2GQFzEWgtI+EaPONZN5Gjs4G/4WsXU5/
f0MTFF7HGuISkxKoRlP7DdJH8AKufJfcoRe5YoG64meUIVmc0VvyrqWkS2oht2prZiVhgOrvsHlQ
R9jh/5ZBH9827odTE1CtZ7TUqyhQFuwWGnPyUpwIpnR6gFnMpXdNI2HmqE44nvZHZ+vn30UqGfY5
WtLt82u+ulgqKSLi7fVVjSN1FAVsBvIcl/2XMRdk7kjnkl9hhRyTFXRCDmTZ68oZhmtNvKzb8Uoc
v9B0D9/uusgvGsOENxn0Ax0jlOtCEUqFqORqO/zHqJphA7tkBJFeDCbyDBGlp5EgmX/KOuSJuiD5
8ekmy/ldzC8KDCE/QYwL1rsp05CT8Ju9WI+xs0NuVaY8+mIUisaT8cd6gVpfktBS+Y0ql3CLY2OY
TpZ0hRNQSHLjCu0vHYhJ65+dgGbtCKF2YUCXC0cpX6srzo1/SN9lJ8WvAH5EQtgjnBwF0EueXoYz
B3xQxvqonxPobmeDK+ZiCgFhO3gw+4DQjzusQMlh7ax35kFIo2W/kjMQzRXQZn7EoUDo8QLyXjrK
7Jr3H67Gy1l/7wS9+vC1D73uomlbeZFk3oCkNHxhE4ad3is3Lth6KgCyX1wyOBn9j70bA50r79xX
JBpqav64yKR2qiVfyjF7FYUE8JCtPv/C9nWrZwTZTmqcbLMUzyyQPDgqBPJHMDkTjSIsBsE5jsw0
LfCW4+Y9c4FlUFX4VwPidm0Ja9ZuZqz/BuJg0MgCqWoCQK6/8/Gw5aB1O0tYXSL+bARGjur9t2WM
XlXXvQmJT0V4yBF32L0ryS7MrcF56tOy7cFilF4h0SJMqhjOI42Vy5pylFNK+Ffj0P1wdNjp644x
Gu9RQKXjqkhyslhkQCtm5Wn8AI7px5DWMbugr4UDaMmYCzLQQDr6vTLVs7rt/1ujb7hYlzgWj6q4
C7bpot1xVy6GLwvWofhnKlIHSMK8/cQ7kF4zVKRFL/3RM97Hlw2GwKd5i+/7zYdyPFlpi/TRPvqF
LWQtuSTa7YBF9ElAdjRcKAWVzI2/4/uKq3aYhLJuagWV40rjjYNlhUVq3b+SATLGbQteJG2tYeTZ
Ww2UhsdscbpEwKIzBm1QDs53XXwXSHLC4WkdvN9xTdjP9MILy72BmP1o/XKgyQLURbcYnDRMipI7
qZ88tm4h6v3B4CiwWNOcQl5czQsp+NcdazU+DGdXqdrVQ3N+r6wYseLdijLCT0af+omlrC5L3Smp
anITopJPW+SwJJiJHvnEbJdGf8vJJaonbAZkwB27ko/M34ztgueKFHaxzP6uMhB+VQdKtlGMZyQi
WW2R6M4XyMCpbDHGAvJjAyAUkcZuuZ+TZ3jpSX/kId5qtdgCDuH74JVslxb8Atlt/dPwBZ8s0MvB
+0R1v2lx7Tos9hFkrigpBvAdbK6vGbctMPV/eaONNqR1ybuB69dwUAn/f6LGsXlhodXlGDmZWW21
85UWDCdePTQlJR13WmhMPneb3/eW8C/DOoSel9oyeuLnruCCAZb+B8tndetlIQOAqhioTX9qNp2U
+QmDH6LXGhJj9btnmd2kwLPIuppXNhKxqfzRwDVD/NhDUKrFs/qumkFvrpbiR6CkkaXj5l5Nhifn
GD4yqF5Nz10Hlgf531bKu0DGHptvhhYS9bo0EYIe4qXjF/98V4rKNOB2wM7MmP0ZucoaUDSXvtz7
oi8WKJoLhnvDwZoW1cdoaIMnG3mhZZcYNjxmxU4Gm8llEcoPH94+MPscwiBoGXYwqY3gJDKIkf+9
QbF2uHTp1brTlXr34KYJfXpqoGEUJOb8pPjM0ugr+wg/M3g649S0gITs0F4Xbayzep99U2EmXCz2
2kBwBzpDQkm4wnfth17KxPJeAKy1pp1SOO9TfT00PCUMHjy6TVPRdJMbB5pKOhksLKnDGN7gzaVk
n4H2INBx6896v+UpiEjFSoBLDOavIxfl1QxJSkhm2JdPOBnZ5u5GH0m7Io95KATwFoXCLCCcv7Er
XOFavf95xEn08tSvXFdccBkCOy52SiF7OvkE6IFt6fAS8lM7pLvcnSLurYlzA4kLCK3/zjPyUCNv
3xZOhQJAr3v9aZol4sayiXz7gS/m9CX+KAkERY4aArsyyxDN/lmsj2vDRys3pDRXM137Jli+6M30
9KyqH/o+Tb2qxv2rNfvphP0TlSQ3etmoYn0qBJLAQrQ9vUmgNOEIyrHjdm8R+1wPdTNmw1q6zgyD
DeYFm0L/yot6yDRZ3pKvuvEsiUmjkkav87cuy4PJyA9qh+W16WiUYWF3usg7QwT7jJLx+SQPP3b6
apUaLxCriKhOEOGL8QN9patf8y56U49Dv7IkBcO7zV00xXc7nOvC6Ki891EKmrowofbMqnRuen1Q
lvIbvVrnQCTTIv0+u6FpXpuyUj3TMJSLNGeQVkmT6hE90bxtX4PNXrbB+D1Vkpj7HpFPZbBUTPpU
Sf7ZUIBhvOUbuVzSHPpIxtt5iDJoP5bFExO3P1NLrYBd+0KvhPBjd2XpBH2ADnP5YDdTyT1p568e
7vP4mxeKXO4jSNCpM9IraAXZIssRh6WjMlVBLi987ecLew7dFvGulD49nKncbM+rRiHv1RBdNnys
P7c9bIaiRaeKWt/DGwwiAJaBg7Uw+EmvNsS0bUqj5nvs+IV/fcLMOowQp8jIlTEv46IV+yTto+1N
+ars4mUnevBWH2DUPMqRgJlHLRIC9LpOXqEPlaktXFV0OJb65oOTP1ft6mZx/adPFZdu3TB5FDay
uhzAOLe3XcQyNHxM052zkvn7pGoc0Y4dhgJvo/IjHN2Ccw9VsXVxgGMBcMgD1iWk1F/NP96gdOi3
T5yYzlEx0p2Tj49UkNb80E1Cd9IOjnUs2mgsDJx1xvI7hvcTJSK29312ykCq7zpMj0wit2fTiswp
Ag1GTBuHe6GyS1eb7TIdIpen+sVKaaNi4Nj9HkEJZ1WJywSPsbyatvlWThv1X1NMzYtNsrRL2zf1
lCwJzeI7xBXIAGiDRx3vyLQ4QMUOsoLY4ZbCykgblbGnPClndx1LyrJ0UoIW635RCqtAxCyqVvSn
PRZgdcYXoFXrYWmiwxW9JJVChBp5rTuCNxN7uLQjqEX5VG6640uUbb/amF3RogJbJXtb6/ZuJmkE
GEaq2eoHewxZ2KkOUsAlhbZvOxdvXXhdb8nov8qJ+/i6pKGmGUAv3sa9cQunOKa9/6k6b6cRJNED
EIpMVTX7sjrLW6v0mLnw3xhP2kbjtpljTvWADKklZ5GQboMh9XtQ6xt3MQ7VPFDrNn0kP1cLwxJr
TcJivRhLASGVB2+7Ld4iu4uRSthVVw255nok0Ndld8q0n5bF3vn9WpGdjQxlmcM/avudiWU5BUA7
xhwHGmHoHG9BjVqIRg81HdzsgI2MNcN7LS2F03iAfFmdV/XipI9nATrm/0Krk2mCLuHWtj97TXDQ
HUD+0jvMq7kq5i6SqAuaNu4GOzEwTreOLSsaLcCUrMXxhjJYUftsqNFhqKvhFOpncfe8kyvfg2Pn
W6XsgBYux7vhBqKS7P+ZcRfWAfB+rO8R3q193+3S5gQfjpCeQlYS3VXC12ckRXVgShKeELsXAJHn
+yFwOi6Fp6AEGbDnnn8/atecX8qqy/d8v4/Z6qLEtq+X1d8cRUFYLPBadYjdkZYEi0yiLuhLrt59
jAv/EjpJyG2pd+GH6LgMDGtgDZ4Juj6IeWBK18IT2o6NzktZMCKipaxS4qZZu5tGeCVnxOOZ9sTC
RW3Xu6nuWZ7vAhqcy/VJuSlaBKV25F6nLoKKBNUj8+Ie6X3EhP0rsRN2jy09RK3QCUfjtC+KdfaX
D7lQR7oTg59bxzkYHmGdFxXwdSRHBxLAql8vZPZxdXSurx4Cvcnf7WlmQumwYEAVFEu43a+bPq2L
Oyg56+tD02GXJUKDJ16Uy4ZkarHw71BEJGD7GBD+0PbGt/eirzk/ycXz4RvcdzYi48Ca9jBTJ3Zp
Fjn5Jd392RNmnirzTQ4F8FXEwYL4wTVhqNMH3wiEFtEg0XIFr7ViSj/2v4jyM65vLLfK2WRLDM4P
p6lbLK0mouX/xAiGV4nvuN9Zqvkm1ISSVcM7TNgCCKjolDalaVZx1HdA2Bbnt4AOLX9aLny0s5PL
keKANsC9BwEEfQqJqQEHLCoDFWRn6Xde6zfbvIU7lNte6442wWXZjkKwk2BymYMf0FywrMfiCycA
82juocR1xzzP3cFSuMourS952qK8ZFKTzNuk5h07WPTVdbZiSzgjX67kob7Xt4G/vH35llEeF+yW
c79da3pNgAQo1OWY8dHAe1W6X7YlW48ima2IIEuprEl/4UKilvQhQpANrlX71n1sCUu9Ky9TtquL
pd5099Xql7lIRDKuNoKT3B48aIIzE5SeQMNyBNP5iPXyPyIBLvL8TGCsTxyNz/mpG7aeSHYOnoo2
LsMBMlsIgO3J4Gtm7z+Lcdl7eu74/T6NnXT5MOaYKtgzSy00Hdm24DVhI0UTY5lllzJiojsBxdLV
G7IkOClCmsMMBVGkV3+3Qm/IHfHGPhI2+Vdw5x/CCorWcdygCgu2B+GuFaNQHtRcezkxs1uNCMYY
g+MnSdQG8Ql9dlFgYkRJP5+iCa8hewJYE8l4DSpPvdgNgDLZpWyfAENDS7QFeJaYxAbLaBu/aPgO
EgWQPsor6I0ab8NIm84fZlK8gpzTze7rRNBhJatasdMQru+xH2VsgeMRY7KxkQmbmCiQnKeNJY0U
e4Lk1b9RZdBq7cNaBY86Uxq2HmtIRb2qrn3WBfdNMDO0R7ZoWlTTdyX7kasjJpdd3qbu07TY1nfy
2HgfWfowKMJe9ynyFQ2BQbJP6DbnYdn/W63qyi2JNxIkTHMBgSePKTA4TUjCYqtjgxeRBhK8cZlb
7ppq9CgeUlpes9/9Xnx6JBOiwJZKwy9tuPibemPR8AHcGCpK8r2mA8xlsle4djvcrcT7md9jQATP
lKJOjazWzebmDL54rhHtjf67uc2sdJgWGV+2mmkHcr8rtp/f7gIWshCcdmB557+kA40nwrrFciNL
AXuDDIc6/WFJ0PgnCjaInjSEcUcRoxxXPHfOvUndjMnbtkWQ714ch82f7EEEJr9sukAlGzkiJEpO
7aLkQ16fnR+8g3YNemIPZ+4MhCs4GQQwjPMc6TnOho48G4LZ28n8EBGTTPkrm6m4Wi3IioFIVxsL
e9+M1nkIsBmOajTxLqyfsaE1tDHBfpHJsnu6Hsc640OVeA7EY3CGEtW4zeIoBqwhbjJmvGHjhOBB
R49cgWdaBbcltJUYH7y34AWc/d9iZ/wZg4xJULFc0PK/ldc9/6iOtM5krtxTQEDFEnuEQCbNfrCZ
TkXdI0bxWi2rR/M0bRkNwaK9jwtWyUQOChxvb3kbbWTpBvJAKZKbw7tPwD3yyzdSYX9Q+D4DWc+o
tPEN9H+EgBCx5uq8YHnxfXNO7YulzCE3ZXVXt9rCpW5r1mf8X7gTyXFMCOiInZoT5qBVLf9y9kbb
Kjgh9W/lcKVubj3IOO+fMjnscuGtHI6oeieOj/goTcogNF2878uHYl8FGhVMSqUJPTvZd7D+EWLv
27RIOE0au+Qj133zvwD+POXpplbeXtAR0evJwqd3dzA/lA9E5HqQgshLUGtqcGIOUa0OlxiXOpY2
0r2Lf9vA/ArGQrG9YVpjOLsZsFV2oVkhpXvuc6fGFuU+5wwh1mUJKippsxaRitZ0Fwg24wwYY7n1
RwF73va0u32p6YM9zp0jIm9f4n1UKMSbkMn6f8XYdixbCHugR4zL+pF7IhtpJbLyz9bM+opF2AwA
mP21kYm6XbOJH2ifqvVIhJIJV3WisYwGgOQ+mgrpOqi6WfwTELBrjQq0FzHyPIba3jeKoa/uaHM6
u4qCsFOcVh0lchXn/ZrvBhM5Or1Bvgj1ir1JM8Vv+s2Pch0P+FhmwpVzVSBeBFspZmWw9cqs1rlR
WtruyMFuYq66dPHPls6hvS1sNN0B8RQbzkdqSP+I87pyjKJR+q5zXc50FwW/6QAEfWTT6vBtyw7m
jGlugoPX3vAu7JSuQAFc4w78EK2dvT+ROY5cIDXBbWhTaIz5WZ8ZZbUKMPXuoqCbcT4fYVHYr2Ta
lVnwMqJ5bRonQHW6jhYF+c2XNJOnY+bwTJ2VoYr8FUj5UkmYrGaZAP2ka4hJuQ4ExHxVciEwj2Pg
VssExyi50oAybESaN4ri4ec/mpi47szV2RuV8fQi8+aONR+ZNKLs2ZKh+MlzdAc4SqOKjH6198nG
zwrUphnj+lQioaoT4R+0jBEX/xB6Fi9xK60AR8YGKUdNcUtov2nVwbY8jyDdw6CyysHWnpbxoOJt
e8wN0eFvNPfkLGORWoVla9yniboWhWOWHwygCBZkWKDmGRqg/fa0vtEiNFX2GXvkQM8J3sir8pQ8
8Kl9Whmkvdt3kNidJ25vlgmqTfxPqvplnDu2mGUo5nmrZx1HIQFgpZvAl7y4IEWrrACXpa28Qi+w
PKEPP0TlFjcYRue/USnaV8qbPjLsqW72aL4xAosk+CXiWeZh5/hJa+P2gggsR9Der4BldvdYMTcK
5XiNvPTkHvTamtYrImdFVAUfKvnvit1tdaWtiEzqcHb8LXzZg9Ctts0RNLBMtsv8kumIBYi7u8ue
+DGhNKpG/NoHKUtcyfbX/7lryzhmmdAm9WmB8iL+GS1p1xXv1Lu6mbIMYe2fdxEqsgU0rcbFKY2i
Qufg6UGM5xYzTzyGk9zUYLJGUCsdoM3qDCK+pdisKUOYMIiQVONNoLY6FORTrZtqeEPnhK8BQNhT
Uo49o53/qzrBhPWinAp6BwBcyXeVQZYm8GwhZmQZ+dCj6qtXt2qqr/TXy5IaastoNoGHpEQkqzhE
FOifFf1fKMs7jGfZb1f3V4g8UNJwvfOhSHqzK74a/xWsps7zTQUq5mKUhC9uH3gFGc063hswAIyc
dynh/0iFnpDEkkHhcnV9fTq/WIacuG93x5EwVJ5Fd+6IOL3AbhZyQEctm4pmVKUP9m8t1ulgXA2m
E/OjUZBxlcdB8ojjkeX3GSO65Q57lZdXXJXCSoxEaBTOC48VUHkobB6k1DTExxG/JXyFpHSB6qSm
kcn2bIruYNhdMLVpUJbuoL+G1ZiPa1iY5fZbkiWn3NnvO0Tq7K0vJbhdNa38PP6h98T0Yv+L9y7k
RLSvJUxyI4onhOjcf/zPX57zNTFFZ/87X2+JohxdaByCP1cwQznUd8QVX9Jn2FAirfOSRe4rl7ca
S355LDk/rd+RZJLM/YyIhk4p4Y6j6Y5irI3z/MS1cnktmCGEBw8zLU2FxY/8be1PHFgKPigx4yHF
qEmm77H5SYTAS6P1SBS7RW5+uXVLgmj90bhGTCJ3ZQJvwcI/RIZ5wQLtsn2wpY9PEKObcbsIWN29
IMdfB38XEP2VKhGYKPX50YY8SrZhuFjBk0l+BT4lVk2LUP3H1R/ml3imA5Aykf51wXyinMmqeLtW
UxzvNakfqnpv+cp2ap6OZ6iMto+JLlF4lJb5cu/oGmwAoYxUFeWLBPH2Ish1WkR8GG+JjAVLcAyt
oxJTEO06UkwAP6J4CLeUJqP6wyDKhRFtfX06NHPaMJuC1DyLo3q1aI2LYsOiFRerj4veulR+aLM0
d9i087n6J+zV77xa2/MJR3P1ZGrErk0wCGkZSwHK1BpXvsgwjuwWEpZcCfXtxfycpgb2omj5ds+L
fAUd07vVd62PvmkbskxwUN54s+kF9bxPlN2WQ8xUGVRmaotTQgdnuzbTDyv6RD13JXr0FbYGeOuK
bGztcE7coXYVASUmI2T0TOsV79qHrQgZZpoAXxZrcJDGNGjw8gjCjw5WLUHum4uPOnA9Trai4es2
2wMd0VkOtsLBKuZ9fwV2e1GRgZ0wsBSZlLc+FeUUjybrVwbseuF2rmprb+JwqAxZwZU68QwYpp0x
tsmdQrWcOg+5WMnWCUm5PudzQcP8vk1wj7DSx8a55PHRtx/guHfS60OTwRhyLYjlUMrWhqVm8f7C
1Dabfz5KM7NrvBd0U3Sv8ieE6UTh0bZ4g4rwQ5aky8EqH3vybhMhC8a6w89w+Ghqnwo+RhTGsTAk
uaZ4GdGsY6FGXl0Iztrie5FGKYRF7xA5h8aXeNbMK+IBiafDhlTd3+x6qr5E2VU7IaZzOmiVIfwk
MWHZ5MlptMXVajFFtAZRN3HCcRP6XvpGSo2F8Smf2hdcV50ghYnOVrpc60ITiEGrwwSVgnSsDFtn
kl6yENJ4xLin2IS7MMsxUtKRqN7FK9tr6WBmWLuEmEzUOMOAoqd4R+6RwcqOnwsphtF1dxbBKCcA
t5HOUTBX4WrSWD66ziaGEqCgCvQH+OCy4jhnXnrv+08BZOG36nPosHzY5Xhaxf9piUd6AzIbJS9w
0Am8oX2Rg9xJF3vyrsIjh4SVJfAmn2mrA43eOF3O6XHBdD2H2oOnnzAJ3DQQLtwq7JKDt+wHw+oa
0ipgsf2/YhrXF3gO8Mkx63fJ1z6ro/fqK4DcMrv5cR30MWkhzTnqRl6uaRgazYVdqIgnEZkteb2b
RrFwpjkA62aaBwizHKH7TR3PibcqANQwbXkrCFxkWuGYk22Y3O+Zw3CwMzkRoSgaKqMJZmWxXL6C
1Y44JLAdLeJSndFUPGjFJjG/c/S3vzwVj9nPhl/DPfM5o5z00rirlE2VG/zL/Wx0Fu8i27TqBe0v
xpU98Ml8FuJk6BxhXaGAOZtEsvJ4BeOEWlE2LUk9ptA79dHAgV/W8btAA1tvQF8RsRe2anIomFzw
FZwlT94U5O1GgqZ1EtNmFXAYlLbNZTdzzqK4DXcJorJkpIe7eEqjubynBhLQwv5AQplZrDoA+OU0
P4co3l9eDZR1/cHOJ4tePc5UpOqMjlJhWpm8wezjRgpfoFP1Qd07VBEJeYOhbKOBet8okh3pEqLD
l/qLyDBiZF4jsQfCYxTChZF82bJhjDu6lfeNB+FxYpiXyqmBI48WQa0jBmmk1+IC1lbtFXk+y02f
CCADcEuU33p6p1W/EGmdZfaUDmryw1jKu9yf+C+dx52hRvsP1mY7up/zid6ZVtno9MOsTka9qLyt
Q2udXbVuaxTmT5P2bI9YC8u8wRuHyAsFfP0wbil5gAB7v6PdLv+l3SzUl7kc1tunNBq02vgqeKrZ
51smlyOtEU6BJo85LYlnqbGLiPs3DJM0S58S7eoqhz/LtW0t4L6c9pUNqFBdvtukfFJ6feSRKHsM
lCn1RSfqRgZtcH1uFVCeKYXoT6RqF0nLQnb/cssJVOiVLOPIdQtd4tDWxOnIdBkRmGAoPtYIGt7q
ARG7oZUynkeJI+Ai3OmSO4w3c9qON+M6z5xuD7E3Rb7O8vcNa+1lMneJYbOBZ4HLICtYMabafolt
TK/dsGCKkU419xi29BMluweHBlanR2d440aR9n/N8GuRkEknLyr9D7N6Se3YT8weUr6/dKbfkD1A
askQj+/W7xUrf7ocuH9EtTy5s7R5gz9CLUotOZ55DmJZFIC9p7s32niKhAmezicDkXrFMEA3jrHT
Mte16DvY0GQdJq8H/uQ39i9U0cUvldLy/eNNk2fgWyjihf8awjrwxJvPl3Xj8UrmnyrGiN0EXm1t
oXpIrRqq8RnVoFguHliyQdseleihdz3OchSn97KAsr5Am45BFvyOMykuFcfQSc2lLhj1351AoHw0
mhKQej5FNv8KVEDr6+8/RUpNUvA9WhBMCRnkK2IP2h+V2aASFgNvQ88b1RKisGEc2IsX5NJbpIcZ
2Jhj3dHAkAwb9zp5k1qKSpxC31OZfFQ3kkfqkeiv5w0FI8CqtW9R1x7tmJydAx3SGnYfIbYcnjqq
zOCkqg0/01y4aH2skO40GfXGZcY+PdWrRBo2+BkP8POWTGsRexYaVHF3hd+GrsWP4DU5OPcqsZB5
o8LMj6XNpN4M5as6/1e6Ltct56A8Bx4S1NYmRY3zncUshSXpKR1Z9FOGzi33peR3Zq5uOA9Lrl+H
NrdQdO8lfxLpoBU5JmF+RdBTcM0ju7SoL/ymRYJk8bd0Muo9iymYkwsmUz1aXJuSiRWJ8Dg8s3Il
pe0MrAm/0RlbDnNaw5tW12zCmlHbvvmz4GSOnGjMPD344OCP1O80mDYiugy9d+EjreiLCSdIf3kR
lbUTRuMKV1jiCyVMNainYijiKDMdSAjwqm/JzCVCNX5SFHqJLHK/o+w7FtzLl2FOCy6GJ1zHbJBJ
gDfRvBxuLsbPXoMQkIY/87o+y1u6SMmgfVXBMv/zdk1/HUfKPAqbM4/CyTKGHePNAjAh7qIeCI9L
2X8ZgJUUA5oIeIi8X+2ZkoPP/Ten2Dy2lNBjZS7aZRybjQCn/Iu3CsNSjCExI8daFdybPFmphcz+
xZeOxw6oQ3mS7xOjtXTY2BYXYGDfbvapp+OsbKtqhJMdh/G13RnbQ+Yf8v9twDOHwxsOenNcwnCv
Ry6Xm65QxAhdWHz0ipO9DqiRb2LOW24083IsWRhjP7rSd7odvkf/Eec+sptqsflKgYBcSZO2A3WQ
gub7yVs9b5Ut1i6OJoAvkPvfuu0JEi7WaO2ClfSdsTK0DQW9bFOsOZRRnK6gQ5Pp3BGXAnBiWahK
9Pf9nSLn3fU/zT7Am7jLotAPio9zaf1vX7/KlSxKxJqEVTI6tyHukrZL6491KYXfF0yoVih7wv0m
ksFGfzn5/IPnCDbaLTAH4fweZNEyFqtfV4Mkt1OQSqhgv1BRdAsDoudbS2w1NdoAz6gT68qlROkK
3+z69KFB72r9IZMFnmnvxPUPchiTIrC4VeL49frVHQv+uamsmteHww/eLReMQ3g7ezQPbDKsAPee
zfWo0OSl21U9d3ONNQSK+IwiSr/HnoF3pJsblreKqZqAKPIJ96xb7giz1zGwezNC9flQrQRR8FZy
BTbetWhqLJJWRFNW89zgH3fTD/JkwZzsbbDdc0/yY2szMSwzEvwMKZPTPRTDqlJQGBwnS0aEDbWu
JDGGFzcPUni44vezBOJI72x6FAiJ1VX5h0Jh1VeEpiBro4Zz7rgnNGczsV/LkNTAhgYC9HsiRwcM
FRZFaJt/lc6zxKPQYc8ZIJ7GbY6U9yK7cJw+ohatHdgD26DFG1aF0Z6gR03NApVnnL1+nqUgYaVK
VKTiJVcexx4u1T4gmrbGRohTixkyRoY75cQaTNlQku4y15tOTN7ch30q0MJEUj5svNIJJ+AgAYAa
vqxr1TJ4WypHcMRYb8mYe3HdQB+GMGjm8ob8dYjSJBcZu8UH9ALyyAZUCW3+6bh+aQVNaF1TOG/V
CrBLswmPgd6MgaPYiXemCEI4ovlsU49k7LP8VqnpQzb6vCE/LfWArcGRq/Y5VqjSyO2l3+vzRsoN
za/kcI9hkRFtjv6Hw66bu7MGEIvIvTAIrX1ytNeFlrDepazDz43KWzD17yUDuLkeFH0ZvULDS4SF
mu73exp/6osBYPqW4UdccJIw7zm6NJks9SsHaf3Uby+Y51dYuG6PIPIkvp3cEc9JM4JqYy7ddNVF
SZCLBtKEuyjbNDX8109Feyv0yYj5az8wuBSvGfQdhXSxrrjK0EVwpL4aTgdxNYPVDbdSNxcg2lx5
6fdo21pIqtN93xIkyBCMOzeBn99bh6ry7qa2n4OTQiStUbt1oBx97+AVOSrC6k0HXnlnpNfAhSRP
v8QJXkxZoOyo8/J3x1tPlnm/hPujalxCSXzgV8NE8ZTZrXzOCaILV5dWDpq86OkjRpBAeMxUYAtk
Vz5WfJzgxz36eJ2Vhpg6EOmUxXqTGoP6FSaSUFMkQoU3fSSs2CPAp0JF5GR+G+g8l6weU0bDdcMF
NQs2D1PtlzWeMoPSNfcYWbaa18E0NE/MiGKyyJ/0Y8YoEoEChO6AIqQU6f6TmjolzDke4xWSo8PY
6/3JqYkxbCW3ClLP+ASEepE7AcN377cjsjUmwmYONf+AJp2S2HSPgUBjyDaw+SpEKusFKLeFjLBt
yaVli5X1of19A0eT0wjp8lYmLO8YCrj2AlqxbMMCDHRFEKBSxJKCYOK6Qpwl82AYf05L89I8CZbH
aYtV82rhefY57V7bC+gkJ2b5VTHsSWcsO1wM5xKacfW8qrbg5jLEQpOox2ocr8WSffcJWZAp/SO0
cojDUTYoW1wGfswaElFbuWuLSmFyRwl1peDgUfWbNwufjASb1ZR1j5QmM+OLfkE65STp7M+S9uZX
E0OyDBAhoy50g9Pyj65+I6HBL0pSU/xdQ3hbg9ljNWCGh34AZDwNQ+E1VdCMp53hZHYPz0o5Vx6G
50mSrZJxBxlFVVsKqR6fg9X0Q2UneJf6P3CjTr4iLdBMxc/9DRPxhyicqPa9ptnndoKSVhHnW5Xe
nUq9jIyl6AQmf8eFc4GDtqd31kzVBIMBq4hVcssiClNjj2QGIZBRvGUoCBP4j6k1UcywbJiklf/9
NMYBg6kDDicjAmnP4Sru1gmCaKpwmqmf2s8bd7wJ8BswKhELWbFNtKA0HhobnVShGkmUFoh90C52
ezy1GQJ9DM5f4oek+v/sh0zuaSMgrQipoJWdSWOUkWa4z03enoGhO8zfXl1en7CERIMbwAyyomyo
bPYGjt0QaF4sRVhyiGHzNhbf9vbhFAjtxPe/tck67NmbfPiGOZrjj5iDRuSisf86uqwzrbRAxbX6
U/UW8CvQmHtDyVFp+16iAhPcGHSOqMhz6ltVk7cEh1ooxAyt79fuyNYlVdH9coJQJgZbIdSKTjVT
JU3MXdF2RaKJsw9DZBQRHk1dkC4vnzG/lGO1ZBpb9GSVVZSb/dDNNKGje0BtkGGyaWvQfdOBXhVY
wrZjkOM0QZnNlVCSUHqnReYZdx7S5v+lpa6z851zINjowor3M5xhHDGhuxQosXpfsz7vBej5EWzk
2c2mNKLyuQToDeJr5dTsT0K1GHfNvBxpRxBs3KJ61eyDfsdLOm1H9DH+jPdheq454qQ9S7SNFxaH
s4y4e4IWciw1diMdzIi/XCeiNQ9olJW4HlPXDKffzL6dAnY9L8kiPycZJbrGWQfLd2fMxUGcSJns
56+tIsPYyzEDuMzgdL3WbpVOgjA0278kI9A8rIF5nolrZQIkTx+LjXkpjK8RW5AjMbnNdSKh4e6s
dz36qa26k537Iz1GodCf67AcqvOHgP5cZmgP6rElnls+8CIlSdnCLBDOPytQktgWyMxuIs5x38LN
0ODzm99EjDc+IuG2i7keR0ffB5X/ct6P68xpCVFaIZ0mVE1MbXfRxiQiRnkegUkN/oQkrG1xf+vk
icztVs2Suo/CJRo2cQvIUwhIUVbIeHLNj01PK7dpaoE3kG/Tch7iYHbBkhdwC9UWs0BAyNE/9lSO
kz81WWdiOP14vsYo+389mwfE70K3/hTOhuonNJJUEPsNs87wkne0u9WaWYgRPCLvLsh7KwE5oxXC
70+q5kN00yVTAxmgb6raN8A/IU2yWv9TAcc7U1xTqCiqlVCy+rjYk3Q4LpEWU3rv0ym0JmPL/m3H
Hksta5w4YVF0cC0k8vDTUHafur2mLfoUtDM4+vvPWM7Ck9cVg5fFfs2K8jIBA2CkEK7RDTq+FC2E
AMOOT85t/eML+9ohnSGkgytF4/tP8Rwnj190FrG+zhRWhj+eAx7j7tlOUabHVZU6lMgE8muKRy1z
VAwAEO8S48F2sKjQZGrvKL7u2qr1uHNCqh6yr+RnHSeX7M6DWSlt5HWDCJijMUB2cnKdLOtgKMXj
Ay6wiySlyRb8gW+GAVZo33ntV97+ZUOx+ks0tjWdo3/6MC6sDPNI7LK1gRzOO0eucMof6jv0pXAD
3VBnbsrxGKGeZjNUVlZB0h/mumGCKgFVjg6Bfc1jZkI4hu84tJOnQSLgjmNZEf6hjmtxS+KDTmXZ
vuS/wq3TlqQxoxj8xEhVdsbrSlwhPy61dzejPxX847B4/MNalTK7R7i/oXj6UuIedZEK2EfMuylM
5iyHAIJBIX0j+ViOkMNVYWz5vqJ8o2xs1CvY9478Hv6RaaaFAGEsKtXGD+QEdSz6QznGwWipxfNE
uPTBItFZFogmtJLXt4L089bHe14Uj3kglBcmhhpdrcqGbirp89by5tGOz1E8X7VPaz/aajdsC38u
LZ3JNaUhDMVfx1ob5mU4Qg15AhFdRp8p1xX/X7LeJBxhCok5ruW6eWaCAoy45u+5L1KPEngZEkKm
u8Z5rA3uf45qH8Pub45PmVhIQZkXD/cga+NArZkVESW00JFUzW5fbgmYGymkI8CzkNWu1x5C7pT6
ECgus7HmGZya3wwyTLen23QQpkRPEchFdkS8w6apDDQhO1GZ+/CMf0Q/EddRvYCsiEF30Ge3sd/c
lAaXotko/pG5bopgTkxalHmFDJolFEuUEiUvQ9CYpBBR78JZyAkDiq36RH7rg7Y6qyDqc0Ksix4t
w7bpgRYx6cPEw1VWqfcqmO9IHS+zSWaHaCirqH6YTxy83K+x3wXhiPskKuGJjhglU3hhN6/ylbva
JiinW8IQX8wIR8stQeGNJ3EE+LiDntWlGL/nIglaMsjZkEKeu10JJdWrLs1kCKla2dFCPndtf9dq
ZOJU04yj2lcq+TRpYo4lGbdJWo9Km98NyxHxuBnYSPTc0fmysSPF4EDX0u4w09VF+C0U7vM66u2P
1CKAfm4bAe1Dd/eyucAcs+K4SXOsZG4mQmKotzzEqvgJVESncx1D5fjViiQcWlYe6tWSjzgfoLfb
y/VERVcgHBngJSArk1Dg8mRl/1uwkqNbt5Vql3Fn0Gy5lEpjhvsXWYW9cS6y+ki1bUqWCM1ePxB4
bUQC+83jV2egGhh9t+JDpzKo92MpTborZOhAlFVjFLB52Si/5VKH0tI5peBwJEwWrQ+HGccKlNoQ
4LqY+/Km21reEkb+IgxxUHjXrgUfshjBjfTM7GKjRnchr3FBvnUhbtDqMrn0s4wr15a7FHpq7QZ1
a9VXgnVseoK9UKBPkNptj/+/Pak5/LpixUCTIy2A+/FklFfjh/7wscESOW/Zc7fcSgXVFQq6bbjQ
f8BqyzMOrWol4TIf/+++dsH7zHURXG13w1EUnw2OR91M8/h+Avse2/ofEcZv9avuktLjlk3cqsL8
sZiUGwmcPzr+Lfh2sdBOWUxjSLLue4FcOpzONM/ISUFiwPvX5PTNi+6sHOTVeH43g5ETHVIWzROC
jlzaYShBJGCTnga5IH70Ct1pb8N2dr3nHN6K7u6vZPFVGbYbwZyOtm62Lm2CMve3equBBWK8mlIC
w3z/cGP7v+F3MK8o+5Bycth4HaCfMPtC/0SrSIylmaKgr8PrefzwEB087kXs8x8R2uTj06TWAvB+
ZHNHpKIX4e9nc5MqzVPaOSgDxBYSOjSVSsXAMW3IE6M8/66cmxmPbgzjTXIaDRrLEwD+PHHkvvtZ
gCk+8z21QqVOjRBYV0rZRbsSLBqbAQr/SdXhsGxkZTUhy4SwrOzrtmrw+rQHRzYe+VkC2a1G1Web
oraGx1eDRFwadUWoXtbVzNXLbqOOnP4sgiZWnpJyrLTbxGtFyviSQGtz6inOe21OPJ08+N0XV4tS
Yw6NebnD0n+rwCUq2T/+wSTrIizax3Hqq3ia34KvApyV83eB6/S1gKNlZ43FjCQP8MHO2G6c/tl3
ODhGMQWwRjnu5jMOBfQGMu2x1YIroSC2wHn7krej2GGTVu4RRpKsmxmmjh+NczCSgh7oGti+ji5x
Feaj1hPQBtnNoXYAsHMiZzZig7mAI6Ks825A9/ypziceeNARTSBt1pWIWrv7lbbEqt8FgjqDKg4t
eWAY+B5GrNj9iYkYvUtB6aB0Pel2F/B9HID60KhpzmEyxtOPRzERYfOHM1bZIcPAiApBDKpU44CJ
lMCVXR8D9DPqonv6Xkv1CIlRduz2Yk7mKU+I3SCzDTXcdP6NaQ6+Zgfl/khe5JAxeboTYEe2jyFF
wtvV6ozvF5o2/fOMKQBofW6Nl/I8VqVZamQPwj5XlOy8U3W5JLmBiEtJvwX0mfLqp7YN/pJWbI6p
znn+3BKVSSmQuPgp3IN0u/wCg4FVC0IulWQz3L3uE5Js0J81Q4cPTarEYw279fSD51o3qvli3+TB
LpTXETdqhDvFNSBUILobT62yc4Jh03g3VhyQi22pPrcj+xaHzt/WmGvuZ/sIXKzIshpxJJeDZaxM
H966vCUBB/iWyEhCSY8lUTdxADel6Xjn7DsGU33ZqmBITfAl7wOzPguX4O/SNIPZnu+ULdRNE+D+
eRH87xQTDQV9Pm/MRTOscuV3cYHPsR3Ou9mOW8p7v6P6mhlrqdXLhfCWosGE9IW/jXuiYBCFTOhH
82/Hj4JwTdWmLRzF6Fc4n/jox4AC2ycNuhb1B1c6pqThOoD4cN1RnXOSRYTjZfGyd5ZJX4OnagrH
jcqOQAMtDSxHAQq7LnzFiVdMNyKM7g66udprLY6GioJ2NOsFjMhLvYyjGE/y3h/s+89wAdkmNouc
Hjcbgec7IqVFmCwtulKz4PncczTJfceRCw4fxlD/Vc2zpckyIW62+OANsMnC3PqkBX2RpJD5aDAc
qJN23GEELY5yozMgeDfcr8YC82k6xF9ahrs5FIaPF+kv3H/NgD06KVFdpQkvUnFLPG1d33/79RQu
5syClCcxwp1oQW/31bkl9Af1MH1NEQHgz0rphzcr1RCdbmuRymK3njbFzngMuIGhmFOMhNjkM7BC
5a7uIySMnpd+fQ6ExrIm0tpE/ql4jwlMtvxFC4S7hqR48krK5Sj9BYP/GCO5FzIpurU4zWz41wzQ
xwCacAEbo1cBlXGUOi8cfvh1VR0IcgrOMg9l7tu0pmunkkCqiJ2iyUK8t4pE3qwGCybA17mpcUXw
TTs7YRjMD9e/tXbXNAm05lUhgVFSpVYUGTh3PtqcUWhCWnnnZ6plgCOgPTJjnQ/kXWuFruAdU2lm
PoXLdF+Cr6BoIqyorqVTA1a+rB7oN4tn81i5IdP5aZenhxtvYMialg9PS8UVCNv6X23GQjJxGFPz
fVfFEok7Syef7JYU2QpXvp8IjbzlHCl1vfHqdfVKnV/zE8z+dIohNNVkWrxTV3ny7GUf/AVRyHfu
2Qf2jUTpt/SijvhOm3IUlb1FIHuU2wuhzbQ+Ky7GU591vON2hy9sa7iRkgf8KCvDmaDqWzJqj/0w
Q9xEy2srkQRuuGPU2R4VFRgMPxPa3Z6+0anf31XYccNbWtAY2fOaSjgMiLkkMPExNsigidG/xrKe
1CGYcjPxshfcDYtVkjxivaFKJTTRwwh+ao/OgyRED3yzYY+khGemI4Kwztd3JW7jEhUAHRGZSUAK
i05sW8zO8hwOWe5Lft155kiOTQQvb3obEVASBSq/pyySCV4Pr/J3+hZEDC+DvlBv6X0hB7bJew5e
rTHxHw/S58HNKLUR3PMt3eXbYjYUcA0+APl9P3A18d4aW9v9fEaKzEqsCUTYrBKOrWRPfM8tP5ob
IynewPMs0RpNwz2laxAdCQjpbUx6UT788xY6/a4iagmNP54hbvpqndRPBFDNyCsjRzZZbH5cY6oo
rK/Nwk6Vf7SsTepMaLJskm8xb9c/Lx8rbuuSIEJJsi/MgbQgoxi2/SmBALmsQK0bWG6Q8VRRPMDm
1jytmujXoTDWYC61Oc+JGFda0mXT7Se9FJcELZwz4OZL0Ac/D6oTkbuMYiSfrD6oHIR8ywofN4Dj
EztxnpCVYqof6UTV4Zzr1P24ftMhx5oN03MjysJrCMq+Tgh4eS1edPODk66W1+MKQHROsubLiti6
Ld6BliM6BRD7xiFsE4ORzbwCxxP9Vlon3qmQlZATDPRiInuhxywM+RfwyX6nEVRkwcJ1R1EfSdWd
aFonafc4CGODqSwykcAmKtoChs494KcIhoNbAriVSSob3bYbV/ym/Jt8kidQO7uHa7puR35A1lkH
/9QHBro1VSnC4qa4L5+i2ddazH1G8FWuSMWwi2HrE+tE2ihgj5MJdpl3pDcKN1frrGU/OXyALV6C
pyJ8+lzeQJGgqJqbHMxoG9hwZYYtwPSUfcR1xSmrfydKY+c2RRtqBDavvLQFZMRbFKpo6JKSRqPj
fniC9nS34i+dNXi/9pSi6PRa1suLOI9rGQdQsa3qg4lyAdpB4RLTumiRrSP2GAoiA5r1OXkOswGJ
KmYLwhgTXYnDgqvo5N4JyDA1yiLaFxJoOfVmcHA5ydcli+ZVQGg/AWfQ4keVCyGaA7TMHp3yjVpE
bGcV32B0hrTPjAuAGtVsj3ALzq6imq3PrjVPAMKchr4rfYn46dCe6uJ4ddCo9iwkvL98RuVCvRKH
jflA56tfuNmxdNyF5GB6EvbqIBaZ31tLZtiGcMmuuC1yChKFEWWSHPwRYEQTXM1XR3GuoKeunE05
OmIF/fmJ0eEF/vtgk2s7oH9tBEO38JDV5Cr5Uvb3mLW/g41yqG7zkhM84OYOY704VnK85fjnUu8h
tnK7kjRsaFu6acZ6lbtz/Xe7mAAnM0Qpk78KfNEvR7BwGDf2YNbFWgBkkR7zl48Zwn0IznJcQi9w
R4u3fSwxXUMGol2Xt4VvJqAkjrsx3sdgNGCOkN1YqVTMSHjQnRuykmeWgkHfwDwcPqxf2ReiygK0
8N55nhdyD6FUEwn76KGheNi3zsPBaOpoIVPMbfzMDQoFwdoR07T+EC5wnbc1S6/qcZmdAIUO3j3d
GhLreBaayp3G3EF3PDnv72taIWd3lv8m42iI+0aMe6IWYKoOnIJwbDDLhITzNm84zaK12AYLNO91
gCFZkk+W06ce+uuXphrNs68T3wGGQ8BBcfafLuja7aQLC0dd9GDGFQjIooWZ7LC6C1dKqyXf81e6
UaXZMlVE+aam4jAtbNIGFNgB1ZWZLTCvqz/bAFn54weXxFTCJTABQbTZEuSC+HU+/9G6mDbgml7N
Idn6HeeBFc50fAIiBHr49eyJQ3bXKC9OXsoMlle+a7I7nvU4sGyNuWv/wf0goT/DSp5X1TJkfEES
NmOtVdwQT8TG6JTNlqB9c3AgHA7XoDFlFnjcY2+T4lzIwfmtmkdE4L5sjIDwdqfQYxJRvoxlkWM5
lHXsKNyuCycec06F1sgyP5Xu0WMjiQrSE0WS+iS+8tLS87mBgtSWbPIPL+NmWYwiJSiQ/orH0P8s
aXpRf2oQf/W6aZ1FULJe3DYT2n2KxOBcy4Sm0/WJRe3xDDYz1SpDfxb4iyRVogJHvb44aFvr1rvI
jeSVMdDldZqUq7lMl/TJ/Y/nnEEvmF1INyQa0EgUy+CKUeXIFUFaD570Yep4D5LZqO1iV27sMOQ3
YkilXEkDEIi+EIyOXlEZjthXqc5vwF/XT+9/3OOcAgTzbdyO4EFyOYvj1T88OLnB9cYhn5Rqfzrk
EOgUYGicEJncwhSxWbTIFFgvNbgwTYAwPb56vOqGnxuONT4zHfCHQzwl2a3e7XeBIjJyOQTkv6Qg
ysQfonV8VDge/VUUm/ic0tXXHHH/FfBOVJHSkPisUv7oF/MQgsP6qTwgbRgJhF0c/ga46IHKFp/4
XwRDdBRMRhwMi9YjzRA6kdjeFuLbHj5njRYmBZ4w1ZPiP9/Bsv4X9MYP7HstcWkAeFurym+aSIvS
wE/A/xYo1Z5AKoxGWG1X6J0XmnO4jCjGwhnnd3JZyXNz99lU6GQAtK/hlzRhSJFnGB0pw/IFE+Nn
5kBqJ7MGahb1ptQwLJF+ZqtBpwwn1NCi7QLRCK2rqaaUeWfByxyCFtNftY3qTf2c7matWMhoFNd6
eFDlLl+YZnlfEGwAlVBLlyOApmXPra1WtF699dbWuSD7Dwhc+x/4lmv3B1nAi1NPWIc+0rrLVJoC
TxmCJXcaNzvkN6W9qzVyd/XAwY9c1oQ+PShUsSCwn9VYih1YkFoAjbSuKOdrlk/E4wxRwz4Zqhgi
bKmIIQjc/i1VArFpkDGIzLz/yM1LmS3/KHZzI1nK8WHIH2RpqjayU4VTLZtvloCkZfZ/EkuIsGBE
f/NEIR6TIGFk4xLn3ggHyMuy62akgQgqtHtekyl84VTLzKtNqOimQh6ZsVdLZbfrgKhhLG18nGc7
zBybJYu3x6toCND+tp1j4iBR+YngBfoxhpYV5tpiwr3SjBhtdK1RfiatPNQ9/FrrfR8mNhr4fMwV
s+nEVCHsXn1MytlP2IMdaX0/hnocYnfVFqwBizXUu70SQwfrQYI4sSvVQyS1e74GoI217FB0uQw9
QObjvUBxQ1n8vd3FbNQiloBgpkDyIb1O0WKZTNxJsbvhsbZEH5M3rMvSiuPfcrvJIEVATvbzFkPR
MCCNja2YG+fAcFVPH65YyvSnepKHigXU50T+qp6u31pJxxKMPOTbkgjeoy02/tlw/rgEgeZ3WWyW
Hm3TPhryFlqn4XYkW5GU7mvsC71Pz2ElJCM8xwbxGc3DdUeO+vrS27jtkbs753x/8r0tDfCNTor9
M6MuXBdR+PDM2kaMQEzue4Jizr1z+Im47fNISdOx4ZUGh+vL7IK7Jnmo8H2lqZX+FFAaAwBuWPmy
CNq9zGt74pWLWqtmPVVgUXKKYmcFgr3JuT+xUjWKyn5IpyrPe7hpO0MKRdnWCdT+dn51MDYuDsA4
ZrrIdZWIW2G2ODswAQfn+95FtQIq8RG6T7iz3W/RSwpaVyXADVIqj14+5BPpC4WLuajbcrecC719
mJDObWk6DoSugNJrXml2TcY1YodFNbqh9PIDK2TK3rk6k1UB0jh0ArClPLBYPL2U36WhpiQmmSgI
2nk7qHLK455uNYYDqNl7jGFiTCZEsP5jeduIhdbA+oTU5Dx8zfzRz0pLFseMFbHQGFvnrqfdRV1x
gPJz+85Jp7yYcbZkEX85122Hfc1xSPcp2KxfM2n7hIYBYunkCO1w7iMIKpv/cDmWhPdHaWj4iOy2
WLg+vMS2lsIlSZuDMqmYNaSfz2nx1vi/tlp6zserjho5bqCy1obaJ1noAYQNDG9j9YUL/KkthgKD
qv1ZnKA+MK+13TlISNftIu+5r/2fbIdMkp+3nN+x/gTlzOnZLbSiTf4OQH5ob57B5mocU/1eH9y9
cxQu7cWR8uEBxE/SPlorvAQt6L03WwKlG9k8Gx0+W23Gl/vSsOKryJ1MHtmF8AU2AiDGipyv4Lki
abV/KNasYh3i87cDxKSVNyAxt+Dn5vK7lqYhA5PfEYleJuuSfFRmOQcvkRnJdXsi1ZqyCpQS7WvV
kA3w6wI3gGSLi1Mv4bCWIW0wlM81eVtwwVyDaim2h7Bnh6ksb7DHhUG39k3AxPdrLn5RSQcwr3uK
zl07ScopOXN5kMQ72cmDJ/Io1321N6+J/blxI0TO0OA1FT2RKsiyC5nU7EpGYk88hc6SBIhKWNR/
Ppr7gjqadtFQRxYn6nCzTD/hyX/zlMCFdsNFetK/DaTP/oozKTlsxw1CsHPOVDoiweZP+xWXpUKN
MaoxwEnMUWT5Clf/P2iUYNtaVD9gHPHbYuPjbSwo0EQqElAMn9w+F8+vqlxp8x0v6IVYeP197yoN
zvtL2dEVuoGxwPQQ4wp49mBn7vUH8oljgefeoUCNAaZgXTuBdBBrD1IlAVEF28smhVyRO0VcWRMJ
qtQx8mO6LOM7JHSn9Jdumf6cTGreJkhizpjg1XFvowepG4J9cwbLeLBu+Jx3/0LiHRdaNB1BSJLX
78ZTAQ3KY8l44ITa92vVee6/Suh+bO7HKs85LQsvg1rUiZwVrbDIRpFYHBeAcIsx/PflRCjkc87y
yt1x0RTX6Gsup2omhEi108J3LpX6jRT+xnh7Aqz2CKmjMt61qQvOR7v8jyEBLdrKMfi9tkPCxfcV
iB64wflUrGT05+7PhIM8T7tHJsX5bQI5aDL9F5wGskNDemtY2CRNdqfxkuZBonap6wYOSd1x3yj4
Fg+CYR3vR4ePzZgoQ+w+4gBbjTfxvvhsoXiCiEhyEpQWZ29cWoNgg+6HHW4zy9ul6S/w2feR+w8x
Idd+N/cf+OPXOJuIQzHI4Py/FaOmmHjHhUDSJHdZE+mCT8QPdY3EhePgXe+3jfvRBjk8itX++SAc
I3IThVDy0DDOdqBbcwi00nfZLxEuc20bnlxiTm5IP29/lzrtIP8i55U4SVoljxSxjYKKv/FKzFJZ
/Iz8R+ulsafW2t1YJnx2Z6nehVJgFuBhLxvb+pIeB8M8fUvUULBUK/w4v3xBj9kmx9Y4XB1qArjZ
/M6CVF9H7zeht8ONRK1SjyEIcsVdR90iezjwq6E1VNydEBMCTh7EQLkYQ348xIi0gq2RvrQt8LGd
aot03tbGoqn7UxtTa2DD8G99L25Il+JbOpafz/CtVgtzf2sQJualchLGFeDX71TjEau/EDqXYN4Z
gimGcWKOaVcy6O60j2kZT1gRFvuuQzVSYa9hP6rIqcMADvlN3yeMxREkSulLJKvFCfzquhxR+sYX
65i89EwmqGxQaPo0Xnl9XuMG2cr9we89ccxw87WCwkhvSGrjAJgZHzwzYJ4swEu7uvwZcILceM0u
/TzTRdv+rX47JesmmXJpdHpi2WpFxjUr2hAJQ+PMmq2LsXHe7W6bx90tWBahOd2F9IyZxhA6jR4A
vkxKAUew+v/OhPbxydiDTG0edMY8l4zcpHS2+qO+PlrkiqiqCZeOtlm7FWwzk67mVimS5pmZVMHC
gt5uwyDxlBgYpz3lb5AoHqk2NQsW4Aud4ZOSFRI4+HzLxF+kGho3Gb60ktHs+a70nXWO2wiJ2g5D
QCusBB1LxUCsHv2r6sdcKU/ykrOIOb6N7cme0lOkZstElWt3MWDIypX2HHVrh+8sUPdxdp2XmcE7
8vx90frgBswqtK2i+5K1LHvL5bRMICT29E6P2fNurJKQY1BUGRFNYwbX94fUcdy4f905hbdXm4SF
nZ//Z7N0W57ZjQucYTGjtnSA/dcMgER5bUQ9Ug+b3OA4/5v/bdCn4OkvFAL5OVB1jmAr4rUSB/oX
h+LgrtX0HfwrSxiKT3ZRUcBCfvbiHphV6laSy2MPpw1jqsUSipVNAe/42q3LlfaoQrOfY7dTHIxJ
qEoCH4WY4Np2M6G7XLPzevzp7chMmChNFfupiK5sonzRIPVml1Ah/iLaxm54XHugWnccC7Mzxd4G
Y6sJxtrO08HuZ5Uw+Zje5nfrMGAtEN1iJ9Pjg/sYBH2fiPSF/b4Q2eNM+axfEGBmBPpCWxj6qw4b
mYhv3z6DFrxHHXTdNxOok15KJa9UL+uJeRsL7GxgJ+uA/zpEvKQ9isPI3lBtVxId91PQF2XClRJN
n2vlbFH47qxmCFNxuRNz8mZQIn8E4+15Nak+cW2gdr23g7UWvv4US96eqS7jLnCEQO+19cCymaEp
sebuZvGL0pXw6sg8yS8Z1+pSe9MXfS7XgvbER1MO1NR2Qpcla37Z6q7SaOfcgAxMMGwW3mFH8qca
s78GVAYgsXlD+hgpduJHn9mfc8iGU57067IBhxBFvze0aLGcLEo6PnIx0JPAEctSOxdcYRMUa+Un
zI3O9P2oQNvtWBFnoCVE/rer4tWaFnQ9VTd6MWHOB1fV0YkmzTN2XlYaj4WSZlxMfx68iiVP0XXV
JxLuisDF4RElmaF05b0WaR0S1Mvhw8nVb4fnthDmFBqLGML+2sPTCoc87s8JC6WmHPiXDcMtfeJ4
uwA/xMCkSkResGNx/UHgvIO8P+qNiMSQQyBw8Rgjg4WDvEabzw/sYZ58A1Xmh7kZjP54fK1y9fR2
9HqXobAg38HTPJNTOvY+ms5yfp6eff2PoqmCQs9fXe++s4FZqm/KvSFaTI9BqrzNkw/YN0gttQJ2
rCJqza8Q8u7RVZ8LGorZV7x1uuKc52vc8jOrvYvDwbTptxh9fU/wzmVa1SoOqTndMzEUaaMnTFc/
ldv6Ga6TBMOTJPlWu/antgtawSGCKf0/rAVLZP3USzECwG8bJHqcA2fpcAfWMMwftrcwnN2k+Md0
N95EvVyGLN4c2WMnLzrXlfxnR6YB4KFuAOyDeg4+1qz1408deXM8YuHdzDbNXWbKp6ZZ8uJyE8UZ
kcTmDfl4tahd+BmfnSn04jm2GEs4kcIxth804qN+oIHfrvMwj3bpU0l9gTP0lJDMqkLPu+iH9qbO
bw5kE/ujLWWzzB7zCwZkxrOIIV/UH9Nw8jE8H6VwtPPxCgu1fIp4JTI4qASS4wnI09sP4mEqpCNc
gVWNSw+Xm/7lO25pAa3FjU7ax9Km9I8POzvRWFvCr+xkXjywKPN5GmsZdloBaYcE0sy1IG7Gb5eY
lofyH2akRTVdZpnaVwIEdTxMOvzSMuoj+rQfQBtBUZRPO2Mozw6WNa8aDxuJpZ+fNIf0g5ZLdQ4s
HRA1y0H2L/lS5uLzwmSCn+TltDbni9s8OZWxln4+1495ri8wWx1LlC1Ber1rJ+5YWfKugSvAzO8f
36OyUyETYEIKbSg9GI/9+DpHk8TU928E8/KwUFFaq0zHk9bApoUZywpKmNePP1mq4E5dypeVPQTl
quHJ0Hpw0x26y1OhYlVhewOPC9lKaXOUDaiJPtCXCSr9JborO0NAzAX7FvPH01nqkHe0+bBXnxl7
Zbelkj8TKVxb199Dp19sqQqWSky4p3sKv4DP/8IOLgzS/h2ou2/P6lq/ripzm0j4k0SyuD1KgCO2
T+8R9QljKnBElGDcqiD4So9RrCI2gCLElgr1qnltWo+s5qbiDGM9uSuYRhed/mXQ2auAqyPW/oia
/t/6cvhoWfIm4jYa+yMFPl+FYGU8PT6AtqpCuyWHQEm7cvaquQ0xeF0zAAKi9beDLbdWxSA8+Kxm
lLEExLpTCKXffV2Pv4iZkdXeF/4cJaDcN9UA5mj81fwucfx9rFINauXJAP1grI45015sXIW4n3sj
itS5rHDObGj1X/38PZ6cAly9ga15KtEhwuck9JSs6gXvGD//WxkdHK/8uH3bDdCSrq+AsjQErZKI
4d30INb4pbIECmWU9OBniHvvKPt3Xhd+IliR/jtiHnDbSPP0SDDLCRcCtySynkii4yQ1uQYfckEy
ttOOckddhbAPVZ4QFhYQxRpA8QI3JBkg9cdHGQS+1gmF9JjvtN5vN5nBn1vc40u5jN41HNHtu+OT
GGeARiSyeqkRLd8L4hPlHvuFxY48D7wjZUvg3yxgTJZAeSW5g8T1zVGejKaxi5iX4eIE4Oh4hc02
sxjP+TisRWoLhoqHk/JksD1eRoxabBtAyuD+4CcVQpuTcNuBpdpdWWJFg+J42lxMphJswDR5CmBn
DdqdYB85wfJTJ09eRQEL8V3PPlH0t1n+4YfYIHEfG9yz63yZ9LuUldGTukvE2DLEt+4pDxcTCbYp
0H4ECho9x8W2zPIMVFYZ9V9RAi9Qup+en2e7+X/Bp4n8keV6CUzZ1eMcCpYCx8jTveys0u8+KzjA
Y0JqWciR4KoHu7beHyJtallSJyXUe/DiswUSsx9JRXqAmQzjM2bd9t9ZCgDXQ1AQBbG7fTnbChKT
4iYZJUrgHVwHwkYQtArqIWkvMjnDMan+FN7C6sw0tchOGMtXkoETYKukdclBj9DhOQeMUUwdXA7E
4vHMlEtkpleEiL8+hNfUI3nPmWh3HnVmqvSAYFLLVuLdbv3ClosGsD4ozYuAoVUkPdPcfNWQqnRG
3XrULRD/htbrfqd3bXM7lJJdi6UG4YnmxoWxwcnodP4Eo6NzclnAC58117/vM+VXvAUIBawWrN3J
Wy1wsc9dlZKuOAUP2rqz3zeGy3e3QYyPGbSECcg9BabKkRgUF2B8wY+H/+UkxMJrv6d+QroMiHNl
ma8jaZtES5wYeBL+wSPaDl3JswHQ//qCB6A7/eH7u7MT77D6ttTzj9xHqAcEJ8QK0rRI2SpO6Pt9
MyhEZXDvkdj5226SJTUH8JwiwenqI2uJrhGwjmfAW7SZmTYTV5qXGKuy054SWGhahy2wt0IJ0KlF
qM/XjrU28xAljOGtIkgU7njONSuznzT65F83eIf4O3hj2dVcMY0UyZtFWrg9dNKeciapj4lXM0Eh
KOWkFk3vYeZy93JNvLxVVwmEnOkhJfl3+sd2NbDBDQs83NW9tNEulXxjz/kJ3Wdkha4DaPP/q6Eq
drDdFLW+TzCtVLk/NmCIBH4lPspkWZPBuqTEhYrqSmT7HrPJOvPTAEW7d8dke++cimbmFGgZlxVr
vYPLj1Ipy16G4HE8QzJG296O4e11voBw471jius0M1/oA+bsGlr9nUmhY0j9dG/0/n6bvM7qO4CH
OeiWu8JMZethtmhR36C7yadza5hr8lBw6VPdrQAlfq1Y3bH/QtxtBJSpr4JkjTTqa7UZSL5sRpAG
RZaVNyNeJB7CHz4kUcpM3SDofLzd+NtR/yfBynaE9PwgOYsihFtCzfuxzbwCZ6REAP0Ph4oT6KSG
ZC0lkmZCePFdANOnq3cZVaAYM508H+9dbghLt4+Rb6d0IJBuVEQKVc2axiAzQv1vHRuBSuJm4yZU
P/LFGgvH5Mh9ZNU1Ys98IqYopiPyeK5dwmJCfaDM6/KZOSi6JNF1tRAH0xeRqgrv2xcuTRcrsotJ
fsyTijEKZKSIBsDV2rrmJG38DacNiCTIBlHiOUat4yqmgZeUJHJvmyw3zrky6JzL+g3qilQRjvW6
QZFvTybAm/I0XfS5A/55qcGxWkKap6xZ6xWRTutda6svVLTGhrWT0V1nULqrFXpoSMTRFdM6ItUM
tjnHM1jRaZ8/vGaPSrRazjRL+yhLyEygAiJM8E63TevMrSCvfr9wGhy3HBuqq2w8E0I3iEkRLNVs
chno8+o3xG+qjzlRFoaWK/gFnaBEdB09Q3t2kQG9RA4Sq+qV8B+5YWu2fvzbfSjLDSSBarOdTsvZ
K3taUVn1xbeSFJMKvwJhMtRJ+2riFPvdbaOt+48V29epoohpEyqZgypSdI1ViYcc+igQq+hH5sFW
T+ETyCQQwbf1UTbqXLPrlyWp8lhGvthn6xIZb3Mxo3aOSb0zbUF+PHXzudKLk5qgwUjq0+1TRCYC
uzDtgbSzjMdKYxTg0BH94gEPwwusw4CSmg1IiNptM33wd79Ui3OkLe2kmL562/qz1KcdVsaWOD0S
mh+l6QpT+ih4cBAo1YFoxjwi2z+Yyg2bikhW3nN8ELNkV7Sza05aExbwMWXeB8MFOER7nVrUOSQz
KPMj1dNaPRtXzZglUhY8klnxkiDoB3V3H/2du/mRTdfP1FMje4pXs3IvsAhag5WSU8NfF4tAHpDG
ZOF/oEiS4hevmq9ATBeV9NsIXyMR+nWwUOJYeZOuKKthn6F4UmDPOBLxS6iHQzpzI+/RfvfK55cB
6BnTTm3Xb5Y/FVGGqclpbhhK8LV7zo18hZwS9kTg79AY+De2G6zzR6kk5QEn8kLxQ9xsK1AJRTbL
OcUfAy/9KktZIFCjJOmtVQeg+gx8rYWUJuG99sGtbzPBkzQZ8Ex+VXC8dCUp3RJIGbFoI32/rvmL
oEMzYjsD2UtXkZMCl/Cx5FZrgbhM7CPf9ibGOuAmw0xOLsjqQCLmxys1xR9BnmOoIGwCzq7NWlzl
se22EjxMrx2iCgzq4xz1e5CsKtki/HbK/yBcbjT3HUApFXzocY6Ms/UbU2O5zFq5yyGuWu4lN+q+
amj/HLfqRp3VjpVYE/b32ZAoko17D3ofJNa32IEvvQ7Ro01j5HebPnYKvC/icwzzXSs8rkL+IMkS
neMUNkvOingsfPFJ8RNqj0WVP4asaYvREydNCfFui82UyLcXtFjor5gSVPsmtGo/WsCfUS5xvM7S
R8U4HPrSolpD/PI0tOokXbkTAYxlGGUixz6vjg0TJ2Y2zvfF4M0CSnsSTNBGrihRpBZHYuxG4inP
J5Hs2rzpxZXDvgsznRCFO3neVnZ02195EHtrSopGGTHhqLks7sTg5Ed4gjJTkK0fU/SReP1waX49
leuocxCdDw0OBzKTgZcdKDGwb1POlghv6PEouB2kbzOaKVvZhuqgwQ3fq1f3VTSVYjoUuAuzktdW
XXup7wxewqeXE71FEZB7vNaQCdYSNZp+JNpifiRlBl+kpCbqfaa6QH+QHAx5LtgGoE4wyYGsJyJi
p6SesqE5PMGDAtsWj5rD8/x1qX7hpi5Ks+o2v+cZluRWNp6sP5dQS9dm552w5l25ZGHFlC2D96U4
8aNaba2SgNcJIVV/ypsC9cN6DBdqGCoYyX00YK/fqW1SZ7jQYx9QKHyI4r06jMsTaIJHhuJUGpXq
Ly0TyKpVTmR3oMhGRcYLQpmh3Fpj3Y7ik/pFczbaaGz9EwctGG1iZXoMs4rJS+P0CjzrBChBq3CD
pOm2JY8kJP7fkHYQZARVLYzomA5a/BkvE9OSRlitxgjuJcWjr9JKHAWwYvgkAKpLxK7jkpg/PPpT
BKE61Y2GgrgQSR2JKXoq6d5DyYJ8gji1KlrCjU6ssl1GLaL9pepaLeQG9Yg+jRBYsz/tFo9ioR1C
5DABA1iLAtWjKz+Zlmp5SZ7rWJh1XaPIhQfXQbDH/0HzG1Sb2jtO/g54UweYElqd4HJ4IhaZl1WP
D/1RYv31FDFHPYzi5+OO+vW6+LGF2t4rWLI04E6sXBgX5u8zlP93AoY63CzUPsl3n+5Hdx5jyEQh
h5qNSZDOn4b7kZUfrMq6vZRHKPFLvrNibihzOz/m7rdj+uRyyy4C6qQg5wCBulTcwAtTClUAadgK
XiUga6VX6TR+UuJbcip6rRcxQyvCltnSUfFp2DdRS7fCo/I7YbQoScVRq8N9xecnMQoPanLinoxy
S4gKf4y9rvbuQpeT29SVBTbJAQxzdSVxd9UNOmPQypGm2lhD40Xmp208DNLx2YujhQM4cimSmEti
/f7cR88zDt1IJk3npiN4ephppFcMch7zuDRlN2xUEMzpnpBNSflbNiMtt1wga75R4eSSnieEQ5Jc
PtHaTFqgVoAmmKJq99E+mRaJtpLepFSi5Tjdb2M1bxZyeTDp3AEuSzSMLn7qqxnGyHbHbNX9FIa1
5dI5rq5wRYUP2AN9qYtAx9jLeq/plCA/vNQJKfSm6K0x+5QdDphSM1UUGtgXUIGgFDqCBkkyFNeQ
MReF/Ib9uGWxWZI1SBT1zIforvTue5sYxOGqDbl9Xenys2GaHq73OpRdyMSuovQ9YYiuumU+BYGw
xae3/hiYxanBWzQzqE22WUi0y1QyK4yQ960EeL4JnOeNmzQZYjqaYn2i8tu+X/JI/oRwurFacOoM
YUfF2WjS/ipLZBICk8g15Wj9b43GvEnYb+ggFgUY31+B09VNCH9EMi29ZFk/UuSVoS0ILhIG0ZOi
6adF/F4clvoxP3IDxvwIHdPgEG2Wd8BQl0j0KpLhCOSgO3ahhN5DuCP2SOiiUvX1GrXMe7EKR9WN
NCzFcSN1rUVIkvaOaV9/14tKYD8dYCCnIX4JnEsN0YKgaJ/VRDZOZnyNllyYSmM4CRrf7rZY6cz/
zfY1FPksEmUrmsyZ6613fGTCsu9kSgkpTrdfwVJYpGmrWqNTKwn8ziRHjnc6XoYFcxpyM07/bOAF
L12GDaCY43JpRyqvytLWf3jgO3wi/eQV5jpCFnR6hDML0ZKa9nP1evLiPj5Rzf1d5muWooyDeo2S
GnntFMgBONa1M5KGBTaetANSCvyByY22vyDma4BPUfJZqLFThwbxfKIUEDbmAP/5LwwMrCn2HsgE
66qg2dijsUNUZQrASJl3zwSCtEE3eIAmBqY820teXsu+b/PnnA2CIxDTjkegqTQonRS52K62cJtb
ytw784aosV/KOUW7wPxP7oc4cUXRb8CZ8iYmrESO0AJ5zo5dzSAsKYXocx3Eikogy8qVyrmPDPI+
iyL72NKiBOCv+4w08o7yVWIsSGO64L6fuhgIvEn48GfMZUsP/HKuV26Eee60/P+YTNhiZlA5rIEj
2Kn7ge/nfRBODY1qf72FEH/iAGvnq3BZsGZbqwlyvqpVoepJLhHhq8UxTzX4922v/2Qu/0XCuxre
TqUQHYp4vGv4GN+OVV4U8iMuG3h/XRCsGXzwV2n7iITfnKjQqiMMw+5fMrEOikWduE3eFmcD+cR0
fNVTCb4xDHdkNW+mkLqWsJqLxjpSpxbz9vfICN0/IP5JH7HGm/JoiMTXMVwli30svVYOwjqusXwH
ipjrDzQ0vM5Sphz9OeqPZLA9oiqRRboC53wwSG87PhXUjDZZmquXfW5EDVNBr+vLdoTQj8Dh56RN
B4ByKogCGYEtee6voFv8Fi5hG79HwvZOgEzcdegfVfr3qQKwCh7h5bHEjT8DYyozWPo5AoVDMXBd
1D6nmCCCYelj6mHBWwBYfCWeC/Ub7EoA8YNq2dvj2uwxlkWXW1y123crm0BFgaqEZez3kGfZ/TdE
b/51n+bCf+a2LdMp3n0WZNnveB3AbiwUwZ3wtDpPLtfyyDDGmXQTiplBIAdt5yEn5UCtBi5DXTI5
TPZ0dMgOUWhneXyJTbM5nHEAyN2DfcKUdhADrVhwkfvXGisdBiHNw0IDMuuCkSKsIHKOseVLS5bb
Z145SkfI3nlYmNqsGIIihYGaHKZoeyRoCPOlqnDcPw1RQgX34NLSA+iLdOfkuQlAshIbfdMlkved
ncDBprbhbX89vOXnfgTN6cTqUneDpg7OW0FNYF6WXMF+WYkkmeqSmeSBB6S+kuuSC9+n0Bm5wXWc
GEXuA2hFDYYDtpUuoGTQ8S2P/qLhxSw0qSYBw2iOy2usQ2i37sBkQeKht44ywgaqnITiT9GZD2jY
pyLAawfEzlJq17wq0Qos29md9jcEV5Wz+Trx/uepkFOMEWZMKk3IS10fxEPbmh/QPQ8a2Q5ZFAMu
qzLjUMA4qgvGiAdZTrhVOSMpdZM5IBj4tN+ChQxD1LfyLPTyIiruMaOh9tpBNMwvEm9QI6BiEwql
j3c/Dyqkb3fe0XjvBN3DvFidDDqL+0calBCNa6TfqBDc39lykJWMKMo4ajuFomlmt56477idKT7x
kU/n0ilZWa+Of1e6ZxjCnIftyN+7tgVCB3/ZRaORVvGW7hTBwoC0wEaVPSlI7XazciFcm+fwCOcX
md9ElFoKIq+AyD0TuBe8Gj9bGfipTszatljYy8eX8G/UYij6pglL8IVXugUNzDTiCL+2fqydKNdR
/HN9B59S5ISyAShUsd7B/wOtXNWDKvDKkF+KCiEelwtuKFgJ40zA2xdcv+7rmtlZiuo5OIawPfAf
AyKA+KNZsNt6gqR60ZGtfi2jTdXRoriiY0EmpiqOKcQkhGfJ+2QTGjeWEaYKFjQx8cT1+7NLnXI+
mPQHJ1Hg54oN2xaqpigCj1s1+yrUzDtCucf/rGyPkXeJRw0c1k35LJsve1KREdTFWw7fueNgYVip
B7pfhOkvPSBMFDmJnA2OrPlGwv+WRyxYIfL4bmCHYsqgcLGv5Aoxljg1AAWo1bn4ASK9bjtxncSK
/0vA7tiR1K9M7Wt5//qaQP/an22byETB83V4bBpbSSN1P0lwP4Z8cPyJZUqNd86f8i/pT7crtuBJ
WT91x8Ee47EYJMFv4Ek6zFpMCKvbzOx+OrNhkgHf4YROPiERPdHmoyZ57SIXFJpqIhF9EiaY6Nu0
mbouEciJ7MHjlVvi0Lto4pJ2aJktDenSlGxdCEKqy5/SjikvmA2iOiXBeclgK1CVwaM+6cEGAvkS
8CUnkwklx+XRWZIr2wdmlv+mZZy0HbIyw+YK0u646kHJDmNGJQxrJ5NEHJpTvVLHfUCSnfAsu7uk
W9Z0yfkY20wtdPTxsHgIRAkixhl6uucEJe8HMF/9gEovdWDnVge1VJCFE2H8GP4nB55cUIfuAKvq
/TOLgQcvVlAA7VuH/4eAEpSyOk0V6RFPUtrJbUgywDSFy9fjioCS4Iu2qjoqF3vLiV2pwiNwuWj/
zPtCXchRiY4iIDBQ7uJ6tWltzy6XUsX3Xgt0rM+ryIMa4X8y/QkW92ktd4Fi9PEzPGZbni0/FILc
8XxgQ4WevbCvBe0LsjgH/biwhUzLfYr2T6qg+b44tyF/IxQhIvW4DFjCAe+WtAd5S1iVrND+igGp
MtghuAdU5YfwmpQ0KgV9goaFTZD9YhZZzvpdOWFs8FsjDknbCjsbqNhCE7+OG/VWOfOcnVEMgqiP
AmHOFukEf7nSjvNcsJ3UYAdPSm696TIyNzJ9mcyPg4kwxZ689xIKp2DVjdYRVL3U9xz0RR05T8OE
K6IdgNy5wZxVm15MZCxNZu1uqxtEEl54kCSY3it8DprYdAmiuedsxZDN84gHV7Z4TsrrTA2+v31o
NOGNKwyM7M0iVmbLJ2OJjrKpi3aJpqhGWhRyjI8IPRuCCx+0XuVaBlK8+vxwvCISDF/9j24DqxAJ
iMfapy13r8hcXHoFqoYau2T09riBvj0D7f0xdREdi24N009U/wEAvuJpWkQTXDZuaW12LjHdUar/
Khp1A8V6M0HO7OlFigeUGmEpI6BlJS+yTWAW8rKy/p8OX+4HwWID1r5ZlByU1JP50+G/FjwQK3oc
sEmrW8XFwxASHwpv4jlJUG9CIJQ2rqBK3jBKdBVK2ZgXnKAzNtkicohShaogP7Dd2O0XaqcmjoPT
Evtu/40Op9H6JCLK4O/lBkv9aVbT6JSwAaEN4//Q6yanv6wtJKoRn4SJ/CTOmqUA/lXrMr9SIfhV
SBQjospmJctc8bEJ2+I3uQ5FWGafaforbZ1DCT8NOs1dF5nhTnzRyqF7GzqFtSEPm5HPD91y+NPW
nOWG8eF2kK8eiNU4LOBE6lYubYJQwQirTztB6pJfN4TuXvx9WbAU73uVeNoibFuWtajSMH05ai8O
Yagci/UwYyBLWe2ZuGGB+Ch/7T15GNEuKXUhTLRNE2nnnuPHST8JbVBnwRpe8sWMST8O4G3Qjpke
eprFlGQIYdBdQTkxcaub4yZKInGwb27Tjbx35DyhIxeHdXDeJU0RQxbLVSeuyWh9vnhIr2lLCHD5
8rkdp5Wn4lFkdiMV+pVanzcjQdu+FsmOaoQPPAoVFUrtFRsowV4o41NOUB4FG+CGlVz/SBL1sDSB
1q3Ze3Xpq0R+H8baKupzIz2eQFIw9mGfkQ4PqyFjD+Pq8+Bb0463e086iLx2iJaAD4e7JjlrjF8g
1iAZryslXPooFYjE5qT42HjqvIVKZ5724YLPIGxDRdBUzMsTGLeQfqmEC1ymJcIc6Fg2NnRW9bos
LbTyvpvLKEQdo9/Y1/Ug9A3vJC3bHkYGFLlo1il0Snu0qXJGzPIjMRtwripq9XVgVUh+KAGQ1d+M
qRIriLg6+r5ozAEg7V9hfOD9vaashJZtBwbL8gg3R7hP8YscXg5wmLcmSWEr+M/c4wgfXjEZs01X
EP4+ERoL4WpHOqG+uuCS6FvfDsC6Ka1yo0U3ireQAZq6sufidbaJjW/aLo2fBYUh6oIBxg/VSERB
hMSzKzF/ocbr0CyGyrmYWTDD8cid0NkkJSEo4rbWbLuNS0vwnYxujzoZA1rfVI4c8FqxaGi4STij
EmFoUZT26p0iNmpvaQuZeBOxiEAGOldybo3GpIAZjnkklxKmoVV1d+BNuKx1Uspwh4hs+dGkQ/18
tvaLgeSTts0MhdI9geS2JkMI/Sfcfju9xcLvPi+gYaKqSjExzerrdzmUR5NbST3k7XmvUaHBsZrA
EFOshLIGlU58CBqZDOJV6bRs6ZnXhxpaw+GUhP9xKMDG8NqFRMxlhn0ub8QqtN9j3w61XqoeIJsT
6WP41PP9hVV8bSvaEYAROogp7mjUWvPQVlqP9Mql3qTDtKsa2IOQoE5rWeryEDon0wHiJ0gADw+U
vhm/LqtEZ9lWXFnCu6BNKAYmMGdkBSLWrdp93xDw7Aiik2M9uoKQpMpZXitqPQAnz+RgEvSkbpgZ
urlHzzKrBczTzi7ixCd0FlZFTfmDH09nGV4wcxRk7LDctietBJ+JA4NPVNNFHzB60mrwFxHok7pN
kjfxa2EK4YResiPqsGPIT5CGuBhXyjvTSnrGdBb1mkme0A96C5UaevLd54Wpo8jyEUx1266h4419
we9X4RBBzblaMb3x+C2eQUdZOJCihRG8b+TlgM+lSXiDYs04F2+RWjXeocdtEQa2cXNDVvkUp4v/
pKT95JFV2I/8O/kl3SFIUvh76pzRCEQTomiveAXlTXIXF8YULNUOBQAM8O8ejnUkk8BIemvFsKMc
pUnA7H8zgZYeZI8qGTDGZZ7hJQbGujePAO4y77KHHPz3iexJX5h0+drP/3T+FRbFE13y04dfq2qd
mlTI88aGk2eitujEgXAfs7CAdcRaIoSZgCdfRQ6yGs1ysFkysUw3ThsXJIvg1vl9cAPgltUQ3Umb
okCeI8Mx7OYxOSkE8Y7gcSoNEES9Ug4ZF80Sncyi5q1Wa7SObffnOtTiwOo519rJL0zNzRDgI1/w
Ce4tc1kMTmUtsQ0MlfImGHJSYO7yfjE4hF2OPU4+qAH8QQK/AZpshS9fOvbsGl3N6UiNthwsPpIA
OvxtGZlktztWOpQ3Tp+ahnZ+yPhnf9QtuC0O54GcndfNax7K+A0j3OVlCK4LD1v0/OqGS8sBowYh
4WRn/yklfTcCZKKdnu7sFREmri39JkrhSFozCmPIoX2rVflXuVLguvos6U7kzN+p7jtdBEatR6He
BuUBr/ReWY92BuboqtABV06jVQk7vWlORnpeBxQlzCFgPt8HIckfokaGZ1pUtkhsNAmXQf2X19+Z
PFjotOWe8+/qliFmHwCjgxlVeS4lxfGahTtWMydAwO+O6rLtWUmH2PqBKGnu0bfcndt3ug7ldWa4
0zrIGzR7l9P2duE1Ghvy0w0owbr+GgXMDYWl6326r/WU35ikPCTCUSIX1B0QKDdB2VB3H/lDCBT4
bebM/94G2dZjOLPJQRB1fGq7tqoZI0tgylwnf7Ny7QX9lcf7FHE3weUKJkJCyErV+7gZivqWOAVl
SvZZVo01PtKnxZQ6T+23o4MYgt8JuU1g0TQFdxXTUibeFZMJB0l1JlEwDNzy8CY2m1d5RycQl9W9
U/ObcgT6nzX9TLZt+0CSW5UhjcAoMYI+nvkbwNRzsh2SrGRUbxA1tzCKv101o5pOzlwQAilO8k00
X2JolfG+/uv3NAZ/AwVfsuhP0E8nSRV0vI+SdSxoKDAiskmutHo/UMdqHFLhqd2j8ASZH1llHue2
mk1PzDNDg8Xt5V0uEFvnOhU2af1VolCGdXla0t873IyJah99x5aAauAwsUHPjTxA4HTBLGtBjbz2
omZS/Q1VMURlGe2fOwjLN2QY8FDGATIKLtfk5Tg1bBOR6TaRXdfdRe/Uw2fo02jvialcAYWbxnBO
mq94pANgLoyqUpehSx6d80F2eaQK+eLfsmKxh8SBis6zhzVdUcBxn27EN6eQshsyxPVNZGsFr7Ul
fgInbCe/xo1M8A/iyruh5f23OGVjsGzAxzeJn9bWdiAdrR26Jx9BiKsVlHMBX9NyZqXWGepaYPQ1
UCDTfWPnAuHxHu6HkEsH++M+AxE9i2nw7SQLhwEbvAczbfBlW23uqjOs6pHmhwb17u7in92NDQ3a
jVK0qA8kYun2Dr3fluARcy8xWAqxvy2ziu3oV31V9Mzdd8rlA23GGmQ4EG4qOE6M+F4NJIY69MfU
RxYCuDen0yK8depqUhvetpARa3AzADonOPIxXN/GmZ+C4XftvmJqtMS5bYqEbAZ/LbyJIkkRnoYw
R+EqlRYsW7pW1E6XTrgi0jFsVkkfE0vXw1hwuAA1Pe+OEnj+Nwg0f0OtGPlCGS7L5KFCDr8mteff
awu0RYKM6ILB7okO2b2fq2sbDEZSDVj3xvAD0VLnzmuKC2GhSvcSj4IySjsActhzAHWrAfIi9Mcr
Zk9GgVgCePmiqoQX9a45q9hCiDsTuKONVI2Z3Ssl/OZVh71it2hMqPZvQn94v9rczYU8ThuP4+lN
LusDIZmC8jNgJuoknc1LGFAcen7zvEuZ7cRB5zmJZWJH08t+c1RBmqRerT2fxgn+YJRgogusJTKo
OVhx+4hzM8wVVTLr3TcpvTq+PpGNk5ciffmiMtci9eoCkZ9T4bdNx6YgGzUDaTBA0z8theYVCOPE
QHCE9/gvgnxvJAnSjcbtwPwdPnNiRnMZ8IPI1tqjnBwwueP24N9BAuLcSBZnQxNY3AMnLgyD6fAk
BXCiT0i1QbXpiYURZJDdqfXYgKW8XKYBVVGOZBivH3bm2GzUP+6rco7e593rm4IsvpQnNUrlA4Xi
cZneOhenQxQBRVkgFzAKr5rDGf1sfcVIkXbZIamtDAH96Pxoy17HvALsatZmPZa/wr5H1jT1PBDG
BoslK0LRPeerOOL1tE8YftrjMiOJBp7hK5ZozH4/67QRcvhuR/63d4gKAab/eGPQ23hq2wZO2sVp
bE9A5MkgRI0hlNlU9VgRu0fDAaxNptPWXWeoMN6xfQOWH/nuy9TqG4IZCKuY6xMTJQn7w39MqMR3
DWulyZS4eTo0Tvp6zAg/8F2kom8kl41YiQfVqjTYPpFb/fw8nbU/826li30WzfA6d2CNZYCbR9Wx
FRSahLyGTOU9EBSX8b7sNp48k6r4zOgpytGr/6NfnwxrJmZ262PZYCRFmy4KmAdr5mBPnxQy8pE1
iPn3b+SalvW8MQkZjX6iyk2vF8f7fEIEehOX2gR7ZOPdg0lyW/GjRYp+GuustEKMvCptHP1evNa2
j3VSJB4W+ZcEk2NCsyoqW0U3maYLGTHEDCHF7X77bq9l+kL/vbX7+JtkJlFBfoJDdA6SxF/TT3Ak
3xnbr8a/S/9iKndSCqH/42Sv487w8CxV71uW82C8XXJra/iHM5raKEaHFsbsDTMkmTsJ2OyAKf1h
dFDCZnDNPC9T7gbex50b0yWS+doAN889Og4hNl/TSFLpgCbsnliXPVMJZ2hTPFfDtD+xgDqXcoOS
iidiNU8hRBPxwDOwF/qtGTr9UQAEdFgUD+fF6h2UPorzi+w16FqfL4IWx5eVT/8lox74+Qoc9HYG
f78OUBO04cWcfv2Ka/ptpb19qyHmg7JoNDEyqxKhcYSpzpJ4aMci34LqHod6YzWSFc2WWwCCCjFi
OeyCpHNKbDnlPEVxLRvxtTv/vNMt/r9c4+kemLQMEfBiLy9aFlU+juwCPqc7CSOtRDbjzJjWNSCw
rTZGvxkqfL7CBAy3fTTNnnzDlumkOKgl9ItAlsAGcYb+eIODhD4xIIb+qg+gkrvW9/VpI49Z+m/+
o2flcH1rDApk6oezUUYm4P7YlNVZlcSMWXVNOsm9dr+J2lYSBDMYL9939V83NqhjQzKTdGqP02bb
9DLXqlFw5P6brnLZlLP1sWWirhPxcntJjeAVs+WI6BmHM+zapOPVFvQL1R1sZv6s399NRNgu96Km
ImE/U4SWXFeq1vo+PqOVNeTENRn3BU/VC4rl7TIE2TNLTm7jnNXOaDc+8d2hA7ANB+tnDaeD/mnj
bTVL1//fIuc5CHBOhxvUvbuAhjsEOa+IHaO8ROj5TkDSfzQn81rQe8rbd+qH5ujUEucPnGAdSv++
xbHuAaeytu/fxh2D5Cq5mbIGj82lljOCfKhrH/1AZmv2j8WkPajUNIQz1ZaEGj7GaYhOL3R+WeoB
vKBzONfznuGPP7Tblkr2Hg73F+NXMHtrPHNhDFOyWzEDT3WvLcZUEe7bnBCHJ34sY9bBPtsxmqWm
j+ojuqGKmrxDI/PUbNXX0Sp7dv/wliDwWK/oT7qrrRJ4+HsJRQPflb4zgBitfxJqbCftL05ykA26
akKv0h4zlzycEiYWNmX6dcg98M+Vf1SC9gf0zwsvlFDp2sjRgH+v1B7eg8yJFuRQFtA8aPslY8Yw
PWtdg/SRzw4SoRndDSHAKv0Jxg+rQkavw1ZcLtSrvyYVLO/nx00+PYorhMOiALzNDNxvxcz8dJKc
IYZMnFPH169YNX5/mocoTXhtCs3WfsZsWRjPej6J7zVe2UdBTfX2vcuoRRXHI3ywa1Kp0/yoBOvZ
67rb+oLtsdfZq1vcTAihASL4B0Qj0c44CDXVmY4EzpWr3pIYg6EKtMPgVb3oPrg1acWpxozVK6DK
yflh6qHl1fslPRieCOETF0n6sBu8XXoYcK3sKZHafEM16aMg9Ln4gH1JrzoacwAvRZtcwcIoenu4
5guo5vM7jXVHsqz8Ed+10W4MIuucO89HpHpgFoMKXkI+7sno1Dx4n/ra4SiubqBxIV8KCB2udOrg
E0dsh22nZtp1gG/yTynu/BHdDBr5JFMpxiOo5MMyCH0w42C0aXwvUJM1domaWa3ozaQrLrHgvlhg
wU3XwAO5iY8WBxR0i+kEE93UBfPeHqC9406e4Bl40Vc4kMrZmMWGjxR7n0H7yeyQrmBrRTzeTglp
qSgck0wU3Qy2kkE6p4jfvk5AqwYwkMtVWl4dkSH6JBDpvu0GWza2sdN9RqWFBmXKzcEsVPfGy83b
8ObOnE1zg5MqiNwXxh4dBMgx/oQA/M6iNNe6h2LL7jRDG7GhFFBBfPzhMLuIq7fdYM2mvyw7NUSb
KZ8DbOsY7ThpWvLuWxppBISEzfK1kg40jdj1mPgfHOv/j3WSnEhGp0Zh6b21N5MX6LppUf1nCHRC
m57b1bvnQN3qGO1SZf4yMVwkKNJqk3CMGYpt7gl979bbwspYQikp5eQNrY7/+wtg9aFP6rjbhm1j
IABhPl/G2uBBunHaTLYxFaGMd+n+fo0V1ITNaPuotH6E1GM7qJPekHbQemIwhse6+7IYOHU5nhJV
BtjBtXOb4eNPsLMCx4bKi8NJrFynXWve3OLNhNS3c2nOSl+5fqOddry0NWbGnQ2md3IcFE5qIx0Z
v9gknHdeRXP4LyZVt/1mRIRNEmZRG66YRJHJ7WXUudeYBDL5UTTjNo+mhOTmwRHzjpv7+nfXh6HP
6NnJ7ymdxb6prFzmxeyWm5APRA7sIvrYdJSpgFvwQbOQdHUzquIoNEJWSlwguwTtrDbG8Tm74ZZG
+fuPFaBGrp/gA37lACTYiwOHC6iZvgd+UKxwG/SLW1hVACku63DGou/paMCkqNydGtd4/1GdOvmM
0B+6hR/1PpENzzcNGrAGRhGot/r1NyFDvUk2TBMyV7WVDNa4gcbX9p5jdRsK6N1hS4q4I8RaqYLo
8ZDcfQGK2JRPF4ST8Y54YA24xglI0t+GJNWiufUc6UCuOyXe+k4fvoMENUlUDrwAglAaQe5hYnXu
dh4n6/xV+kcJytwm6gJR54iGebhEUENrKbnh7gftH9HwTFVaeDBQ+qxPyhM4iT19EUO3xYnf4KsQ
T+MyrEqFCX8NhD+Zv/HTfAqVjUcGOPYuQD9lctzQxz1Fu94NiLxp7yoD/BtJAYopQ0w0tHd/NhPU
4cg20gMTLtH248PXkl1Qvx4PzyR8+obq2O5vIpJYrOtMvDx79fWca9DrZvALJHQ9np6bYWsdbyEy
s3xtAyT6tpcu13doe000lIDIoXLrwAB6zIThj2gAclyKGcZQX8grQKPtaU6AWJWhSG/LtBf8aEmo
irH+ji/TRs+A63nNEcdUS6rnte1HZm9zlABz/2+/tKlf7P+7Tf2/+A2CbwnMA0N0p2F2mO7ye2ov
tpAp4GVXNf1QeK55glHwh7zQkeHWMp9PHbCrY9fwBgey3zzKtAanuX619uMZ315fGf+u0mO4Ng7D
wFJT0z9OmBSZCv6kDEW7jfVQ/ijYDaKXqKpynUN0+XJvcgjyyH6f+ff1UAZgLa6NLAmZnqV1w6Ns
sVJy4PaanpHIh9wvVQWSSrr22PMe0OtX8qF1dSy1Bq12veRYUyLhmE9uRgnUndkVxv6gqak4XOb7
2IpAzL8xUKMMNt/WaQL9V/vT0rjtAHcg96KzpcunD09s7CRpCbKThffqRYj6cU9xHU+7qtPLvlNF
wblwuJMu7bpIgYd/XeQcKGEvnB0QbYXhHQ5+4qb47zBM79wB6YkM3Kquq5DMQKnzHgnW4c5IXmve
7XoaK4Z34NAGOrozquVMPkurZ4Y97kC5eY0+BRUEybpWT7vtxB4eWA8/GrNI0KUnGvmGqoRnCVbH
so0CT6SZVPxULfLRLmN+YM3ES3hwEO+yTkKNq96nMgNdpe/jmmIlk1wtqAiJOh7SyggmwGSVptT4
xLDQnG/qrYm1rymbzWEyzbSIT9EsLFERFrLWUw1Yx0Y25A85ou/Hk69V26mbWrgUC5cOal6Q9FC+
ED+DVENE24e98VgIiYmT48GqXTYk+Hdkn+QgQaJjSBwmorxnCjIlMXCrV+bnBh0b7SBIQOcu/KIE
3sYLT3cE8yeC1odIDPqc8NfS5dHB3fSek+LBpGg3w17bBmY9oZGnDnrjc6Qoqnc0EsFukE+82jEh
9/6c/U5VqMbwQ2Va7C5VRUUntxIKuGEu02FStBYW25e+a1ppQwZg14i4H3GFkSlYp7a643kRqCRZ
duVqD1qQ9PDjKZzgRrsJxY/vbOr8UMSNTuaVOmgBM1a7u/Lh8e5g1mK2CHoY+58q036nZSrfcDIh
lJjh+h7mnM/8MOjBxosFZiHBriPdgcdIsK+jgy+eI+OxGtY87x9wNTji2HmjL/dh3tT0EdU3VgGW
/CnC/gHZfFHiZcQvu1k4hOAyCAMulrxcNOFkF2VCwz3Fvmi9cMcvFrW/k7SERIUYW7r/6+TzAKMa
SRFYOwmGpw+xOaL1fpPzsYPLauftCz9Xomcqzb3wqb8f2IdWpXx72M6F78ctfnfB4kwc3dwcfAuO
rNHyklwglPyuEs1yPjBdaUc1bFW4U3vWYz0X3TCMTJGqDTYdbN/7emqa+H66nC7BF9ENpvHXIv7k
wtYx5RLqfvRYxlURru1+9cfL0W0TMIQqyG1prCft3Fbe5pca/+WBi4p9+0ZZ37L7g3+8cbVDqc9K
45zS0qiQ1O5CEjM7sEFhKlM8J9rrSxZJUQ4Hf0PS67/owApWOUqIRJT55bqDVT/Fd/fbmjNP2GqE
6Vz69GnmVI1OVJteJeK7bonZ39e1emkuf5Iy0AEO8pyax0GSFZU82pLslcJES2zZo5HB0HIP4Qin
cLzrE3Ni6acr3/JTlf/0X2RrhAyWJSU6WrXgOEUICXpNUOCPfZHEiugpnckPb6cT0UXEW8Mo2PCw
wqs6F4ql0bxlwWDCcBD/m6D8POih8HSUq5sLv4P4vc1q12+AWVhM6kLSwA2DzFRLNYs4M9XR0pfW
SU6PuSA7qwbZZdWYHdGelu35eRsCKGqgrOMgV1aog4Rme8v6x95oWLUZpzu0kUit9g++HKSxfpRU
HUqtfXHK4paw81Y5GzhR+OgkZ2PYv1ifxWVFPmDsrTNL98YNgBz5N+nyDPohIKSdSRPDrlEjT49L
qC9umtXQA7eJ1fV83GyqNPi7AKJWQOvaWmuorvwF0+Nr0uKriy0RLqzmgcd6ETAEa8utS4YBNdYL
0RTvmeUbSj+jVlBva39kGvM0u4zntvRXjFOdIvXSvSbpb+edLmIZVBj05g2OmfszIiK+kNP6tvUq
+QdSReIV3OcVxdrFBHDeeKcBIC7iA/phdOdPX+mIiB/yv45rBGWQ4+R2YjPfvasqSSlo7DfhJ24M
RF4LkFwrr88Qhm+M51JmOBnWi60PqEQaYK8j8iT61WgrBz7JRWtmhYogQcBX1Ah5xkYzOyaUEwrC
NSgu9KQL9JEs/S8rjq5itYjmqfnuAbQfxyiwrhfu/AD6QxTDxqUqs3sq9mc9XliNc/qpYeOm/69a
T1v+6ly61V3DnVVEaYz4flcrcRJSZmZXHpXAXFkvIleTPikvZtG70g1STKSrmuuFteITw2+fjcnA
Lw53LeaWSHpyUbvJQFhV5Kdtc0SxnvqLbPHb3lO+SN7KHE+Br3USR8wD7KoRDtx8dDxqqZtJsXtK
Smj61oq5C7iu2+YKq6JdAyJAVw1zFvcOrfjby1+NfDUqtOyBo6WpyxqiQDPjPnyem11aRVWx0elz
Jrf+fULpdwwvzjZ7HvR6DT/38jPJBYjrVCO9cIgteYWjXIa+0VCQFNUCyU3ZtV0rQrHJZM4TmJOO
joCQw1A3QdGZMUVxRqMWMgVD/1Adt0pM5pFh5QS8yQm06vktxLRWMAIrYz33fVRV7ON0fImB8lNk
9+flCGOZAS9Po+xDelz7tPodkwUBGiMuXjN8wTCXHDsW+O7SFUkDPHqGEVPAYyN0noIzNONJfvfu
xjS0/MRPbEp8kO+rgtyStt6nJasii47i6Z4MAGwKbNACzEXgJyXdpYNDFqTYMyuVfRzt4b0CBpUX
9Ac+S/cqmqMPU+VyQBOx4TKVJfFPeP7iYWTZtxilUdESlqoHrfpJU/t2O+UAdXaWyjzvQAJjSrkB
agY5cuwVcM2+YIbkCVhIyyzG+pfLcbrk20GKKjlmfey8FKVvCJy37O++bua7xphvtEAuGxisb4Ro
rSf+4dtzbpNgdGyw85ZUPNsZgRKM/yF3Tln17e8X4sYkagJ9wCICyRjiThAYlv3+vKkUeHTO1Vzr
cr7a4GOsITl5isaiqFxSRnC9jj9vvOqdx+9qZ5pm10dxhXecdr1dhOpFQAi4vA1Zrw0jUS0qAuL7
VxpgtQg6mWL9wR0MFM2s+F3JTT4nCcUuHk/tUD5KVfgRaGcb8xMyelHRhPQxYfMDoppRHpoiGY0s
qyM/Y2uTXUZI41OHhRosXPM8qpD8ctiqsVotpaCgA6lIuU1I935jvVGaKibdGHF+ulocML4BFO5m
k0x/1K/k7Ev1j8PM5Mprg1AEAXZjmrzpLH7Wp7z8jORRNEh253Lypp9yBRPrPnhijaOkVO4Csf8Q
Aad4fREr7KyHX0yQNO0tVaJbRPXA8T5budtllgqNXLhfFmEqYVVR3EnYDoi+gzLd9lHlRqSAwLet
jAkuuatxrxl/UTJZW7132YISICYDaFzbZrTBfREBUwUfzFqZLO2eww4V7HW9xYvwy6WgPDH+JkXP
Y9z0sVTBQwgHCdoeunwmAfMyTedqsBsC9861IQLg7WWGbZNoDg2dAl/4YtSvab6ZPY9duuvyayP6
eVdOYgp4/oX4d8+Adm2FMC4n8hWwqHUxjhNypmMvcCoGFz/pBcgPZBcvwvMkkofQ+61J1Im0NWmH
BF/ZchcBsd+lLB1/FJ5ugwNB5C1KUrRXiO/+5xSy0tslVlDQKwqF1e10E6FzGOSAr/8be2ksDi0d
uw8xAg3c73XxqbT9PIf1tPq1K2vZryFV/jKL07l61eLADS8DmZUox9mBvla0LRFH45G9/xWOxA/q
RvbvX9DE2UuZWniizFw67jN+GLipVnCNR2xi6KYFvc3MYwAA3raG3IFQVxL2063gh5ZfUwjOvkhH
ohNfSUa6bABuhYJGqqEkiF044WcQFgBpvm4dQ5+3SzUppDTGZJR54qRjVkOOI2RI5AWaKhSwQ43f
BQ9Im/8F/j9grn4P2YgVSI4los/XepDV/XDeDjvWPhMzXwOcHrQsa5q3yfrkvpDeTXzymx4A6BMs
UUc0djuY4Gc7u4wdJbJtt/i6X0J1X4QehwoKuoocvOXE7IPkeS1Bhg3PQZlDw45qXB1zSUWvbK9D
sk1ohIjsK1Jp/lIORrMP0ToLd92NRYakrnMK6D+UD1PAs0jexyxtYT2ewdt9n4iLuUVxL5Cagtr9
2y6spJqx5e10OSwZ7lllfPyyBqtAVt0A0F3wh4KZTLBkj43zbaFLNeXw6oBOrniJCOcNu/HGp3fa
aPDmBAlr/s3KXZ46XxSZ5fZJXqSV3WRT7IAyR/0/6GF8Bd7FTIa91hfq2+nXvTCV8adfPFFWFmFl
APWSHuuO/3DXibKXacM9xrGCKp6wrY+RKZ+DvkWyaORja1AQmv1YhW8hTUNlrwssS/gKFOSWARbf
+sCXl34B0XsW4XTItZh5cnNA0jhE4YAxCX4NWkLN7fs4NVTcAQEdmsbbssxacqntz7X53Dr1fn2O
HwHk2G3GxRmf8reCtORgN18aD/FRKtzSY2Ow+66POQfkkPbwPRHF5PPC3EyODuxGzS4mzNz8uDvE
Ae9yUWPyBpXJwiT3Wr6sVtSonnn2/f+A/DllKWx4YCOuCSz+8n25uPSpUzstLB/kxInhORZ3Nhm+
ZdXvn6BHqUVLIRj3QI4yf1cuo8c/kdBiRuCfkuE2buImf4utGHVYXCv8j3ek9RXYlrQSkMjBnE+6
YvlJTV15PeI9YxE/N5xxVbke/AgNIOu7LTjtLmsdoKqztkUNjbyuAXrp7+9+awLfdV7VyALIHkR1
1g/s58BAvcSII/0aPDuaA8lRbZOuLW4b+cz39ME5jjj5xwngyezpGGPl6M0QyoMoy/Y5i8gfG370
7w2g9rBxzAY4dK/c8eO54Y8h52giBFUUG3NTitxQAC0TR00h1OziAwBggmAK1pFCVvP9Tv30v+v9
YlR3k17jKRUb3JL3MnwAzGP6lB1qbndIEJMhb+2us0t9oXZGrV7t80jd8nMxojRj6D4KlkmppcF+
RR+astWWKhdQj4qk7CwfDEwatGWDVBdvLTjVuQXpMeh2JY7fW/LZPPic1ii7Vtxli6mz6FMKDU4l
ONDMDmcPXmpHSJmkDaQnfrphE/Dc/4OvsTogw/nPskXEFXdoLuIUccmGcdj9/7ie3HRJi8Ux2xI8
iZPCdnZyue55NG0xf6kWXnYGvGP0cumSpbPctTffMNoZOMjcNHgJJzgraSAq3ffQdSuwQ/YvPAuh
wYAe0ZSpqdZQYMXpnRVkIWcFG79Zd0EF+502v17s3W/HHrAq69e4cMAMRHTaTEu8po792beFRni3
MyP2wol3dOdR7COsbTLBp6Hn+dhUpMf9ROyAWyXOIEKJXLdRH0J3EHDh+YeMLmQwtDLxSVBWuXMZ
9zAid2VK8xtm8WXeKPCFRynSRaR1GgjS/9Gyopww3LUjpcigA2xq0Ku6DP8Gq3h7GS74ySl9+SQM
xJVLxhQf6d9ffEccGboleCVKZiSH4i188cOe49bsV/oIg0YpTuNR2d0Bf/uHUyhcxyKKpa391Hi6
o3Ulg9yAlQYVagcgNIlErNR6QOg3WpLXzNfiW/On9L3B8Fmk7lCZB3fWSJiKau8CyGJE49skKyrB
6w1h8QEoeNAlsnlzFwjqlDk4B9RCMxRVblbPDFUlaeU+9Avhu5rK121xeBnMfQcNJYCQivqDVYLy
cbX4WMS4jZCwRJghydHBeDcpgddHhuO8HnVwGIs0469iP76VozrBYBruZTUhA89ZOtuVGYglXFH1
u8JU0HQaw7DWUTZ1Vtm/GMHQqdHS+QuvweEqI70kRxDG1mCLdzwCiPhxNXQxivxrcbrtMONt6VNs
ttQJPdw8pBHho2XI+XBF3kpvz2uE3QsQNoG2Tu3wsBgNMzdqKL2QcHEMOBQ1bI14SXIj0WRtN8Vx
V7kGi+JFbY9/XizTyorkGTCcJHBbPs4CkpFDswuFrRXjYhZxYDer/KuuveEW5zonPpBWLK1r9zAa
s61VJMZ2Nqs/w8IV8r1PsxnEC+A5ETW2xySm1+MEvx2M2ZAToaafxNvFzIXCvWlUepMB+bfTXYLQ
lVf4nqgVhpf3FgFBGJrREGKZq1gpyVkj8uHttazyyV6cOh/0runzfRWFjJjuwnIqaZIVFXlDry+V
uhU81qS8hTs19GxB6UwHcLxPGQND6DkBIx9HfuAZSuIpp6Oak8SUNUcwHGeKH8d3RH0BEPqLJlr3
VvvMduqZIDu1L4e0zcdwiSn+sffa8QjxWpEiNkWonaV5wSV0tVdFBPQdOWYfIcFAXQKdTJN4Rz+r
pTI6eCtiheEtpxoJlZ/cKitrnQmFgFFrpLGpfpN3WsjEH1uCq2r10qxCv7MfpbHWuUJ6lpknaFBd
Euz6Xh391+5GO+ex6wt56UAh8ll+3SsplDNmLAwDln6mga0WqgdvLPXRnS32rmipyHwpVigfW3PR
AHE6CNvNc2X/OAQqY3FVsOaVFrshqf73WkAJUls06TlZQfZZFxMuUryHPCehr2z4y4HhJI2Hh3Yz
Ig9q1aRcHIu7Ru6HgkaGXTXEvE7re0jam9gQmDMNAGs/AMKvi38ONljwTUzRM+0CZbzndXpYHBrG
rft8FK9Ln+VYU8T1i0syYZr4TkcyNKCkhw7La+vJxoVJxKa4JJf9nlz1Oc+bB8Dqu8fWui8aZhS4
54Afe1iFNqdZdd0/L4oTq2bP4Qx5YMI3M9mKsuxzPW5mSqMXJogrciZPySemkDZ6wd3x/oD/kB2a
U1VbPN+PFR8guU1iyKEkvycZdkZZlkCqm1ALXoWp+YDRnIC3nKPcfpTq6YGM25lrlSZyJ/JelLcY
E4dBuqvqz8BcXZ7BfKz2SyJoT1dh5Z8YeVMhDH2sO6PmCDDN9NuGRMnEDxckMHTjYcu2A7FAhy8d
HjlhYlqAsEGkIaa7L7ThPfdoMrOHStcQlIfrqMFIcJJZlbJaaDL+dTX2Q6QQrIVY0v1XGz1QnwCx
YHblpAbq+dMA2IvyhZDd1QDqOPmMCwAY45eSxzu64mLB42wojISqR8z0P/rr+sVy15YxKn1QlHoj
3ZFB+XTPGBVGZqvE/PaJ7H8aCd1ia3XuB8R4as642065llfjt0dHUOn50h50JPd/RGV89pif9aUS
EHcr7Ce5niX2pJ5GTSiXxV6fSAD0QPqBEapEhDIxPLupPFoxTp/HwVWAkU5dTpg5g8iYPDO9ac6r
aOUWw3ZbJgh0XRMVeRFgwPrsvTH4NYpcFqPMa7A3xEAeXGtx+CwlLR+ThO3L6NO6ipK9gTCKfFpT
GRYX9xkftJ9o9gSFKawXviX/35k0G+o8LXLnNjaxCZougLaDqNhc9RGyxuFKRNl3PB+7ViBQhQ6P
UcyKvqmSHq70z+0IbCrMxZhP2+HLVum4IPka9SqO8pnDnqas9olIYbk6AvOC/yHQdS079xIf8Q7F
B+nLjbw1OhSGwcTH5Pu8pZUcAdvgLWDsUtCeQyiQ0+PYO/vlp6SlCxEyMCLrkONZKfnP3kYyB0zE
a2MU+LQv2O25g5veeYO1xgej9wrQy4jpZAxejOOrZWswLtSv2fJKkQyKGSK+fHgoPgDBH4YkqvGc
HVYO6PFTrwKN4BWS/2XpF1fVsFByYqCNfi1cbzyzpHXZJyrAhJ5yO+I1NulDk57JFjihETFvBil6
ywhIVT7d2Kn+Sf9ZW7qj4ySY7E1EDN+7iP22A6UVSxxspguNtzi1I9K+u3xD2v1E4oEGQGqtLjFs
MSlf3Gts0N2mz+Vt0RGrAYnI5gBIhocZWLhOp95OUyNpp5/PpGiUFv6TyZlEXYHVeltwi+ryawxU
Hc4YcGR4wBLP932qsqJ430bNDTaskmFLR7s8o/BjLPkPdj3+vn894czW6NRz0Lt03ai5ntXdhQh9
7LlzDz5qXe2s0S1dWU/kzVhc7WY8l2DAtUBa9FJEt6LDtLO6/JwNXVy6hmGhGfJZWV+/X1w98G0C
jSWE6N70fptfTAuJpgy7M7NmjdO91PCnn5TLMAREDNfLCzEW/Zma7tFahuK2dAgesC7gs2P+OYLt
wglne3simLLtjbW3yQYYdJ1TJORdONZvTaJKAJ3/zeJltdr8UokVAsD98EKWFqT5WvOlMj69/W1q
rXXDWexAE/jDn4JF3ev3/ZbPxJzFiWapfaeGnFB+H1X2emZ7NGLreuoUL2HA7G5sPeJ7SlJX2HuA
kwst1uckACYDEnep7zWDH13116DTJwguYH7chIGInUQa35fPYRmSrdQzzTwH85Xqp6X8gD4fwurd
/OSAS40H34dywyAZ/Te6WwIzpRhXyNUX9H4i1QoPfcLk6HEd2CEpM0zseckzwS9vhHivsYj8DdOh
DtAuXklrgOT0x5QVWqLhEggWTZ2k0DxPxpMZSYso3OVjqAbIF6HvbBiHmFiWdWJRAB+QU2+6FJ30
Ox7g+Vb4GlLetXSzqh3uE5MQNir8U1lD8hKUg8BaHDi3nZCP3wXho1r6KTfjshjEz1jPTWTKfCiM
IAMaQYb2aj4P9ZjYend0+tzGp2CGEOtIEEghO4GxTaVPPHg6omG2BEt/bF9YxaowOy40LnV8IlkM
q1zpWOy7ULvs4tMZLpkAu9I88OA1CVUIeDN5O4xeJYHoHg/eYnGnFeAQ9IC6B6svYutgslMYVk4Y
UnCIFKq7aT3m0e5xspns5xoTHAkl7tVNZf5hmFUqYG039dO3xpirGsBw4TVbm43EfDHidu1xe4dh
MOQzzH04cFJ5aRGHbiPGxPbTxm47BkXTU43FbCJMPMwFeSUwNZOwn1mMAglST5OlpHb/atgSHtPg
YjyjVBLddXPYsoSyzTYUq93bcQM3CL4cTbRA+f+dK6P0Drp1UD/Phv6Svt/VrQ/srVNSt1UUSpb5
n52DfhMLbYCR5c6t67RJm8AjsYR4oWDzvAXjUQnkL8nMja2VbcThCXWHNG7N19F4zoV/XfTDTK+7
1qLRiUvZKCM+B+YhIi4am09Tw44FLeSt35rzhChA2teV62gMP/Q8nQk7a+OV9EHJjWgSdr0koX98
9hGxF1Smlfem1r05/FMl8leDfatzjwIGueO355gvkfflWyPvBlav5AHQ7HvmrNBhmOIs7A4qufE/
nWLuQFs5dMzP5JxrHu0lcoEquaQYMdwHX6vVj7EqoKnSqkTy0Ga4XM2XBoHvEtj4mw4kx99KJkwK
mzIO935FzSI+e20HqeQvSzTtrct4MbODDO5Nlyb/dKz/cqHCngXFMYlg2uTYPMkk5LxR65kT+2Ho
3FLyxvT9SR1mKkl/YO9yLHn6wvGdfdyDjCCjp1Tky30KElQhQnRpk8dAkgeYvgno1+AqvF3HrA0O
VsjlhNZiorhx6gCHQJ9+IHZPj0dwWaB3gGV+XYqDIWVqMnHFW3VqdyCcK2BS5fKuy+Mr9KtRbLst
q4eCmiO5huq9gdbji46HcyuL4m29e4nUzMo/yzbQIG85Mk61xYfiXKdnOo8g87Nf3JSdl2txP5TW
EwzPlwF0kbOb7/PVTenVtOj175DAseqkxECqkBv4OEHvnL3C5QYU0KhZYof7ebuj6YzrPl3LVV31
dw8AKed54AxdEAKLWix0ym0ImlKh4pa+18kXeDzv56KlvHOfT+JVED8vr9UaaPSHtiw85oVQ7lAk
zOLLBInZN5XWcxB0CqvPJzzqY/IH965+fTtbMNLXZ1fyfrKLpq5ohfSUlf8WD75/CpgIkXvlQNCg
awhJcb7U8oXMFC4JGIPaV6rkm1DuuCd23End5KigzbMFys39wxM2zTxtMSoLFYnG+ZVNBO5/CYqU
N1JeRtjKTm80RbXdh/7WPNFJrE2Mid4iettTFwd8EpwPYIm3CoqiRAz2UitTPkyoQ1PpENJpEI+U
KCu5xnwCx2fqf/zJJU2kwZhr3hr1vydPjvXdHr9DwkNsfqCBkFlegiBkapCnni25o+HvzyUxNDMq
6ZFpz6b5co9dsbH2haOrvxMV8aKD+HtqZrgudq2+lqu7vzNilfNndFsEYQ6FBUNHDbQKsnF7u5B7
Pu/XhIutKxvx1aPoqVoiWPQ6Rc7n7IagB+tx1Kgpshf9W+DqsUwU0azlLRb/RPOPZJvdnp5DVWmG
80axbcI+t/6ACd5hVM/IESyQmISQqd29WN/mI1lvN/IVK7gbtfqJ5Ei+juVeR/PnSAeLs+Y1CaN7
KzgfsrlSnEwOU2f82kwEhxEIEJKLbpuKnT/V9cdfx8+bWRnGkxNrPePCL3F7D92VT9m+cS3MlffF
t5U9MArFcg+9kanm4/2bYLitDaGrf07bpB6+760lCGgJVTMWmlY6oBD27ixotmZxisPqyFZV+SQQ
uLrbJuT9IOLIpEGmTaDEaJH0EaqthnYJYsytxAOaKRdfBy+1hrKY4Dn5pdCYfKzp6OYtCnOi7QVJ
lbsea6meuu/BqvXjW+yVTRcidXcnR2oJQ5PtK2MdPVj//QDXww3xzN3+5ww5moMMLHfbWRSaR9MR
MD4kWdyHZO2jOWx9PUZrR886PnfJo2gCyR6+5IfwLJiItsPeoO19QIg0DXjffcWmEfR0oPNQGD2z
5pR5R0IMNBzRMd2PUWRSQiRs2Ih1MnplmNbTx1wxDPQyVHXCFKPI9j3Z5jD5QX7V57Mv+lMqTDwe
Q4vA+jwX+2oruoupOjaT3BZwLhxBAEQnCTr2FAoLQMhmsUnsebZiiBN1WwRYMqqgLI2Eq7au8m5D
fZL1CO0JtDRMCl394aQOLwFfyS7ou5jEyZvphjEwEyDvyeWNZ03+8JCo6bif+rqx5jACANw17RAg
fRO7T4uBYHxCNJl5hrqQRvZ6rwfgleTXf3KrVnjztdOGRIozM6OY2NP9+Mk/c1yFLt8xufxf2nLa
DDaNEuT1ObCq6OA5//UN6Da2lwu0Y5Y0m+2My/cPvHd6wcF6bnpNDD3MZLQMxCpl3pzAwl2/txZp
5MUR3ZKUrHiIHuwGTwXXWr1Vh4z3jVADjullLiURhC8WElPbJXHuByuumQGSY/t9knQgcZCrXrab
kG3GduHZH7gsIoUxVxVLHqjuRc4tQfVklbJ1s1tNPLDYN3VM/+7oENAwKvuP2Je1z18w8bhOsTpV
4ijPdGjFFzw0Apva0XUYJnEU1U7kTPyAHhVT2cfrfNRgvLUCam/yGBVW7h+VxHESScjfnRqn4AWG
AuEbib+WBgj+f9EI/joH8VAL0BozVj4ZnNYdR3sLbl4Sy8Gvr9kdEzI2AM5FdvCzCToykbQTYU3b
KLzJKJZQDDeAafUYy6iRN9zdb7zI1vwfSZxOeYiW8m0aaoTD5Jnpy3cKR+sFn8q7RSxg3jKrmsDN
T/69ZcWnW8nVjG2bQTrQL/Ipg6H63zFgq50NLJ9a8GkRSPmLXXBeiY19m6UjxP79LDODSj5OiLvw
oZDxNqu7ILm2rmyDmT5Vv11XC5W/DP5IyTaUs2QbAAii7E8AOPcUG54SnZiwE7PvESNnb2Wim4tB
IiA/qQcdOdO/CThO7XWLJr06M6RUSVGxgauqBJZZVYjTYJruN05FsmBxst/Ui9C6JfYaJeibGELj
Mr6Gev8vYf6Co3MDgxaCEJV2P5sKAdsGDa3xHBGVYfrzq8crh/0dtrfwA5G+PAhAqV5+Y6/df/hy
XKHL6ey4/cLxbkrWvLeKw2HVKjJr1BSp5cu+Qvhg8Wck/tWw5ixmcjZGY7xQCFRcplq9Z5v5DD/E
qoLlw5u9mvtdrF0QnMCLpkV/RZjAECQEzzhqk/TmV7BJ+qMCWcNLOwaOUzsmlfGMyWKTfDzwjGfw
BYSd70DjjqIs4bktsriKdTEUlhM7i+BBCJFmlXKxXkGfgml5CtzcUSFKZNJn7nm4zkCvcR3bcC2c
rC5ywT3bT52TA/dck8VHzxCgDdJS5xJ55ESNbKLXH0w37aN1v/VgMfvzs7fqNtCz7bF3F/Nu9eY9
XskNIl4C14Q7qLFvmbO7yNQ7i5CGYzlPHNWWMxwmAi7aoldueec01JGllozkY2OPy6topebnRCIt
b7jvf6tRVlgw/SOligoI5Cjj57TSnktNwZ+z3zkEv8APQHkbYgBOpbwwC43Au+V0oDMnIAUnLyOt
/PnjmG+2+cwslDFh/oFMYltTvdmVXoou1o1kSQkZaIHVGj6/ejq75IvPlX9JemX2fSfYUd2x5V7O
h7WT4hHrSTaVhrK1R7XmInOmp33JEnqlYxwol/NZo7KSayB4zEmD/MFT0D8RIsdbMjRnq7kvwMjr
5sJ4bjEawmyfQ67SFi5Io0J0PWnWEjDwHyHUKsqi/DvS0YtkYp6/fFmKIvIW05BaMwM7TBvJHS1H
TESm0OVgol4NlLT+6wBKAyCf0tM892fGAHVtOyhIARmQgyMF7vjHNK9nyFi7kB96nNAn4PbUIKFs
DuXrW5PY/Tda3/Hyn96a9/MHdjhYMwet7Ky3zkfSxbMT684grV+IzPr9cBb/Tie5xWU/mGtArxzY
bLcgUbfgwU6uEmSzQ4RZZhowzx1E3UZsHvgYEljRGg7WfUE0ZLV7e79m8wSrWzVgk80QcquKlohZ
r+T0gzOYNJ9V7lFmIs0lXX+Gsy/c78b2MG0bVdZEnHhjJOdf2iHT+kGWgaEeUaXzrl8C+bHZq/iV
YiWgwP71mTLyB92RgwFsQYfqTS/YgUKV4PA1cYecGEr/+zWhP3/AVcr2aJk3J6WkVaIfcBT1n8uv
uxGY7S3pcXOpEbJSA0cXKQbxivaVNvgOP4/YvpJS/QELfDyRA/8NPwQYRkDaMOFuMiRhhL2CTHve
1zlqcSJwb8tLOVoiJ5WWZQ0jqnY9eaUqHrThq4YGjHk7mZ9Ft5b/K0Ql0zP/ZMZuxqk3X/B7Apr8
cCD4QDcf3jnad3RG0g5wsza3hsZWRJ34E4uBvRFb6F9QTfR5H0HudZpWH08EW5OBhkHclW0o2+nv
YUamCkThkis6S9/c1CYdlN4bph8otcsr6DnwjMNFpnTyB9PCjdfoFEdSBpeY2nJN4GHJdh8oMHr8
U/Auivb/YqlInskKsnhF4aI9dYeUd3KQ22XXFXsuJiTHwfY0C+sWPbpPr4Y+abriE+w8TCOBhZGM
FkVzLCrH5+kiQhePEdB0aIpDuqxYjeePwBBwtLXYBRzPkilzJkTwoQz0fJVw3e/6p7D+3gx0489U
fhJwwMusFBtZhT6ib9u7a3OHNHSC8uGKWRt+47hu10GggUGQ77uC/aX4JerYsBH5vUayqNR7J9R8
AtW3woVttDsKs4KHowmt4OSDcHXxfakqNRkDitNGB1Pxut2GM6Zr4p9nRukL2VEFvtbKb43wBjBh
lonlwZ2eeFFmdXvHz/xYyn2vpjJctgnNLEMHodgdhv7/4Lvq0MzvA0MHAmNjB41dXatKmyBTxKDK
y9NdVcYCdBAX/oJh32u/UT77PKzjDyYkAr7OjTko9Ps3qxunTIZ8G6kVzWBX/oWuSFSYjNIFQWWG
4ncX4v6/XKHKIhxUeWXeLfvM1ksg9pN5+uqX57eqhgGaJw4wKPX5Gi6sIdUuCzia3fAzL8meIMhI
/kIfZhT3t1RoZAMy8uCtO+0t2VvROiHoCxOkUzb8I4K4XdvqIj04mw9mSHeEE/3fHiVkwG9yKhPT
U8otsYieApwEhkbBg7/j1xxux4Ydc6e+4v8x0ZbqstsTyLzW2p7Z23J+/r1rrop0AOetMXgXbMjW
+u1gtvHe9x/xt8FI6tKczQR8yRMfXwlb4mxUdkpGtCkx5oGcMz89AoUesdD9lYiDA95nP3EPMDz8
IS5n7nhIrKvSEl4/cxvDNQXiuTp8fncT4A1gNYyaxXZPGCpu0kdk+VlankEff/DMwyjeWEeQrARR
8u3U9pppXYGWgANBCVflCr24RvqjTNmeEw8WuJEG9qMJf99MemxQaSNwbdZ3FMgypsHbPWIJc9vD
mEphQ17bSzNJiY9JV9JHPN9IKWBLR7I0P1paxyQVg6xE8u7LMfg3Q7x5u2ir6NQ5TVUZmn+GW+e0
jLEA62+Vs/Aj2moy72WomtU5QvY4NxJkXzSIMrluHBeRJhkyW29NadiJX6H3Q7nQiSAKxV1Wt83p
yZsGRdPGb9IOjeUViKvTprbpEyGy1VwyRaoh73WkA45sQjYqUBCZpG4YqpGGpbUuKW7ORdj9xArY
r+tVuIAqAEC9++xZ7fT0x3vTXCtHUUe0eB5Dz9rbck62jUnURMfUpIuX+WVAGw4DdV2u7RDn9TUf
u546tkVQ5yDVp1rj44vVvmrRmwYEPlZPGKI96rlhtMNjCLA5JayTu/F0dYf4Xz2L2wv2t+KLGk9c
wFljS5q98N5gv3e06CmgzaoX8Z9o6wl8DiNTup6ql4S/sx+/dbOtYhAulSOhTTkadrzSU+jaCpiJ
I5kVyfEw3fmXqGbIfBZDdl7NrXk5ZE5vsjnrfVYKvzuLyZhyRn0ZuKgOlwPED2i9kTjtzhrOqFvX
0XcvqXLP2Ah6fxqlG+0eKkF2rAGbbwi5R0dOf4t+SlCMOLsc0IhkhByYqADonrpt29wqYVE6B3y7
D2G7UnH30qLGkyhJ6r2/fziT910pa6dVDJ4cUAhWae6Cs8/P3oTsl2e5pS4AJdd2ItA7dKkLCVkE
lVQKgRLVsffo4tg7KUAtv+Mg9+/Jsw8tj9LlJcnDkxCndA1OpGqsLbMS5XkXp9Dqi0ppKKNHycZJ
g6euyi+tQenR+8ymxc9pnk2KLcrktJxKT0NIugrcWbNvjwhnMmZJIDCxavzQ0ucpp3R0qzStVu7c
4nHgbH57ftSmiTC+Sm3yPQ3u509GA435b6gFf5Bk7tdIehfy41murnxeAMRzgVwQEE1K/wBUP6tt
RCGPmmmY7qPNS/XhONAz0oOE1+3D38ZRL/8FmT6qIILVEaFgUxGuS4g0jOTGgWaZ1jFNuiPLcZxU
PfbZLzWCJQ+B/G8VzPB6Neqab4DNJXQqSdmUYDp8CYTG7E1MRaTI3bMUefU/K0k/WG1g3kUI5o8F
CDg5aDAOpkadVbaAMRD5YHlKoFI7MrXdirXJyJmWVMTo1QI0CO0k8NsK4MIoVEcNWjmwKGu3pF0x
TdhEF5+VUV3xekbVeLpEW6M9ZcurKJCd4Ph/emnNkz8o46YdgCIWXJdHn1bjEoNjX/1QmxX3ihUE
ZDv0nG84hfb91sttQngGppqOMDDEcb4uyMXuZh+zn13cdiDe0sVCP3HMgSRtafz8A3xja/2cKYqY
KP+J18V7uVM4vEktrcBn4TpPj/SSGVN03Ay3rCcFjI+BNDHt0FWqKDa0LjHtnZ+iYgzFsM9rQ98T
gmcNO3XzcfJTQKNAc6Y1nxpHWuzUpzj7WhpULvPrHz35k7Jrd3dcquihlhBfrL/C3qfdbRTjm8ZS
fFHFrYUgJ4lOFPsBcFkiUhKdZlAaakQWFQFE9Oas/AI42q8iT382s4/mcjtdhZvEUcCL2/TEiHVV
NAmURwx9qQ7JMt+RYCpZEIqtG34mHexWSlglRAlfpTbDWhpxIlZnANP4kUR7vOfxsnk/FtHnspCh
EaUQyCqER84iB7zi0bEPaZVJdWi0CU85Qlsoli9JmAnyCZyGI4I15qnKzrAd5MMRoErS8MVNCV7J
UOQJwDg3xv1sN5I3RnmI/5kAO5K0ThSBPpicB8YF2BT8ewybkyCouyjsFu0dEbFoDMSaYwuhOpdE
4fJX9rGkTeHnT8MUIWnNI5+dgmCKdtCKgJCKTohfA0pjnFma4RFYBmdgbUz/CiGvObVZUZDw8YOA
Qa3vT2nQ9qKMIaE0LD9wTCeC2iPsQAQwRlXVkvKz1VKpZIhAwXCnYiwr5MvxHSJND6iRvsG0lsB8
1zjOiAx4cjmBUukaCaAc6FMTX8lq7xtPMhjEXv7yA2Hmy+GYutN5suynQQjqQFRFwbvBbQIKh93P
xZimfTbUcH521ny+KqdUPyDbXJKhOqLPN1VWarj+q1nzf+p84T2dghtvDvx7vvm58vYU7GTCcYiJ
v/haYdIjEboMR8VH9UgGWDQ9NPuVWZ0OKrWG1xETaKQz7Ii9smh+kG3xaUID/8p7Wc4FkfgP8JQ2
xCJLi8sd3FG7hqykrjWHdwnQxumpIsc08OvMyT2RHmlZ4agBEdqV7TlEFoqFAulU6HiSuyM9V573
fxBpYQ7xRgWv6oDqldpTheKN2qdgl5QRp2stn5xoxzt7e4RuV0dKEs6/8XX5bGs9B2P8DE12mpwW
SP0+bHIIcsvhzdN9uFtffRsqmoQz14FHe64iw0wGhdxAe5DQOrsSGO2wpPqsFy7185WZtaxd007A
E36jmLO+ctgWni4noizF/O8yT2TM0FVS4MDb/lGU8kr+Zq/4u2IKonAVo7s2aF10OtM1drqrtnIR
qlDa1ONq/AvoQB05/c2YfT+MZCcVb6oHIa9v4zcFDx7CR0YCMTs8tZ3J59Ad5q2eWMH99EuK4R5s
4QySqjEVvQaW/b9RecDouqIMzwfSNZh6fflhqrrYO53M8+3+gj9NmQfhdf6i6ZuXPjt35cI9dpyH
m0unz/5N4An8RoHlIETgv3TBxdzzTKH9i8Uqf0KkiEITXwiXD/Q9ixDq3RzZ92tepeVyMVmeSMiD
gKNzGpNYlbsKniJ3LDeJVoLvzAy75WltkibqjdBgo5sZV5sl6hHzuj4kT/DnZbXE4oTXcULBxrcA
pwQucby6EUt+eTXarURce9/O00UAZI8BUibBudtiN9Uf0ZGdRsWsYEx9XW80aJRz1jdKYztLpjr7
V+VUpZnZBfy2GKHyUjtL+Upb7HL1++JB2cTIIfZKgk8xj7l89fLDwrBOnQ4WRmkIu9PXyNpmOvut
jtRBcX1TE8f/Lhlr+cYyzv6ihf+YOzRw4D4Yynn0R+nR8fsBZeeeC/Ih9zcD7Iw0J0PWTfZ2uhlL
gU+QPvJ3CQ/Lo2fiCCKKsLOpehtCcT9mWF+ad91vS1tn/gSbFUhOdsX8Q2/OY3T5ud6yIBW4sDW/
L8I1EUPK6N/bv2+MH10Rw6MWx9V8HC//bLSe1oOfDb4ewj7hTJ28AB0XTw8OxaSd+nv/xa5/FcaG
U4pYepWLrLhMJvaiF4muRlfsgD8mLpXv2foNKiln+NRgyp2C4WuO7vk0iNvyFN9JnkWGmObWqLGK
Go1RtbaIpRaSOWm4IQCQaN6BN5porWR9IUGqHTPb/+9wdtUwMn045GRqV9e2hv/J46zlYzVstbtK
5tsCr1RMiuxl7I65qd1sERmsEFRQAKiM/62qPCqjPXA+7j6dJgK1okkoXtF2l/mFSFKfup6yNza1
nEhqasSxMR5yjw8rMZPYRqC4sbsaNSmLnKMWOH8MOPWaHApo0NJnT4iBmKF7DM9TgLEJ7nTCmTmJ
lRhjhBWSlhgZTgwkQE+fVSpWj4npg++AZeipNLICtasTf3nTocYnJaM20p1UDqKVy5RxG4SDIxeu
6ATyLlzBlp0WjpEwLNQ3LP+oXC3WiBxfzSy/LSC00VXj2wsVUAXcVWnP7ET8z7qV7FJH10ZtEsbe
eP8QpiafjXgZ8gurlLsb/5agtRnuOVFiULCW+ufTgm1VVcgVtVaMASvQLLZJJIUeFEAseDPVwEgi
vPMp+hgYQVbI1aEdVWGXjVhfLnp1VkqMz1NT4BpWk+gn/SHmHN64e6Ibqz3taYkJGEfYm9VgXfmc
G23T5gR1th7ADyRliSslft+MnaUf5UKqvJHz6MVXgHzxqKZ/+1FTGOupdJHQi5gWsGsT1wzOimLn
TaTIA/VNe7DN+eRYNSAQCk8cGz+Xzw5hOeb8wliWWvuqid5pF30SBN/WUCj3GkqnkM2osdPWIFef
4Q9M8YEJgh3LDHIJ/uz/j3Jk6ZG/ee0Tap7X+TUrjh7MFrC4lIg0DR9jhgOXRwjYRC0g4r6Y3mvO
fV+j1gNb9QhdL/EEkllAm0jWAGSRYNPU3Bsr2r71s6RaBcfKru79X984M7utKOFy4htLuqVzrk6t
fx6MluMGpCKgHmrI5fXXLTWmeNts57678oKi46TQHmnLRnnFxDSLgec7J8jGxJE9MkAtyxM1BS78
AIu5KCom+ISJJKn3FS2GOXgKtToO2FTPCRO3XS561L1w55ReO21xoSzWmogqzWK2WT+3aRaevmwe
FYQoy8gPlIcMs0X6MJsyYIU0xgc/ZWmu9es8J5PWqC9L4ZQdLj2/dRRcJLz2TXnCPsUWvsh9u5Lx
VN8Q4Gir+CDitXHhyahkiNUPrcVS0FfVA3kYvWEzZqxSoL49curRyhiw4Gq+20jXNk+FZNGzVm+H
qwIcNNz3C8UTPrLPS58ROVGq6kQzoTEPTOsYcMBV5v6fveAQeDvwk8EyI6hs/TbEtZ8Bn7let38x
+3jDj63+MRGupp3aCmg1CN36wmV6BkjoBNfm7uTt33p8vVTptyxGmcoUTcNeFTUgto1f6gQzioI1
m9iuWkBEYd8t/QnqJ8OT6qbedJHzwBOFunf1UPKCDQIvaCaA/61weFvuaZ9aLZHJ/XjX4nf2SYwb
IFWuLm87WVBZ+P4CT/8rr8aGLy8fMBe8XnSMczU/dw7KdwCKRkV46xylfaVszzwf/asckyI0c6Lf
Tdpf0wyzL3fHFhB0ZLV9dUQJiVv52liswLMyX0EOKzVemNjVTIRuetI4bEjCNPqC7AGCgpxlzrYs
IkqbePX7WyEpXnukVdd7x/aLszm304Ba+vVgKFbmBXuYAbSpnCrt6q/uSPm36WMMzHThjBmwV7iw
MIn+246VKL1KagEmqxskvSWvqJPZLPkPHBJ99eNsjYhHDtn/URrLdp7jCUTdQWnyJUkzRW5Dd6Xb
IPKafHh8tT9IE0/1XVzgo4WfTEFL7f69yjcnT2NmgrmLM2V9xxm/C5NfY3YDDuRKlqPlTVsq5bY0
XzS+rDTx6B/Fl3sO5gln/9zMsD/KbgtmGRBLA+E9tQVXjzgMzOGwFB4oeA42BwaNAqSAPNycQirt
QP5BCigge0aaWlwFspfY0VODmfsGj9PAdeMZVgGqSBP3+WC4Rk+gtcjeEkwFWw2Ux/0GIbIJim8x
Hd4JViQ/1jqYMIan3gXx/UqYU+EWuCpt+dqQb154nUPjMXfqi1glvlZa7tb255U4DlyWZWY9ZMUP
ljkoKKwqgyni0HDdAgRRHvnIAXwEu4M3FXfK7DuICFvb1q24ihLwT6IQghnKG5ZJnGfxSx0wUDMf
Pw3s5X3FPwT8q8VmubGSTceZCAwE4lcM9Ldwr9G34TVGGzm/wupoIWEto08yx4U6ineCYBxeYWWY
PUpvAD3+vkZtLejCmfs29JrnKqdQ/3o1TB/ctnGGAL3jSk56rn6Tf4HTrKgtWSJrcpSfJWsFeVwy
FA0vxeC9R3W16Xo6NxVZz8g5CdJc2fQx1KW9YB+RKzM5EGUlbYNE3Yl3jPewSHOREeSG3pnMrtld
jtPoAlycV635Oo2zuQnJgbaVra0DnV/MKWccL8icA8naSWVTRvo6wZykdxHXdCxginWgmDSo6OxN
J5xwa7Pbsqhz4D501GGZJA08S9IvSXqF/z0Ccz+zglHkc4lVnmLailRViCA29QsUr7zwpy57CnVk
VVfQ/rm5QvOhqtPSHL91lp0OFfidq9LnwnsCvPURO837ttm2cJlNzl6a4mQfgw71IcwX51e2TQof
jpfm4gUR9+PQGE4CPJTns6v8Aad5S7GSpCOX1A85M3wQNdiGJEdmnjYfrjh5FTDcZ0eJe6CSp1LF
ZECs8ZLgEtqao3k+pFFimF6ZDNJnRWOrgRe0yrFWaBTsjUkuNsa9uVa4ZI5/G2568mgMmHjco58g
sIhJUsTEBTHibVa8ncG8/VgZ1H5T5OhCwVi4LaIP5mSQgkNzxFHn7MASXM0no6mc5Vu2nrSPnnma
ccPUqVSyCereokF7k9BpRVzu15ELIC7Vclfd+kBf1gR8ZzY/5mBzc1v5me0R+aRKpoR+/sB2vTnv
9qQX3vOjA4s6RcSItWB6VY0kMy8neoK99Kv/sASF9R7+Kh9Y8fgq1KH4/PjFLayfCCdOPj/UQdqc
AR0/zeRQtQPtLK2PD8/dnqJ+BIk4n0Bhc/kXjr1xSorqGODr8IJIRCpu4eTl+AsyYOcAaTftdL/2
vmJElGsP+eGE4CGv0iYycIfYb0a4dpitri/lzxX6RIJJknwHiKZfezOQd/1vu7rzaw3m4ZCN+Q0F
ryrz4uGZtQbjnW1orytMU0zIkI1w0QwcvAJ6DakA0hLIRcSbxI6xfFpE3RpfPw5vOsgzEfbAnfb3
JUdyKMqwNgUtlKQujaAa01wpSR+j3ztc/F4ZJI71BtqnYMyKF136STx5ncCCz8AK4Z1vWRFNe1Pd
slT3b8bMThcYxu5HcybjE3AMbZFHKm0tWIMM35XVrunVPI7OP5Ux3fszT3K3e4l9VOFzDfNufvyE
w7Y5rttQra4xpw3P/LTN1do4fCTgLnxtazlqC3Ifo0neSYjfsBnLteJY/HPcbEYwSOFOxwT26bEv
DUiu5hWBcJaWfKqA0cmg1YG7PRw9U8TAFSmGrSpmU5rqvILsB9Xs1QWHWL8wNS1VyrX7HIgRHiUh
eVMfquHjZuMWTtVPhAVRZI6io7+uyThZuGPO+JqYCoYaskp8FX5SG5tGRlWJvBKf3BahQlRVgTLk
fbEmYKrkZPd6tSFI+aWo71gi6B+qRytmDGs9/i/2SCEB32z+A3grUXNOfhRgIvd06B3kGwdzEtFc
h80Kat87tVHSD44eoDSUgu5NiKapq+ZDxa1LCeT9obNCD1c774ZrZu1c9gpLNawGoQutdmGp087o
tXsMSJEQV3L+4nmIH8643g2r/nvk55BlMtW03FbQh+N0bKzEnkK71PmxZu8FHp9Q2SnR5qB7FAU1
8Q3yFxT2/9K1aFyyqe61jOMA9GK8E7n1/vScVZUIfofD+7vyA+ynGZRVjNVok+2/J/d1175wcPMK
HVEP2V9Gfu3LbhBieCA8Rn24XR14FiJggAl7ihNLR/l9bIo0FfV1u1RoYwKQ5x4dJFHX/uYU75BX
doMMkjebLTz+Tje0VOcTxRvZACMirN0HZF+Q5NWdGJ3m7GtlPi03SGsWe5sitC7OqIxouWmZc5f1
LgNSdp4Omen4DiSa6A/8QYqzybsD8PL9rvq/L4Zm28KqeX7vA5iDHifuJM2QU2HP3Kg+FKxM6Y2K
ocrVBbIfsUW/kmnYCsB6m6DS8MnUUG4EYoJg0oVvc1ejyb55a2dlDB/ev9KERFtqcKYm1si0K03C
rRAEQYU0izkNeaitSdp86ioVR1/zENBiTt/wE0G3XLo+m+gpR+GJycrvdlw9h/Da3FVLv+Dxavix
N5rwz8Y96vHjaCsCnpKn4cxrdQ+BjNEy+YVpGgQkqtKIaRnTZ95NBh0bFT8UtGpbbVFKOJ3TPniQ
EX1QoP94PsyFTzkcn3QE3tARZ5iC6LzEOFekpzyz40Byr2a/U2jHiXlHn6bnZzLj1z4HpmtWZt4n
TrADInBhEM0zTm8ooQOHE0iDsBU8vQ7Cg+1cVNIZMvyT9bQIm6sau/xFLrspvXP1pMO+3VOqIGTH
T3XTVt5HzTZ9Nj13d+iSYNacFmhvgS9Q7U65YsmpS2cd0GIiVHqhIGAH7AgBlMU5swzfFuHhvxEv
CTmsX1BPIygf/RHTN2DaUPNHxHjGhx/z2z4HBSqCK2Td3YrsOY56/ZXsWJsBDunzvTkEdiT44lV4
8Ic2cZ/g5zrlFIkk+eU/D2cd1wwMN/UEhkljTiRbc2jORkwLk43rvob6ZaWG1clnQZOQhJApM168
2NTsXXRcnmFAo10Ha4V6p0p0gEFEeIRiwrusSngpmgBYuuwldWOhMpd1rJ9bPohfm6dtm2L65HbR
EBCmNioXe8OyQq1h+1XKVkezq9+iuAgmeJpJb/0aE7Gww3ImQaoi7p28AMarCLkUuve6IO+W5uj1
LNowDNsfPJKUNC54yaoChboaN0i2RsGtZKW+i+fODElQ+fXeGEH3zFNM9y8lLrct+BEAw6uEC6QZ
4Fht5RqGi95/KxupP8qMkpBaI9ASx5ywFDjaHjv8pz0SfSA8+tEhTVgaDmVNdADtdzLrfhZ0Gly9
EjtVv6E4CjTmS4rHKZ5H/4Jgsm7ZuDANUmtaMd22WlCuXJwavDde/U8Evbo8ORhenxgNkOG/UKHy
EMcN0r+ny6KL/4K8xBrnwlf1EeT10FaqIw6b5NSoI9a8DwqLmXjbhqnQoeutsjkQULeI6fkm+VWp
o2A8lQzp/aoLVmvpUkIFlYeZt17sin40XLeRIa7umT2L99Y6DmgrW5DA/Ehp8uqE87tHZDQnoZCq
pDI0MNP0tVFIs0siKOX7UWSh2KIY/LuBmBVFRIfF5lu7CkMLJ0yZ+GcvUd/n8FbG58lpbwB4vWZD
eQ/qtfGMsIC2GcR8kVGgasplF6pFU7A0lN0pmhKA9cElMXeITDjnrtnnDLjT9MubYU1r0sbEu9oO
ocRt6fk/VHOwkqrS6FSt9Gah8ku5tjpGDAgNFjc1RosNTMHiROTG9xx/XfZ5U1OslAAFWsHAR5bo
+R1e4+JTRuUl6ZMNgj9xylHTc41ZTMAUvjsDLO4agphJlcD1ZAtp9iLYFRUxw6RNEj73WHXGzBf9
s2wY93/lLnQ290XRotoc8m0/6c3r/pphlPzOQttIbLxILz0ARxa7e5D4FGHnT9niboQo+xpoEV5B
ioHBoxhVZmtX7BPUeba3FZ2dXQSFd2v3jMkHcXT8yc2nKsI9C0ofaVNvNPpxOtHl1cZoIsTlc0lv
7wBQ3EUjmDNaXg/t12+cO4ED9Ww9xBiv0CFuCYKxgLdx0keWgPTlJ+UfGrC6H+2r6lVJyakHP1S0
PpWpXkM25jtNgwj9Y4fCb6S6bhdwDjXhgBYmpuwsmaTGdWU3xeb3KZ2SFx6slhFlfdTXi7Rg642G
RNDiOeRM8eMfGbKdOv3GNI3LzSN+xZXJoE1uWOGFCyWKw/QCcDvL/KlOfbVqFNUk8FwtmfNifDC/
NV+gRnWaru1MVwMDaY2Ei/7fD1V6QOtBghhy3+bCQjLhFUK24kctaZSEY+9rSnaIV+LMvRIx4POd
EifVicILPEacO+Xinhox00hiDJV9bjw2POLEumJISdXt7XC8msI/Iezl3P1oStMrFX9kHUnsLJ89
v9FsKSerXLTUSbz5Ifm9S5R370dhBNE2Ddgy/uoj9lSCSokjMD4ORPMBcuF3/STjqA82CY/5kd2X
kHs8LQF9/geyLNN1XgMbDXAGl2o4pY0y3LnITyfR35S0oVMWTr5WE8Ucuw0xaxtytHgLOZJsmYhp
yJ34i1siy0kXRQGTiT+G8b91VEuH9D/6GhpGHDsm6Id8fUSdgKvuWTfCZrT6951QXjyIP891RJRR
zLxf0N1DLY7pKPSynanKv/YHvndY7OUxjtAhRcJuLZQVIunCXkMMBLRQqzLqsMk2OJ/QE8ug07Au
WTRJKJDS2xpwABpeeEpzssfLF/VuM820ZrBVz72bN9nGZenTO6FvCD3RBYwMJkohD/i8OmKkgrq8
+vbpif4UK7FjXlBIKhQKA+5pth0LJeRoE0SYEl/gbvpwuwJt3PNnP560u/sdCrdM/tJvPT7gcBDe
+KVCev+tVw4QAAn/cVj9K841o2xqU0E5WotGc/rWmIFZfJZzFQPMUDzgwbyIuMTx4lirLC8Lp+v/
dwh8Nw+jqNJVjfxGWkGLcvOFcz45USsRZpK8YWxJxbpRdzfF8exyeMCksGf0loVGaADLWd1vCC32
1e50zVClVITVJM/on1ZE0RrYOuzZKva/pqerUkaOGQ1U/Fs4mZgOwKt+BMxYyPinQcvxEkxECkt0
lkOnY2ucWIGcusDGfoTr+MBmdmqIbtZTNvu84+NGJcNukZfdiQbPYln/JG/5N2vQF6FTr9fOIntD
64JRZBwduSY7zN2zA60yvOkOWTWcKjE+i+IFq+q1Psuxfecg4i9M1EddN8ODz+BRQR25XEci9Rxf
Yes75T4PA+GpttKgHWvb6xue228jR/MTuDo9+4Ubshwe3ou15fEmF9T7BV66NpE6p4himJEdIeFw
G4sglEJXi1s1N/+TiKu/KdzczG0uoxpnnQrKAH0qr8FR6M9mC151Om0e6L4uO5+hpWBKd8CK3Mmn
zFZIsiUyiiknSjO9uHeIfBPEXvxgmqttFbypEiUZJdZ+Q6nRpnApq6Gy+lFg/hZuzyECWL3VjaLt
P1TbaulqbTeyk/M+U6KlXvjSuCDbXOC1uH4ADVO/jc4QpruwTDVVWQD9YsFexW3AC9TjwnxIPzGY
SHUhlCVQ9wZljWl6EBNfBzdCpJ1/ZkXe6PEu+wb1+ZyC9ZQ2n55EP9MO74+79uPeeVTmEdiP0lZJ
urkq24lOGukkcJXoNe3OmHq7JQziTBZyFoaXiUch0rcuYGFJriMv/INzumuGmS8qRt8jXdrtJC+A
AmuGs4HLzC+9L5odZQBgaQ81+rH+b1V36wxKHC34pqq/Niv5pzBZPyCOfWN9RZmsux/SaS/gKIj9
uYUc/n9Jw7RcGmDNrOY3M8RUyWTnDShBQbRen/2sC/rs9he+S/hhkRyely/UMaLwJhxSIU4pOrL6
RbIX42F91Ez+uX4dv0Pp95UpvnSLp4p9YfCIyOeqOLrZAjoLXaRpatZ6Aem1DnFCBv3TnK545GFK
2GlXRCgvOiJzZQF4Rn9vTBzjRsoOKGIrKxzVm1pz/fz2mUz6VG40IWGF9uawAU9pjZ0x8ue4TMhM
NzURW4RCqyuv8v+gFBMLAXCCuuEFpvHaGg7bQnH6yMlrTmVRqcbjsCxCXrdgI4yRx6Dh3bzJorRY
JwqQqWJ0jTcF8jUxKlCjhgvH2WzU/Gw65+7OpgSA6s6laRpNGOWnzzrEeLfmLK6kTPDM7hZk1l8B
s19fDrAlE/CLZ+SZWYutQqMxTalU2KouJUU0YtLTMyKYqWEp5enxGi88Tdk5h9aUpNIAwEI36DQP
jO2M+6OynE1r6rGYFasA/kup4wH7WIEs2fgHyJ/yw+DoUuETTrWky0U/qwzDEab1RVLu1VbbtH7S
hqElNzihkRbRnbGRryM6MbWl86maKhVz9qJTkLghEOgT4+1sbKa47quf8Xw3nu56YaOZoBpHQkGE
PFFILEQiLZmNnbIQjoBwme3DYqu3FhmAL2kpUrvIov371qybNrpm6hYy/d/uL8HNbbzNaZR6Kzo1
s3ZtDJVZIj9g+7h2Wy07wEB5SAkqOUV0slDWAbORQJiLPKsnUEJGfmmJNu1UCnXze9rkxzmB5EQA
8fobRykOtdj5n9DI/JbdRUE47lLlOizlIXEdJKIdWSJEmY0uNa6nlUO7NHO27WlhznG8k1QDg0/A
daX9hdzE89V+SpMlhf2pMill1615D97Qf+BzksBqkv1VuVK4/6LVJ/ecM6nsiLFvvIzkQGbjduHp
qY6J4cxgq9JxklPwhPi75P9WJABFT15IWLHWNYAgiKIu4EaXIywmd4TM8xdGKtZT+JxA1Cl6ykta
bc9IWqpt0IXGeLDXVFfSsGMUNC9h7AaSX4I9qRpUJzrY+rzFvjd9x72gba4WPzHvMqMsaxspYmBw
BTMxzjl2hV1DikdPvq3pVDS9kfDERoqsdVYDRDdcPRN6Nw3MUcHDEb9CTzF5VGw+KNBcyFZYibbF
pNTgvJsNTiGBy6D05ndUm8rLrN4xbSIhRYj+RX8tYZeAS4slxK9dC/vPJ2ywqtCnWFT7BhvFzgbZ
E+FmuZ8J+572UsbaAP7d+LO5gGXXU0kFc9y2wYIrD88RRxdqN2+xjCMCFbW+5bZUj6z10ECiwiYm
grTRtut4xegpAGyOt0jEMXF/OYPwj5U79aaCnrUdaKE8hHE+ei6o1aUiA1DlPlCmxSycnv4oORw9
aRoxGwHZNWcRhnTcjhMICyhT2zQ6QCXHnd07ZDIDXsNn8Xy/hzewLxCOTH0LjeOh2cZ1SSRrEVhR
pBfthjpDA+iut1WI4bsTBg3xfiGNdmXrHHvBMbItRr4LgEE9YtInNRQNK78JJQ6209GlBg7jyZor
jFx9ABJn9MgXw9DTQ34tGt/R0s+wWzv6v2jbS7FU51xL1HdLiWvBrJp6nOUCVaS/4JPf/UPxH+mL
hnElLW0Jk6ung0IqEcJPAXtm54wjOMC29Ff+0fwSBfNe44n+ikQAapWKyZ2DYJywIdFY9WfPJaQb
/Zj3X2ZFSik5M3x7n/EIuefR6HR1TAWIVEh9TYN5E8wd0OKv40dnRrNxSKiAnGrAf2XOUgzODjot
pqODU7dhvXVEGoZzITVT+FHKFc2P1mEm9ZU5ClrAJ3SSzS5NGdr5NyyJK+CpV/rMt26W2NlgpT6G
1VXCPE6ZIruokhl1ewZ0SThz9tt2rhhJR5eCbozmGKb0NkI9tn62Tu5jc33a8IuyDSIJCA/37p1j
SVDOe8q4KyjGcIN6E/YDV0VgmM+0et/1YZU8lmCqovowMu9g1UMi0mFYqCFM6glpNqLajecRmTxA
eJo/zvjIU4AVCCakFoqcVg8Wq3U2yJoYe0AhoPU/QK4dY8MA6EGIwkPtl4SlPLWtRETmYvFJDZuF
U1ZN7hOVT3Mc/E/pJDhOBizkI+fAaGK8aGcnNltUOQBhil8nf/vV4siS1YYj/UKF9bImDkfpkewa
AVQuzQR4ftYFxODEPYup7v0cx+mOYGR55cJ+YNc1sScQwO1qaY+99J3HfKIR9frHxKvHeemUvsnI
UzPvIubjBfL8aZAnQOmLCjUkmh2F3mb5fX+QLrnAE2n/i4hZ3BlgFS26FKCa/8W+pkHWK7Vln9jE
eCyUIA/17Tzvk26xmNjn5IFIGi0F3GT1HkR4j41Dy2FM1eFHJMa5BwGpVkPiHyhnoN5N3f7QD0+L
wcVNy+OajskyDGsjpwRoZmgTHGsvC0szOiCqAqktybeZzxcJu/uNjN2mVADYlIDdv5nmtFbfJgbj
z97gX7p6fkclrGktREpuhrz/15nqXoqren7ghDjsHNpNJ7teNqjUEtkgPek6qeRUgaLp/j2foJes
dbDROF6p+m5E/CKwCdhX3KeuyfUViUTCbqowujwhlZXn30HI/p9xVWZK97s+geldZZgARjc4KvhX
Zts0RFLo0m3egaFXmj9q9zZAPnBKvlDfPeypodKz7YlJ9VG2WgLml11V7eWjaBDu/+/oivgyeyYm
0qV1Vz0IcccCrfTSQ4PWqZix+Jutkti7YDrZU8Qj86+8hQ1c7cYGJOjO/cdgbEAEWYNJ9iLa5PjD
aX0OKOnVy1/1KbVmZNeQoqrMPkznribXT5np8gQsdr4KEmqaKchZ80bAqbSW96dqt4lzYaymTwiB
QSFElMtwjE9QW5Q7Wvv0I0Tv/u4Sadw8/0nf2bXz3CgBd58G8KKYXln2zM8Z6MPhd+H1OM9l1giC
foebN3/mG7crd+pTfP4rajDVQWOvE//U8UZo9O17ySpCDbC1MtSSPkDm/5bs1HJIN+j3so5AhLDs
cIZ/RNivmgH+NreUAtE9992bws+qFjJMti4FbN4Bjx+XM4VznJG81u+GWztgfVC7v/GWUdmugW5a
JS2yON79+jsfLpBXqDh/rT/bBR5NEPN5zT6zS0t50DkT+b+mJFSKBOcJRHbO+IyY2eUaq0nYlvLb
HRsi9X6YJBuUStan+oTU4ziZ6sqUVzuisoUyP0DRXf+onIos6+T9wqr7mNZ+OL99fQY3VCvkw/l8
raxcumfaUygd4NyQ9a2EvIKrTj8aGGv0r99T061nSI16A9LVldSRlkA3ZpCJ1+8qK81JqWjkDL9f
3HS7dIipxiHpV5C7LNn/l+7xWoFPk1F30mY2ynbZYzkBTmhODeQKaprsTxJTYq+j/xcYUfD9P+DD
3FA6QxNlt5ibOQuhZhhbA24fzkO+539nciO+jCo94VlOAxJyySCuiE4051gkij3V9/gESSlKY5WD
p6i432GsojWk66WvynHB3ryGiQB1cDhOi99Cz/tzb/UOA6y6J5d0q/cJGewIqLOiAkfBqCBjcSCt
JrQthA9fKpIm8v537RQ8/Rbj9zSDgJX67eRcZ0GqCi6+kvoMOa9usbzWUOUOapSsqJKvpuB5WtCo
xhMMY4iULbxYUrUMBWfI9Ma9U60e8DC3S618jI+hhUiLWtONzDSDrOliO1O7rgs4EE7U4Q/USsw1
+u9ArVDZE6wnB47J6u9KtWMfRA498weHIamAP4t6rZTFVTe0wALMiodNCzFceOMhCUaLLUCrOgDr
/w7JCHWHv14CbP/ofjILlAX/oY9pTUsWw0nd3nK9+R3Y9kSfn0QV1MweMRS203PLy9n1UIzEx7+i
vP8OLjPMeGm0vthwBo0ri2/B20k4FLdN1Z8Fw0R0VRI8I7vO937tT+L1X4JhY15mOBE8Cn3PxDYQ
HWNNXofad82PBVtlyeS5gizcwYIQcT/DVUeW7ey1uBRhraFjViHCCuwcHEosePB3yI+mZJVZqRar
+a8m5kam90YUW+Tnx/GK1eRPcVP2tnsKRAp3FVVEitMgnrqpnT0Ohe5PFgvUiCLYa5D9m3Vkl0cT
mGRlQLUdAkaC8TUrkMIMhkEU8sisbysph81xHgn3/GSBta7Ypwjwnkcha4kdn4ngiMZoC1DRCpcq
PSoS7uT2vxeQ4zmnPXxrgGtMaAWy8jd6ZTkLCiysdGq88maFNGxPQaQ7+pgXjrd4so9RK7WaGhnj
n57j12H0jkL1WA2d56AxhKOqg+9fl0rNviLZJO0+7It+YisrzsJTBIcuqEE9LLKcY+2/RCTi9Tf6
f+pqs4EvsO7F9R/eQK+KavGSJDBmNuuClqwuptv5o3ULaJmGxV2k4xSs/snZJmaUYJqaYh0ZIrH8
XBxICc1Js/zVedpu21eF6QcQSwJ0hHPQtplSb/cvMsg5SoONjOG4CMtZGDwGzpKW4z7Zv4tb27Il
hcKCUqK3uninxSj5OFIbIP4O1jyIh9M89eWWjJWhqRr6vMIAo85ShPkC9uNrgMwb0pOHWaufCbpR
KKZwMT+OkIlAdauPQHtlO4LYq9xeaETEfi2ZDD1kFWIpA6eDDVpTILevEF4ZM9tZSD7wxZKVSmMF
Xy0PB0i7mghrNdiDOTtc5dNHO+z8wfjhM+3jSb4/NgJ0NHYr0CWLcZz+EaWQnHPOrUEWnF9nzEYF
KUipRhsLMQOCax4ZmvyPKl4T51NqapNv0oS48Rm3n2CmI8OOBKhb+GUzs3+/ikevPCxLtycXtOXv
uqOdcmiRezUGtql2bHFlhlcFOikjBI/l7lvS9Kck+jd0Mdz6Afej0G9rzEUb6dJZpRc1v6ikgfpS
ULxi6p1SQjBKkIRztRqJHFW8QqexETskrpRYKNm03pX/Gb4MU+E1wl0YyaCsrPJ0G/Ivb9yHxwjX
IrKKLnCulfP7Bb+s3HSU9veIM701J7ry61J16Wwum5/DtjXGAnZOatAWPMzjlKnJ5r1z1SVHfdGT
KPM0pJkxu38r3CFkYF2F5/7PKFjUnoqi5mE58VO9vcReVKq9QAeyw811NFrO/JbmPc6yJpKVSAVp
q0WTHHcPkYaA0Du3+POnjF7mkTypk40z7xiN7okdfqO+pzpQcM50EgXpumu6BwEfzwmbgPcN75YT
gsAikYTfiqLvv6uOnSl97wNaYG43U6zmI55E1v/z2B5UD6acdD4aOpL13bjocxapub9am+iTrox7
qRiaNnJlMlpmb5xGoDZHMPwMJla3+KlB3fuh2CdPR053wTAgUyeCl4E8BsufB/7Nj1yMkz4FO5/X
VU7JXWDRlFtmc5jn/SzBEfgCnp01KiUvYqSQ7UuB/AMYy98VOkmRsx/6XHr5vP0NYDD17WB/Bd6f
MoZkm886QtBcIIir7Qmy4/8DD+MFqy6LDKRwYXa1rNPqvhuVBYq77otzIaH13rYdyhcJiJQVxBWw
JfK2Pwld4jLQ/HgeIcamyKde1+JRIsRuo2Z6zCYwhnlAJ5m5mGwEZJMKm74Zv6fwsoLDIqexr5uP
OG43Jq+O9lxaV4OQNpblZdmNX3/nflWsPia4g5Z2VZ7CivCH7TfuJ2/hWnFADCjeqPqeczDEwhPP
Vewb36DrAhOgHg4eELrOmXDJKsUlQAT27Am+3w3j43vA2ovyKm16Mh0Tsz5OyQcUH8TjiVFRIzLi
wfIQhrd3ks/heTjIlbtI2XVCDZ5i0qBD0iAUFIRcTnGWPVpJlqCXyAP8pwW4RhKzn3MOMQeYkFZO
VRYMDoPElS/snWk24pa+fTMhUwIU0bUWqaAMuvPAaOcAzk81Xyj5qTsi3uXvt2YYdLZe+b1/FBws
5VAd1HgnAAQ1+wPXGoLpqmY0n0IKusjoV1NYVrPGAy7v2SU00WMWk8GoqDH9jxRmFRb7yTSuZthz
g21QwH7i9VUVXlYhz56TVm8Q4FaBPSb3mzfmoN+zMWs4qlr1/bCfhkgADgrtLpXX8AY+/aBgSkM4
LNPtt4SBwPQiCRgcvOObi2dIASj6RffeTOLbZsjN4tCt3r9AmgZyvEVUnjqq/DBYu4TlDuedeWLr
MsDUeRLydsGh6NNJ/sIA4OM1gYdQxpTwCjMZo455xMAVOJkwxOmgz2eqRCxb4zuFVdGlMW87XSXR
VRnxixjsN7kGMn9hx22sbvXiOUHVcKSYebjT1eJq6FQ3aQhWSdvTw5+O5TihufOGZ3hP7ExMS1rC
98Smx0hg7UJR8bTGODIPGRJFU2yI+7SFm3SlAI+b42anh1ptXR6FZLnCF68EgOz7H9e2eC+HfYiM
EwZ7qzaCbwVqGUu50z57gsfUlbuYHer1Bs7tOevSj+Orn+RZ+6PCf6wtFaOWNU0OOjAWyKx7u5jy
NvBstxGJi5duj0Re38qjla2DtY79l8WFkwvWOxzODYwY3Rf7sToyOqFKbBZzKJ8Z4+kZMHCzI24K
yUDw5qG0BNlw+5U1kOPb94D+LW3Ofamv2zotvMrRRrUT1ebBpvH4wA8iyV2+75W/Ang+1YS0TDlV
9X96AHzDRuqPCNnmv1lhYPCUaIKZ82y0xZxLQ8NDOucQTJsZjoQ2sIrTDAW64Hgywo1Yo5H9XFcg
NErvcph/hRusnOlVw3WFCA5VCqvTKnvLk3H/IsHW4jgJAcwptCF8sE0FLcpouwzJZeTmk9w65xlY
JDP8lZWBbbKGqihKtMYWvNgvY7ailHEBgt0R+U1CPX4s1/kQt0g//a8StoYypDSQu7IJ1e/BHWhv
UYGJIdKEVo5v0aC9p1g3wXNuk7bL9qZBTWCP9rgGws7xFYi10Ij2zdXY4TOoDaW+8umrOJRu7HMT
fVeJPktHCFOhB/11BOYt1wFjyFZPd0tmq+T5qbyoGZ+SzCBSBU0c00GyKxdZSCQ8TCSEbzp/PH0R
+vn10xctg7+mlok2JQql48RksmXP/AXef4VqXM0UBjWUplixl7rBr2UttX2yRkw/Rl87A14CAcNo
sLiAQhyAiAwegHP2sj5O77Cv+Qp6vvFDgulYR2xhljJp5Cs0OTUghIXqZ+Z+9GPYUWWLayIEiAJA
FPylwDylppqx81SUTJPkRCSIMWBjR4WBvtIvNdGSePckv4ONStNtFwu9bSpMUG1ahzHViSYzAsBR
aB/8vtW43dOTY0FGJnshDESPMVeOmXvxjOYkDPBExUPVoYOSdLPInC6ZqSV4Kmzs9GuuvICY8UnR
Nz/zYG6MlayjmIV+YDK6C0awsZwmlio/vXRNtcl6leSaRAn/HWOxDAkuLL/rTFqJkJxfugbL/g3S
k0D5FXnGnVryHTzpFrm/wGDHXdzXonDNyhJ7FMdrKabXNff8kCzrsUytGKZqkJZpYL7q1WZYkpXc
vCahmxocf7IoGdIFzrujiMQu/k0mPvfbg9QPEbK1RJneacxMRcWk6bEN2098bThyhB1Sh0Kale4s
zbmzFs0LYyWtiIFSiuulPdi77oll16JE32tE/TM62vg10XLX3q3eLc6O/csIJ8GieEVuoFMRW5K5
9d+bvHpx4gofaD9y/S6PGfKrpsvrJTfsvBEoivyhnwkyF8O+IYkh5pgad1vhpMnXr2xkda0YxvbS
DL3vB8T2FPnI3e1ms0ryNKtDTc40UJZvt6pOhSpZQHiTyrS0MA91pILKhlIkgVjz2wNTcMTqTzJ5
PXSiWyrcn8Scb6lqvPpgBdgsQGOD0a3mLx1WuXn+sLbtQikS7b/AhGIB/iv9piUlEH8rdIRA8LAm
GIDj3M7esTHV8/lByXGBTVLWdlogRc+qsDsWThMmdRskcTiLxnyBLgHK0ff0Vh+NtAU6V29OrHKp
TiU95T5bBIn9qbxV1JFG6arFfwx2ichF9m/RjyThLTcmySfgYfJUrU1tQfO8Jf2ErOLhaoVb9pil
KA7Yxw5TqIQvqUrs+ld+e+9risQqDY/F9jHn2dC1PfnVEh8JSUXTi5R6DAWJEVLTTVyhH/BxxPxh
LSGxlAHBsMAu7lWWTQxwnaMLwTyN+kiJHQPH0CqY1PSY2KUu5wFbld7ZpVxwGojRdTdmg9ZZr1Vv
pQrPgnk2ZILiJn7mhDQG15KS6PnX9v4UO6E2sLovRGdD1q1VhXvHhNHUVDx8ZBm1Sz+6X96BXOU9
qCGhvsLKcJuuqd3njG7tRDdpk7d5eAva7ixbrAHhEdOLe+5GE+UGBSrhX8/3A5UN4fGpHOMkuxAr
Pxx/0Fy3m7W5T7UCJUN9SDtYHWw9zgEaO8hgDRIZmEdfzJhCNDnJlPTxLnT7+cTZgLh0gGLnGMDr
1PY8JWMI1a6Pv2lYR9/SGmlmbLajbd84SvGBKk2dGLxS71CGTRKPctIFIq9cPbF3BRHZCbm32Biu
HcfrvnHMOaLnZPXaIgWxI5zQafsQ9nEZf6UqL9kUfgpLwRSTGvUQgPp874QgRmPDOq9wH/fgAr89
+mXPUKru/sWcUVbKRLak5S6aa/23xkjFkpYr5QHXn5coouokX6x0LNmVylPhF/BwtDFFMwq75NiX
j0TJus0aTie7LI1XMDeBhFU4Y8FwF3FIn68xZdttELZP9j2UEgaxsjrZM/EskcizYE9Mlm9Ffa77
a0+A1a/6+E63NAeMO1Ue/xBTr1d6rafyDAtYhlZ7IrfxQ0pVf0OxeBUikW5QPZdPEXyBRcmnChiS
ilhPWkepmmAKeTHndrs1eWLYz/i99SzlrlmAOHc5DqKLsvilfCyGpaY3fjX1248lF27REbL8eneQ
2lfXlrhdyFzxrcHiRBvZ5Pt66f3jc68myFj3Voxrc2AvKjU10mBCj4zkUggGqWcxdunWTDwlaOCp
gbEUnjRElG1K9OVZekkzSNmW6CVofNmivk1Qv6xcPRpJj+subAUZbaIsMmjcDPcEYkDGhKhr9TGt
hTN7mz0MCaetAlPMA5adQ3bH3GhAD1HKwct/GiYgbQnoW7s85Tr2BQbN/9pQMF5G5Z14qp/onGuZ
7zdC7FFXgErObkDW0HibV5XaT4K3TCyddboKpBxv0rJ3tkrGjaSKaQw58G9OmbdcKo4dpHMsgHzm
yRFbS/BGLlfORC/gpx2iHIpjfaGV8xuVXhDIOR4DchpGKWe4tTDMQZXJMWO828bFRXHta9QTBZDq
Sz/Vl68SEA7qMEuKB2DOX0PjwtShJ97TtesSRdjSJyzfl46DR/CFxrFCy7FX9oTOUgg2BbiRPy8r
ncoH8oRAHY1p7nsxgwN50IqfFWadbpEiVSpfSvMhSuzRQ6CVUu5D6T8MSAWk32G2afkYvDcvB6Bq
9Ck3X8UEYgrtmRCAHFY8HK50+xOjDmE5t4dnB132IHML9WNnullP6Cnm5lIg73iFyadbXxuoBj2C
cZ2wQYf7xfpLZpkwXa3PpPFbX9mD+NLpw/abm1cBVlvAmcRYDhLO91YtUKHJP3Ls4/Z+uyYDo32R
9VeRr8aSW4e/aQ9TNK/BfaQ7yfmfwBIdedN5C5/lbm9uwxooIIuTTjxqdsSsYFXbWr2iOLTVOEmV
YlHk9bp1LJxfrXYsFu1nNBaRkb5e0V8Y7uoiv9jOJa3NJtKQlaGZ9mAHnt6OuUhGzbN1EHgfaxQ9
VSVmBOExx23mgCiPZqw7PhdU8rtUymNUMWNoJJgQ89Kc+xXlS7lIofCznWuShtwkn5EUo6SYGZfF
WLgq0CbiDy77Qcz0l9Bh23FOt4XjCFiowbfVjxFbLMjtTma9SLPMyN0qmCEmMEAIvtShD7yuO6Rh
q01Ayqm2So5Cs8N805gltafQJko5dvj6XW3IOqBXUVVRRX+0b2MzfzX6JLSSwig2YjdmwuzPgHZp
icgpOJo+EEUdOblO1TPTJbmvrDXYvkpD6Nwo/0B6kBry5dkNvP2qz6e2z4yzLC86+sxvQakfET9s
5fBJ6y4EhAX+YXkJPCFsZhOmyIyADSiQXRjvlYj6MLKU51jkDMJAbrJKQoMfwZNimCTi8sR9Tr5M
0h3NYhs/jtKcBjgev7c59xsQfQNIoK7e1/sqzbO6IaGnntfY+rsLjp/uOSLv2H1nJdC4JMb9+hp3
jq6Mo9zv1iJezTUL0MiY6YO4XfU9pJiqLAZRk/jNt5BUymz0n4xkrZZmZM6dyMWgZBG6nnZmPlXr
RTrX7/YZ7wwny4oTY07h5kJeKmHOW1mHGPipiGmRTFnWWxhGE/LkKJm6nkYziZHd9khPomsB1Dh5
FQ4+muZaKqtXRL79LA/RPlYfUKbCEYu2ecCraEpV4FYHPgyNrquJ5Xcjizg/X43cJh+j8LxKCBm7
5JkbnAlG2nIqld7ZcegVm7/fPU9smdzkKU0Ab3402/Vmffn4i4R++kRhnzvdWzMfpTYV9mHkK/4Z
GyeHTS8UqlG7sCIDpjXZefCAbxZrBqDQAouZl9ymAoQ+KV++GwqZOqrCpd/pQE/gPXCebjoMuTFF
3vj4bODGfISqmaxuuhXhiw7LgMBc5HE8LXoUZ0NrnCaGNM8J/HmIFXjTShlvFWGyaLORi+zo9G8z
VdlWRteRXIz2yQDX9J0sTx/l9T4ssjY9aLZSRbBA5GELKfhiNzM2rY53vp61l5YWiMfVHbEkMbTw
DzNtDXOsPuKyRnHotb+9yzlJdu+6209L9djMjSGk9lJHqEhgjE4C3TT3aYRIdrYvU6/9BAFrOcOK
yeJAujbrtJZnBVk1j+shFOX3yYoz3mVlwFJOFCR88G2CklVs334o5zn7GJTRfjteTSnX7sL2UB7W
GHxZelU1iooDDPmUs/NdSg0QSi5v41vhJ39GsiVer0R6PywlERf3d5g9Xh1FMlGcvfJtlK6mY/Zm
OhcAlBK3A+t/l+aq0ePnzX/dipk8whCDhsdiAW52BN5UHp3+VP879ndVReCOIXrMTbWf1Ti5FtE8
RJZcmwY8qd8Uo7HohKuSaGLeU7Z9BsOT1wm8gR2YcZUfSVBiprz7iLBgFQcrtNSCk1b+81tMcvLj
IuzS4CRi/vRNFTXPVE+Mes8Kf2PxVt3oZmS2crEzIzwkx+XS3zdqZhVpOPG5czncGwJ3fPVRIQMQ
QngK5S9U+wsJAg72Ux/fM6ckwX9fqWObIBSwkwiVKFGhxa2FM3TRRGQWYm/krw6OiVKNgMIkbZaG
vs7VyNRlReYszn+LszfI8sAiM2TuddGgOQZX80D6RSMKyCB6WsX1AX7kGL74pJonaFygvuXMppF1
rGhzu5r37jUz3srjdu5vdEBxgxs/ccE5EACMF4fBM9V8rF3N7TWSedLcqf5I9f3/23+LVVmf+U55
LjNNB5ixq24R7LIRC0xbR6qsEgqDdRjU6aPo6EHfnRubIoBS/nhQFv6p3757IeXu7JrG+n7+lwaa
hk+7wv/wT/ThShlciFNIom47qSE9eQ39/xRMUX80WUQud28mPoVETgSlkxsEMuR1zXHxZ55XcAvk
nilj+12N4liQOoYu/wqWd6tzAvOQmYGc3yozwVyp1pIMH5drvuoLQDhHy7kEZkM0h5HLXUzHIdrZ
6W1NhgJKFv2zwvYSRJkB5sFBsVRU+q+nPytm3XzDX4N7kz1BDu4Izu6rw6OlHMsRqDi/0VK3zE39
hFba+RrcI81dzL1Qxne5toY+te+d8IgNVsMUJxgpjnuV5qDTxNzmPuL5CBOS1M8jbj0eK02LfsZV
Zm39iNr7mxRWsKW+XOIFTbuKnKcuWckpwtfEwXESd7k8WKjFrJAvoHvi41CN1VHXKq4SMb4C4lI7
j2B3sywSYDxzcHrCUeHZxiW40RdWwFUjYLeAP6NW+trz4fZI1Jnih2Hs3DxooEdFVHsZJw+Og3Lk
1CV/H2u7wvNIGO7GiGV2D9/IIZwH3lIhY6p8n1EBrXR1JuLaYtLuR581Gl+NvjKRVZgrSGOfENRN
ef1uZUSk8AIibDcylmXP++vm8bVTHpSe/NwKTC5UdqANaNm+qqU9nzkv4HZ2LPwSPEKE8JMUmiPk
i+cIeFJ2YbuMZFR5Xl4yxKJQ3l4EZMdLHZxGa1x8w/1MWJhLYJMzwRlKVaXuEm7vVsj8vv+6Ctda
tnZFN8XWI8T6Mwg/cvKKlnuqFf8lViZmy6XBKqqihqlzbFYLv9rKZk50RtNQ/D+mzTAW31mX9UQx
UKiQz5gfhsNVxCnOjfO/QdZ0+N/l+d6hT9WBzF/X6fEIdnz6CYDezcaXVk5+a2FpbLRoWSIDuuRe
u/A/R3DX/luM43gSFVk8jHBNJqeyBnIJcm7kFFR2mAePR2c4zIJXw+ade+TmAv8zOQwwwYR6Xy6g
4WLKawPfKmvUIdRKh+R1C23ZFZud9cQDnzPkvcnctkiqldbQZnfR+ZY6hy+WhjcLTiXxy5LEotyn
NuANwJQJb/nmxKFFiA0AKDrTYtN1hoRxhjfB7zpxZlGaBR9I7PK2ba7EhCR3/7C42Qsb+uLHm4Fw
Tp7xoTsrTHSNngfdRg11mXMVELR8VIpUpTJRdlkPqhyWpHHh9tNXAVbkp51MmmCH+71JCXnPLGzD
ywF4wad5bA8cGm8dJdgaGveBWBaeT3BOHZXeaLFBJDcoLCX4SZyUO3tR9ZpSxkyAMNhfZBBdN/9k
0vHIHsWJwMAOWVwuLl9oGTnv/0IEOOYcK9YMMNeeuvjIe72JG+d1Bo1dVRTO79locE8sZenWl3P4
e52t/mmxm4UUARE3OuF3rYoKABcRnF920b6mtBhOIJG9XSPDyGvJNddlX9BuRrbAegSbiQZL8qpw
Wz33rKp4v8/TPOhOMEgrPpj/LJ1MQ4JL/deMJ7u3oQeGcEy1WuR77f6Yn/4t2PWdnJawZsL3VqVQ
S0iD1STs8FFLMjGNFAWDCfgLFySSNIT7Y8R3QJWpLz9VbA8xoHawCxW6qh/3vvraQpHW2vQ6uwC/
jhniulU8ks0K5IR5o2H34qHO75pANHASPrnEDejCZo/9tUK0I1Lj4OuUdDixV6XOM3h+MKaEyr17
L7tkkDseU12HTQz1VJXvI0ZtRrH12C2q7pg29cbMVhDLMxyFMeXlskn2rFU6ETcNkp0kciFnpwg9
TRX7zs9fyVlSuXRnv2vEUidcbKTSTR4j2PwRH0BcROXo8fnevJ90b/ip/GaUgMLVck0+yceBiILv
0dAEO/J50D8Ho8NNDH1B3I4pI7O325Yr9pWOEjBh2hmPvjWVUmxPMR0VdffwTfmvqb2E9LACAvMd
JWDj1dG3qA4vyrdkAoG6/PjwDx+hPrYGQn7BS50HwQtxWxVaFL8NLumBJRBS2DYAizXCAGUlDY/M
3esrCFLvgSCgIRqQE3bVvgyopp91E0BvRwrz+BsvSkb9a+Or/SG4BBYXqEMSgiBNkpXdCb5jblAx
wGhPz8J0Y9FTsFj4JvNA/Dw00Z9A0Kxm+OlWd5+7JdGlda8gz8iirZxbmzc/+T3dNKFKCIOdYtju
k01ngoZ/lzShi1anHLrzto2mjGwnr0IBnuz3MMIVA25DwIb8br+gca8brlsKWQYt2s7nhLxY8MIt
prlOt/YHuYLjBupHIYeDtNF8iXNabFOAjxYRnssbkABmdBMvIabJ9/UjRa8EGEf4VOdkkgSx9qYD
FdTc8Z/5SDekJmYTXrN7d+/jSJCpWfRnGQ1gs81fynrOyYn3L0atdGr9RPbdwtweaP+fvDnkwAsY
2kupPgxb5qXZ7T7YXaf+YpQwsgNSl2WiKplptI+1FOngMBVIrAThlezpF5q5kl0MUvgQsgbXgSyb
61xQl9iXofK1KbmFNT4FuKmTA/7d05kaQof/JN7UwSI84m2oPuIT6q8w6aCNXqdaYTEq0xaCvOTS
9NACkrrcrabIvmPonF6WxcMKY12KbT3ymf0xVTENlzN2QAMYt3pfceR4PFOgbG8vsNGCV2h9A1ox
HnwoOTHlZeKDJCTxwjwBBnOvn/U6vkQtjTct1nYrXLWdeCP26TaSdyjWwJYFhXQyUhWJMvdU6TDY
aGaTR6KrTVa+eVFBMurRGfSAhVWRRP3ksJSHvnMnc15ouAd096TDqotlJX0lpPtV4BLj4V3p2wCC
CVrH0cOnOe2yfmOGjm88EiVV5Xt7oPTBY6NGvsmrSXuG6Dc6inkLEWKKi9pSLN3KJW9xtYFW3ZFA
VeDiELG46wfa8wDzLhEOFTW6MQFhGkeRxCXA5/PIQmXvegnBb2WDDHMK1tAWRaCMGIgBn+j3wx4b
8LAUt5Is54xSsND4McQuQyWg7Pa3hGzYBJDeBZiOqFM1KUtBJEP4XwvkEAE2ToFf363xtn0k+l9n
3EsBZoKeGyxIMoiKeX7VVYSFJPxFyXJOcQBV+uG7cx7pR3/MiZbG2wXkfitX/jkGPmUKDlX++FCt
flsCIbv/r0Ml5s0gyba9e6uX+eqDT+vIl2IXIH5juuVwVxoWp/xENeM2c3oIg0GaePjqzww/8Sr4
itmvnBF3LfgoLvs+4TGJ8bYS1jO3spTKeoqIwlFFEoB79stAQHAcp/2CJ3t9NkS9rcJp/zo09S/v
ChqQNp8eV+ucCXElNI8NCkLUk6lXqRO+5A+Pvlc2JcMMT4QWEZLn9iPqZN5Kwr4w7cRRCS0Ii3ez
Cb5CAMhypRgG7Q5XVJ/zrW6es90OJ6W9VmMb5kFmgSfmMn7AdfGQBFbLrsjEAV8BP0zCXo1frD2M
9w4U4ujqgA7OdluTX+SyZn5WTEtJmcqqaTE7sJ253AqyawMYOQCK1rzBGpWBhLoVaeOb+i3C0nVj
+V1YEMg5omIsWzkhOpEtz+NGKWcS5bPpkGtcyAWxbYi7/U1StG2qyoEeGlhmndz9pv9JjyQattW+
Ws6wgV1dKX5xPvVtsgXXTmc1XN3gANXc7ni2ppKUNL6L8pJTufiQ77jKD5XYsj/QHxdxUO+Vzy5+
dWjBU+//JB2CtUr6oA0M2THAtdI2+Yp/VOOLLR07E1TdvQiADFeN0oOkfI+UKYoFpHxOSgsf/FDd
Z85Yem5SvL4UyZfDDDER1aHawDO/bwUKlS2b5jbc8BJwaVHZxmsl778oAEIox7y8aV1HRnRamAd7
g83zZJ8vECxrUsg+j+Un0eCr95jK8fh9mEPDzV4eHscDF7/NaGtpBH6ayjrwPpJGXGR9qtXOFLHG
6rMbplf21Ujmlrwrv+i5WOJCjBWhYv2e1Ki7/QJWDpO+g7at7iLyttRzoxoQSHo+Yq6ema/EHw/T
iasY4ZOIzlACCoK4QQxS9gEiVBwiBBAA/W1/sJYCICFIhk83Q6IMWpqPcr2nPtZl6G1a5+x/pZkW
t9VTYuzmjzoH5lj0/SI5p9tVaiRDzohLl1I6LkfHYv4aEkXG6VEQiKnad7kgFysBTDFNV4yHhlx8
xR9IUqgin5oWE9Tu0MfqulvZCB3PJ5s3+S91cWhqzYaYgGL7TkGEKovRE/Nrz5lpI/3r7jTwwsky
hdMq5v/Q4oIqqAEYO/So/vxEQhRwDRYQXtSMWkfyRss0UYYxz0wctjRBi4Sb6fUReco81E+LDyls
ZFeHVpk68ezkZ8pXlgPJU70abOdhphL1PhyZCH0mhjmorlFiZeyndJMF3EBFXky1/fKw+yynBjTA
3nyTUAYIpLKs4wWw6gA3RaUDS0I87Lbz9/mNp9/v4kR6MJWDKeVa8MhYKfqwrfYxzeGsixUG+jlG
++X98ZnER3gQU3lQMya/gEQFemNxjsSwHR40YhmfCjKOTgISLFFVhUVXR0Ad16ajVqU1btyG2yf/
e3+fv7wZjwfnNeqGc5QtLgtNiwh3JC9FM1lLzjjqY9eg2XA7e7f8xrh+BCCTVCCdxDwar5phs6x2
gjBAdbOrWKobxNqb847XmDhgqJaUrMSPfAMcCr+KO1BY/XuHdx9Vbp1eAkFPJsWAv1pXArxGnz1M
h3BMee0t04w+thTLi5p8jUmJjCOLJQ6cFBS0R+WX3sBoZaZM6NpymdYN1GV1IeH357RsIfn4u73D
smIh9GgIkmQAaMF5ZInBFv9TSi3799EcFiGnTNQXuj85ghRDpVB35UAfoSyj5bMVpRnS8wdLlUHT
CjrY4cF14qF34wsBm35vqJiy+x+jZZYoQmM4qWzaR7YjotznBQKRV+tEOJJBNA3t1pliIYGvO+MO
18FmHdOa/Wb38Ctzs9eFDTNzxJa0/UAqJrBZWANbzYRsJXADztxpdwm4JNtkDn4BC+BistZUMtTu
QRBP0Ebh6kuPXaAEYNr7cFT7iAElNn/l4zY8jonFwviCTU53/M91gIHhmD9zB/frwllxJ4qLOvuS
nEQeHG0WugMZD63+2Etj/uwVf/NC1T4Fus3K6RlG0Bw/lbyKlMqynqCvgU1DgL6Z943X2+XrnoD6
j8NZWTelvrnwOkcVpxPYoY8oZ59F9Jh8Pav6J50J3swU8W2ThKDU59jKBqTxv8CZZymr0lvm3+LI
FAPL/VsGdE2rLeN9OYitCJ84Hz/4dGCu1LOVa8mHrDaAB6LNpl5pVTFh0KjNZ2PRPBWYOSVnI41N
IfpTmRDK2pmBTBup64hyWF1FDzHciniFEJDk7rS9GjA9iZMdVOFkSC0gasYCFa+HZqd7RAIvRfId
bA2BIa+zWBXBJDuubUSSDAXjxilSd7eL38GLtiX200qZ1Pk8+dkavl6G+P5qqmxZp9tqW6JxqUE5
MpNo31bPmeHx8PCeMp6C7bl46nfzqHIybm+hUehQT/74zmWusJ64Jqt+c4Inlg6Q4Yra6neud/DH
vDTZtwCfHDf42O/Y7H76g4Z9b3JP0E90CdI9z9JVgQMIbXG2BO/BW9Y6njKpQNL2xLf8rUF1a+eO
V0DnmL4hkZswW5HJrVWhNd7vzy7KsGMIcoiTufKyy/KS7/lQ9C4FImzV82wq9mtNvRZKLpHOluVd
IsEAUJE7Wfa3UUzleWbcQdHJevtp/igI85AG49I++h95hnN+hkbLRwvzIreadQncx5+2iCbM0b0I
mXvA/39AkRao1R4GSfVWpTJz8CM3Tk39//iEwmVvD28h/7lENM38cDkzIvyjL1pgGQcMcGRU4F5i
pH2P6eZ5DCYdgMPAjVaKi3+OoMcMA9p52RUptfSUw4K2r7YSWpnuUPZFV6RycgM0QiHq/5EZu49M
qUWmnSN7ZknRHOdGkzX0XWsZMLR9iw4h0wG++BPD69s+gAyBbTw6QSCagCZF0MpOk7ZayATmQt9K
BWMVlJAoNKMZ4jNBREWuFheZ0fz05JWAY20p7ySroI50KvUQAXGtNmVewbPEJ39SGIYNl8SXbcHp
SBkCmiTpOYonDN1aUcLFECXNuraW/Q1aCGj8f3jiJNLyflnR1xHFF8NpptqzjtaZ+kOEeG2Aw64D
RcITbphvcrMHl4s+aRB7xLFc7ui2Gz78OyWC07nHOL1nh4nteCTp6kSuevgroKpWPHbcEskT0fU5
2dDRBAICGeg8XjLQKJ2hIfdJjMbqe4Z1ohHddG3olEuhZ7wfkheBgTGUjI5K9/i+q+SCrpmQ56iQ
gzt81m8agx+wBHpm4qqL4rObatgly+V01AhfvxrvZIR69+VgiCDkrPZukT65mln7k9m/nAorbxBL
RViAhwNvktcH0HQhUHYyU65LURPh2XfGwo4/+pFzsW3beqj7yP8qXueMy7fcLNIT1pyTp60oq3Pe
GIj8zQUwm5RJF0HLQwhw/MS7vm1cFFzQJ6jtjrm+zrTqoCnF3oY8N6K1G3FUHrRMtjRqIPVawUJe
2joQ1+rTpP+b8yiROJPcC5S/a5CdrmieQdI9aWmjgIVHAwhG6b5MIuU4O7d+q/bCuJKUSZjPRKA5
t+s8H0ErQdKwV5AXWanqLYLqnawhdVMl+sJM3FMJHSm+33M+mzTTKqvgW7iRhDi+uwa/xZ+L9EA1
kw+/H0MRyysbl5oaFC8sO+f5r4xPOYpL8+7R+JiaG6fJaFOuPp1/L5fzleBBHPp6li9ofZ6nEgr4
Vw2s0U9EmttfWZXFY8+dBBAX+3Re+s2XnWGsWijT+SP1nHQCgbPaNLHkcv6IJmk7NMysCj9izNAw
ehc7pPsDckCb3Ljp6rhpZFWQF/dx0hkdStLvSoVOjyR6Q6HWUAJto8DnggXnlsXmWYqMhSP0acem
m3yQ8/7fcyG2yEMcl35eeLCQs1UiT1EGoE97wx4jApLcDfhD7IvfUCne9EUj95ZL1ZE4ptrH51QQ
mQGwRL5z4y/SEzrPTI6ZbGgs1SQJvwZ7ycwIUoilf63PX2AnHRaQh+rNulNr656jWdWn6uvVzFJt
C98JI79ZlK0B8yPYX4SVwlP9+vDPAF4T3uTmZgidPefgze+93eCLbWnuju1lCzl4/4XhxfJs1YBv
vp/95VjeUjkmsZBy+Hmmgy1OrcQPA8opAXYlAZlyscgBZabvAQO3QQYWPKmm3KLw9m+e3pO+B+D+
kEye/lHLh3ooB1QSHi0HkZ/9PT/LLoW4JshCffSoRJpXbSxB178aQsQmO/7rPWiEM9uOBUGIzSQ7
+qFeZAS724Vyea3D0BcpeO6s16n6gW8c2p/pufaUHOJjUnmaS7H2RAnjyjjVILDNqwhxEym5mf7C
AUm5znvAIrP/xEnjnogHJExfsiIXWisJcnkspishXcT/bbKPGX2hwINQfnHoSb52yh2Dj9wBlr2i
udDGT9ToluQhTX/Kko3Xk1btu3AkAqrFGdUr5umvuWaMf1pmvMN2B+llyDUjH3Ng1ZZbMcAaYLfr
mniO6SIIWNehN6rbfYetpw59xDhMQYbRD3PFF8OmoTW14dSbnkspJ2C0ZcxR0HNyvkvPwBrB7iur
Ru7Ihreb4G2PTjd7Ohgbof8rE2jR889S3PYbHXb5WW/Zikd46APY0S6XzOSUyPm5cWn6+Kxq/Qda
etiZbX75GQHu56PDM0SP6P9EE7N5jwzwKmlzngSepdmXXgtlDZNOjEmFIeNe9hC48ggZK30kf3Xw
YSAlmvptBAO7YtqYJMCFXARyNlFnLFQmwLfPrG8Jey5FjvXocAWoes25iGO2k2wFugANVDm18Cm6
8MeYHos+b2ozP1RsgbH5qqSSd7YjS3GvuI8XLB79F7Vfi038HS+vN94uwBdVtrfzcYDfjAybpDRa
WAN0D5LnuyiB5JUm4gmd5t5BD05dVnPi2q9ei3rJARrJR1LiNQqz04G6L8OMCsT35qjx8g+qaEuL
1PhxZorMuS9VqkboSaQfzSSbEpg/QRSQ8z7kTap7ZNLjfo/FQFEYoCYMuiJs84REPPPV0+mayYzf
gfw8rm0FmNuftnWEJ0UVg3lsYv9bV24wHsNeSe0dHNloN7HPBr0hiSgK2aQmCS5YNw0WLMqMYffw
dj+7lMw7MVrLC6ly0VKK6Njfe8PZIKlWPVNWXyP0bOGTDUhurJkkCN1932BfnmZ1AyU2Zsj/fPtA
96cpSY4mmJejO4f1M4ZY6EiBiEyRFkixUcv/GjAD1/vxkHnsdHRrN5ub8gDb9JpvWEPHFWIrpbJa
PaxjOreIe43BVwU24OELtDJj7TtXfgSj8ogMwxFVpawFmfWHko8FFvC3WvLafT2bdd8Bjnk+EqTt
xwLsL4mszvljVBRm5sJCqYc8R6fXe4ejKaZI1mYTY1VE2WvX/GH1eZOaE3uQ9YYbMHfX6/X+AKfK
+q42DLxUmduBKJ67BUP60PuBnL0yQ/rjSCIEvn+DEtIJSBhlrXgTElzSS7C1PaULVL8X6xGggEvh
Rc9NS6Ju19I9lsLuE0JPZ6a8AyPJQGVrhyaVdZmcidyMoeWkaFiJqjkpBWrE0aueupOaRj3rSe8u
SiC3P7YtHAdrUR7vZMJ8FGCWZuSBjWZRsCQrakGx5le7pnhCqmpd7wNkGEVwQ1bbfHYkVfthbHWh
oDz/CXVZlCKCzSkA8mou9ryDJlEU4TB5O+AJjjv1B8542AAJTTHSD0v6GCRiWwU8x7v1KIiLuqP5
jxScNBcRmpBepv0jeHsF+U65kZWGUZribMrpoWAtrdtbl4OXcMOZIuuC4xQc2baCtDDs0GcQjxuH
tdGloz7Taw9e1TiZD4ODjPtQ+HAR0fRCdkfg0L+hv74Ws3xm3ptLNwgqkw70Zojwu8CqVniHre7r
M+fDkXZH+g4weirrSrrzjtOfXnEAo80QrDLXZBlN7WuwIg1j9s53QV2AvRN2CEfFR6sMKKpOZpir
oNk2AcXiW/sT9w6/cXVq5PzyfIBdUHooffUeBoSpglw3zmaYJJqqdEekW8XDWb2QHOuEUgWNJGJK
Prfed9ii0U/s7QJ8mDmBicnzpTDkidjxiHLimFhTtTxyoatf8PcswwajPPVfOkIGyU6JDmQMJW+u
rnCvXoMG+Yqouj0PmLbXrN1xVqsmOTBZbmvM+a3F86leypqKgJYSiAbM+CtSUZkBGPBCd1EA4pJt
+C2QQKr5X9smK3WT1P/bVDLFANmr5n58uA1SWKK4PhJm+np11yuyiagXV8ClG2qKH3PuwaxupLwl
1bQ+LjtfMp3i73npbtYB9MzdeX5VALZlFZb4kayXoiGY9LwqYC+PSVwwUeSP+RKt8dtWnzi3ftaV
CDsAZcVTTgcvoT5hK840PvtWipatdOkMO6P0csZVr0KV3Jhq1Gpg+7uoMiwZ0pwAC3bP5pwYtlGx
x67Uk4yKcbZzfVuzwf2OrHZKoABNnDqhtfPYdeN6Xkc2Iw9XKEGtncPJYt7WiWFVaUyYyJe+nwTC
oASaldbBqwBROgL2y1FexS6ehlSIDdV9W8ukm0ehlllewZOjbWOBIpx8N11JiRjvS7JaU4xNOWoI
75gL81EH/A0ZDfln5t5a5i4EZ5PRZ/7pj9csaQUPdDZF8ZCyy8yOS6ID6HphJyQRCqGHJNRxR2Pv
OwuWQIec+nb3xwh6wWJEFNj0FRnE1sHL2wfiErB2o2B8DFNojc6H7/KoIzkT/G2NdewB1+LYpo1x
XXDZCLLf8TIRFNEOLk4VbXbaXmhzCs/0SIIKLkn5XMZ15F6d8FmuJl11a3TIjVn/aSpVov8hmII4
6ZulW+Y+nuTZ2CQl5KU6z/KlOYYjaQAzUvugD27B5z/0v8O6Yxybv9vwewddGX0NOwO6jA4P6NLF
1Ifkn455OGeC5PlohbxaLmmzzbMn3SjLJ3RhFqgBfnrPLmSTFZ0Eyjpq7Z8Em5oOXG8gVZDc6yWj
Eu/MMtVRFTzgGBSsZV6ZGHv2DAeMGLTCJgEPuUufGjNfGfNFfHS3nmIrDJ+qdfrLo7v/2+H+ROoM
q7yRJ5sOL5uhq3p60XltKGj2fg46vLrpgiHw98WzhdGghK3MRP8R8KkOgnt6QzCQY2X75l6lYWqG
oBPy0mWw2ot9E8+qgLaUqvXuqHLUMX2+GLxU+yC5mBK2NX3MeVATq+3/rN1gqwulfbSYcofNXeTE
wmi8Fk5mlMTmwNVKDKyg6oPQUjDbXgoNpDojRr4IHqcIiOxbVztfdRxfHknPB2zXAkFozLrPkxar
nB/CQYiYj+ul64Pdl5I/d2Vjo/+h/DE99sHRCMj6dxM1nGS6Npp3SjyBQFw1WhoTlsToYCNa3QKC
FETcgawiUJP1291AyDcXq4TRmObjl2EQfZCBL9gHjjWdcVQZWO24v4i2uqhATxWS1+nOMT3vFJZe
GBgW2xSaWTyL5Pi3A4MIHGaCM7FV72PuBxRvg62lN4BYlUo5Lppstm6zrllY6wMtQ3vHA74bAmT8
MUGK0NP7pr/GztDFFkQtR8Cm6iL8+uId7iNw/tfNb0yMWIgVnh/aswJ7yrbnRPDoQnQC0iQX+12I
414/WuAaYtmw3R10INC0+2fulgSvO9Px69ZJUByoO+tQtd0WMwP5Hgw+NVcnko3EN2in7Pfrev/P
RY17txyw3itECKpeFDkp3Yqe1O2LctxoTO1WM+y8E9snzwIfivrK98nbCASyJd8qgXVKE7RUhYF/
byTD8C1xSitEGtRpEmZvTRmYpMUR9N9ivEC8Qxa8/GWwOi6X3bUlixANZRNZr4uhTaakbWJoIBL1
7iCOlpLTa1So7jWElMWnwujHsiKIB4o11q8u/eLhsvGEZDA5TakJzPA6LPEqg4JO58IjBl4At0MZ
Xc7TeagUjXn+E6Q4q6aiI3jhL1XRAqfCSVB2ULB7SjnXIV2bWBtCDvcsw1hZaoaPJJawX8ea+wAv
TQ86H8CxD7QBmM2720GfXR8cPqKvhzVh2V08WbTxFfRsTpmLZMZNZs8mw3tcmnWJHdQxkjIFdr++
hDUdxr0V04LkSTTwjsToKYoQVzu+QLPudx3gCqmnU0L/BwAoBLbcmcAN7I1J+sgsovLvow2lFWOT
aktrGTS5n5Qa6AhFJc4khUZhjPR9CQxn4yHL8tVUBuaYN/Lsq6BOnwc1zr6iiLD6UggBfh3qah90
YfIKFni9exaDdydg1w/7ElzOuE3mD24XkyQ4mq8CidrlTF5k5PbVV/gQy3sRS4SRPAj3utPVaLQE
v+M/G7WsoW6qIKPxROGU/sI9QUsPit2K55awwmaJnn3ASmAKxZpLw6OCzcPSCF9JUpK7GLSPQMYU
jhtQ/YyKbjIV/wco6AJsn2qOdEh4gNdcfn19rmr4IYPD69eBR9MZ46rb6XKG3BFi6+D+Rx2oFs0B
JVodxziRRDmcFKB/WDaH1h0IuGZknbWywKwh3VnTlZGtzFwKV2WQceEbfQFaPqpYfdsGuE4+Fbqk
6MHbjJaH802V0pxRAtvXtrw7QUUW0+Zj8T4pemTuyEzwMwv43xlFT2X3EMwn7py1XGUa7rDGwd0i
TV4ux3uMp6q5oPoieR/lBZtvqaLMO0wPRqtBCzRcBi1rw55M38PMMi9wy/EtT5JKdzLrppq3Hs2p
PxFQP0454mcyK8f0FQm/bmWqcnvOvSSLf8/hD6hwlO+n39SKjpIbtglNXcV9GBiWLzvhLqTNIVge
Q4N5kXlBCQHNMEv2veoxkKTFlcbJES6va26YSUkSU238mLTC+YG3poaML9KiVjfFn1F5weVN7e+Y
h2k+S6tca4JuhrSO0Oi5db3Azn++GyS/Vrn8E1qHEnckFYkPzkhCMN6jgOuSWUlCUQ6KSYQ/tTp+
MtVvMXDP6aI770tCvjdKQF132U/kvrIThqbl6NTFoebWzrPcVxTRfr90bCIr7VWkaoPri8lPXRqx
6HHL/v6DHzNn6mTBlIST/UAugY+T1iq1+xQV6lZMWyEJ2B8jvkWp8tWdfehC12S8Bw/R71o0K+KU
AmVhFX0Ql3/sUnTQbF7UcNbjselG1nT//zH5WFv3Sl2cDTCqwdhYr6OY81+H27anHptg7RxDQqeN
aZd6fMK1IML9wqm6Y0H7uug43WTKH8FXEfHTeU63Fspn83xaui+B7LDZqBCy98xRy+x7YdTK9Jgc
9nrHuwcmTXuRouUT52WXCaSVtiegOI91PCU3ydSMTvwc7ZBO7d016w/vVXxhnusi2vAqAdYT2IP9
mf98C32XT2621MUIl0T69G0rFqAxpriHv4rinJ1aTuNtDhBc+c4qvxECVgGAgA8Wv/s3Kzr2Elih
RpYpHGiafTH9WziSQAeMfKH+Sb1txx6nsAUkZ+1om5R71eDcX5gKI+FS6BNb83jTlc3OZLtpOcn4
Sf0xs7lKn33v3MaheKy13e58t7rZyDwokQz0+kx0TXgHVmK6LxsuSkZGFWWCy6HWNNp0BJA3/MfZ
hHTPEJN14Vmanuo1+Z569WffPprxZuCk8VIiRqXC0sLrD1SWKn77MobRJvRBK0sc/XrIKZEVnyk7
WSEJDBqgAAJnBXS6rf+sBwVhs4sibICpobS6YH3f9wp4gPyPqvxbuolwZSxrg5rTPqx/KhWSsm6o
I2pEWhzkdSVp3xJhX08lBOARnZVp9ucXs7KcaHK0bchcyKePKwFro4pXmiGAqpe8s615Iz82Gapr
jc2QpkpOou+rEC68cPw/izw5xrfTsQiDSfBO5DW7hkaxjaLPFZ0tGImdmIIYcJKUERWTj5Ss3Ge5
xh1Wx/iqmuc30jnVCEjdUQaJJ/iNSvl3P8HRei30NUXTOThtLDAhc2dFu64F6rW2VmwePWSFoKpI
ex9jwOWZaPRkoyjOa5JdDCSkWDgfID8E4ai96gL+3vtXNYV6NyIKlu/we3X+1Mab7iDOsuNVrkcX
4URwdorIkiH82qMADRrfz+Jklsu1uJVFiqug5PBGj4qPt5Uk21ocRgJN13FP6IPTiPcOa+EwwKNS
L0Zwx0Sqi85PhCex3UQDy+OZhBe0vipHHA9innTEHE3qoKxcoi4kmGJDU1Fk+gkl4NWqDsbdza6J
jzrQ38Vfg1V4CwmZUkh370SimfWqygn23aHhDW/LpGzv8vceQprfgYd8u3S273y5CEit5Owejeap
9jXVbkZ7KR99CVK+8hULZP95ddakCSNGmqMk5gmPVf63r9aw08bX1uvwRKAKDE6NMAZfCiQUMSIC
C0I025crDkelo9knAqbek31LTnetIB0fWL9KETVTwqb5S7ovxeHomhEjeoSXOz0pvf8KF5zj76YK
GpxnuwbSlAzOclcNLr4B4ktwu+FpwUK4C9NnWietUu9ntUdJC3zpWwn2KxzxeRBNnbeCAabFofNu
qaibRVd4IDJSWfKAKuRscNJZ8eb8SW7qGTf9dac8i9wrB4qh2DTYcr4dgHcFrBZta2V9PFYekZrQ
fGJgnsFS43sGcFPJGn/KGz1NV3o5RQglH43scJHPHQdBG/1SVqpRMgZcAZRBvJqcGSz58ZvUF+BU
AO8Q0u8p4flGq544+yPoZy4GI0w5RAudnDce2Ay+0tbn6+sdmDUmgkzpQ1hsyrwmcnkWHEZ+rHug
h1TKBAc41mYaTf+Y6xXS/Z49RoBFi37+Qx4hEQdQ8++p1hbEXyEZCEWFU0k48C9myZbQpVUYqdYZ
J7gtpxA8sSMhSq+mOD/NHLO1l5OUh1N/wiBjBATbC6U+yGoe9nh4xFZFVUTXT3KnROSsB1M6Hn9y
Lc8gwphoESBdRXUOpAgFDn7444BIJ1ljMWR0EGreiM8mgAu6r99+6tW/3kwng464c0mdBybgTZhe
qDZfSEupj/ig+SAFYfiFif1hI1nIie9hfqkNCYIsBEJNqRTQ8qWtW84pDI4LtF5zJGLWOjLu9GXR
LC+E0b6rFVlEuFjgqTNZUNVTHuXvoWjCOBW5fsuwwp1TjgperKVw7vPc7wfun83CK2TN//1rb4p/
m3BIfCuyzVJ2PxolFBXW4U5m/1abujat4CexG/b/2Q6QR5uPgCJ41aVZ93WJ7jkwilM3no/ttEoC
RgPdbLx5WotQJRZse4nyc8lZh9StkfEVZTS75UXxlSgeaSni9lgV5FofhYywhjv4U5zhvrJC7LPb
JS8tpHmZiqJNpGnrqGJs5sjFhgWHR5FjR5PpeY0oU/JrKknydw7opGzPaqTQFw5OKLJv5IFg0D7h
A7uWRwVgNXfAv+QuwlD/L7lAAgbGZ/0pvgh08gFzcubq60spZMkcBC4lZ7uKf24a7wv1zjVYAmAX
R3AZZWc9l6B2D19y+vu4I2Y/3mQhegwB0JGV0Oxl2Ydxazu7QtAPBoSugJ292guaumFDQqToZ+iu
qERNNUWvdmoQl+dQWH/ZWNWp4hg20gZf1IgSVxr4E5tuhjLUjCSLykVo2W1mFJiNPKbnooXmPGFt
2rE+CwpVabeLqT1BjJl+tCeubRGUKV6YU2le5KqyZPuQM24XxR2fLzbdCWQLU5Iz+ywT/KaKWROM
hXeVguRDi8hYHkb1CZPOg9qeRXpJmo4JdiZ6ZmphMzMJ1ViBXY7R21YFjp26QeTyjKDANV/1+VeP
Hc70VXrwRkDvJFqIhS9HW2TVeXzdZ6RlKhD8YDrRrOkOQtxJHIeQ2tYTdV7yan8y0CUYBjy/4Toq
+gjMD6ASnkqsQzDKJcjQ30HsbgGIPev+vDtWHKInsd7wSOzhx2byfKTgTJSezf7PzG9sYK44LZsl
mu1XfYwnMraJf89tuqIlUWZG/9ahCVWM93n91BRxEqdrkNG/9uirkHqVUwNu4o8pioJsSQ8PYEmN
mHMuolpnTUsXrxNEFtyEfCfIg2fbtRShNj/r2L2ONbBiVbYfSvSwk2+0aaOzXLHXJ8chYRebZ656
B0c3ztOAZEAvC+xN4NCI306ummbVciWLvWad9mZxtdH0qjz/fYpkoOtc6lJsXShWEHqJOa4ATFPv
MgqgMYsK0P4jBVBghJBtywDXuMiCc9sAlTwkRbxBjFdP3wR35gD8NE0PQAjRa8R3odaMFvr+UYe9
xLuZpl7DEz1Z1DNpHpXV60nTRspcF8nYaiRxr/llUi3glXGsVid9BjOsC5k0XzGKExtGIEb8K0zR
cPnvW8uftdMjRM2VRJHrxgDW1wtTmKvxh7skmpR+7S46VHjkHzvZhaTgT00OztIPjdtF4u9n55AT
15+FvE01+hLdRIRijiMQPhTKyI1AYETnHrv2/npY8a0pjyjNjYhVVC1ozxaHOGUehvq/EdL8S9bS
V8ibcAXJWvqnUJSQ69hZo5R68nGwjx3j9SrsstDYqDzcXfbgdSgFJqgDFwQ2y5w6cEk9U1BTQdmE
mFAMNg2mFI7QH8DhGdytAhfR99O27JtC/5CtWNx9ZIcLaIVw/2qsWMWyju2eBA6BYb3VT4gGt8o0
2jWcI9S7/Cm+pF+hr3wYKRci6Xpb1CP+JvDje6vDp4x5S8W8VkxnEgzVUUQ9Wu39Ds4nSCzBsTV1
SyVWHBdjRXQkUZORD0aoYdlMQiBbGwPacQXeXQ5ExkQo4aP3vWLZrQNxk5u4rHHbeuzCvY4W1Sho
1imvzn8Kg1DFTJD3NoynAwHE10DMAUoOYp5jIUfwcoE53EtUERVqYMnstx0XN8YbGk5VpmFCK78d
egx+thY8z7JWuDqJr1l+85H+imwrNpHhZB/FUhlK2Nccfsf4Klhu4zwNoWPF9batJYyo/ZbWU+CI
OUPbG04FdBo6xN6USVypMl1/PvP7O/8iSI/YyhyC4nOeS6xCzqMX0ywYWoq57Sj5bUWxISh4toHA
g+WrIDM1lC+Y3wu8iHxGoUOPd2QKQ2O9AlTibx+FX8mGthlMreeu3hPBLsOctaDx25u374c86dwL
msHeUt/db8DzvkIB8UGFOA6d+mv9A24sAE+0BTAh7TOdAbYzC6B76f0yJKalfJRJVqL9RMI6y0XE
18tmXoaf9BVc4o8ubCEMBW6Ca4nUwOBghCunFB1PmRlpkMrfDoIpgGn35NlR8CuqhiO79RdeZyRy
dPOsn/+yQ+xHql12RHTiLkLeLtY8e7POB1XwjR789MPyS0yaEn7kB/twwxKHYD/XlJKzyqZi+1C2
7UPRvWP5cJbzrb+HRxOnPmQJGR46iKlOe0+I3mPdU6L+SpldBc7m1Cb4G4WuRMxNq4jrwn3a23jb
tHaOrUsLU2R9ZXktM0gt/kik5y0s88tEMrsO+bFPXc5afLL/IuB6pmLjhmhjk9VqPw5FkDdrxgRM
8gzMCaCiKEQptHEXPLTsPt0udUcvOb77SAPI6uD9nYaSGtxMGKkTQZln9Jpta34mSncoav4wZIHH
uEA0kBtNr+7PAdGM0GsGLgKZ0mKacg658EoD1mZb8oDNvof+0BpVl8anMH4kIKa28SCZnh8RaiS0
AvlBCs6mGxRf6bx3Bo/FiNuhCeQauM1NLhRUMiCdCcr9pon9jQvyoaVeHY6DmJribHGxWEEBWcfD
a6b01LAViFkb44qt2b3cLrzr0jWOWjISbd9TkJ9oGdNFUVP9KwJhupdtFiqqqIazFD79ZmT97QZm
XBuZg9U76b/XsmK8JWYIEHpLdRHvcyfN0iA+vrRkspoJmOnAOSUNl33tFrncn7FJBuCTM+8lO/sR
ji2qcKMVf5j3/ArNug5BICyzY2n1d6xkaAq2FTzvVFyu7TJh8ZsZ9CcFfAJmZ+SMBb8upGoxWE05
MWPllMvRBQ820TCBK0N3oDv6l158QGuVK9eGOoK9KhdIXSGl8TCTjteKIDQy5nEM24X86Jja3Lod
B4teBfOMDTIc9x0+bqUt1snf5RpR97GjJEjzX4UzLtVRzO2M+Sq9ywgsKEVgPWtwNyyovHnwOzgG
aY0oE4Mzc5TVUHjgMWuD1pvGRwSI1Y75unfmCos6PASrjPhd/Sg+6PWTGBxUu3Y3oGwhkoMFhWO4
xeQrtyYoBWdbAhIN5DvZProWn5eOTwhTB+igD9pOEe/kdDai3NAPEPLt3rLx2K4xe6LnJLrQ7OEn
xFGU+CXs/03UaJyVTDFnDG7mJ9RGRKHlJur/YWpxaR/n7WkhzruKpMWek0MzN2YNkBRnZc4FCpCg
KUW29/FOIaEM8KJEejRfsv5kzy1idy/3JC3kRmrv0PI39c/+k8wqYSR7Xn0lVbc8GORx3eikOGtT
8WyC6aliQgKA0eWf0FWpEyW1JuV7IxCwGhNilGofPs+TZMuaE5cVCmDHgFVnwCUGYAAw/ebnDQYZ
GYmHeJQuuRhPjzpGhwJGbUDIEkgu7bS/szVllIE1JQyVcgmwAC0BqFjjbw3Ry+Gwf2Abx7E+rtq/
GyVe1wQ8bRERFfqTJMeYriMMIVCRSeQn3gY5thpOjg5b9hVheLAlR/znU2k4ERJYNR7ky+estNem
0AHTayQlvMVDNvrb0EmJ6oviJvzxf176XRoco6UefTaXgXKLYrXr3SffZetEZnNo5/sQIbLPX/yi
GUytwz4eYV75tqylaa9nR0k9IkVPkkadvRdninQjoiFurHiE8zDHOXCjrN4rvpqW5AocfvIyyGHx
4jivf+hrQrPsdSpuLadQ9z8/hU3JtVhT8lgwwxAsCTIKnkJ79x+tH1MA24Yt1rv7xYvkAokZvk70
1C5v2cNPLhg3XwSg/NIC9rPy4n7Z7E9846/E32eHwyyjUlXC5mkaWvS9NvK1pB9qE4npSruvoBei
zngf6qKgLiOWZC4VKRHeVhzFSecbLetDoH2FL7GUWpRrWCCpt7MXkH8HE6nugX+X3+wez/jroJJe
6IJTDos0NcDCVaihVQxzvmugDbtmMIQ9jAej7ifnf/7PZkOsn4RUGrCYjgCe3sKHngsp4KrMaw6T
FrfIta2y8toxDWmuQZTNs3nDeE8O0rbbPXm8/iJmysQ2OJ+2mhejlbBTCMjSGOIVhO/78wCSp48u
9fQo5jWfmYrA24n6jXgZ64FnMGkg80BsbIfkyR6kJuM0JH5WjAJVDWxM+/y+hgOWnFoedasEfWm2
ltGuiY5baFQZqBzloJXqeKYVklDuaB4rftc2Ql0UG/uRqVAGbSBtnI9qGf/6maz9xy7Tzp2ByZ1F
wjItZQoMQE0thvzu/m0Jw1PotfSBupteqPoo7i/hpjuDH2wvrErxDtk+992b+rFxjmaJgUkp2S+d
ozk7brwJD4iUzqYrIF3WIvOTP88rX/Cd7XrH0cpPjEn6wjwnDAgLJaxUSxYJ/ERtfA8Cep0b1Iox
XQVEcc4kPB/qhnjLl3GwYLVdzrGOkCbX1WfSDB/LinWaURY+AgzV32lMvtQhEYZyqo9HJ9g8n4hl
o3hR/WelN7d5tKxuOq6fXmzAhQ6tuun16aBlUBE84WcnxNojpVfY9yktk4aaTFiokgUxseAzMlb8
BZggmTwYPrGEXVrYivlVAugzDaO+/e/Fij/67pIYBsS31VZEqozAv3F5BHofMe+kCrmBb6nEvR+j
FXm2t0TL8OWswRwR6Y6SAS7YhLde9ZyY7sO2nieImbSbKBjKWwJ5WY66f3Dlob99DSfpS9wAhA51
cVQhaQ2Y4mn8jyVPLruqR3rL0GIWU5vokQkmug7s06LZ/FjbhpDPZRh63eys00KNbg8bN3dLct48
HD8dR+qaaUpBOAR2+dzNW7RTzlUdg8koCzhM8WfIbKYluLf4dKJ3ltTcIXAU4z7r+dC8BL+ySf0z
FcPRdDah5FaeAvXGF+fD3DXdnrU7WuLsSF1e5voW4vuN1/35byjN0sAEDCV2U0VZ+JtNnFMOcU9o
8W5FAvLRrXaM/OFMTOp5Abs46TItpk6TsKSfs9KLHNcvh2fRj1TWLw0lQNh2FKqJ8yx+Z0EYRrUU
+l7GYRN9VZ8jNT7uxTIjKbtfPUyHSW0avMF14dOVRYKj7uvzKt29L2aT470PwX40tx++lfwUC52P
qoPgwFXBWMgH77xa4OKei4WeWiBgwOgkTyQVMTqQbSpl/ViloGyS60rXeN5HOxdpvg0MaM0aDhjc
2Uo0h7Z5slPqVmaGN6avuILzIuWRzaoQls8i9OgoSHt+AjvMNDbHts2p6lcn4cMHkW767gVvjcsu
NvRKr9wjyffsbHEYWdrAnEXTjlcZmSWniN25P6ABMyqXTLOfvohmT2WdX8kS4z3sWgJ1/+Hm43qe
z+qM56/BHfJ1kNgi3DCWzYJgDXhDa9PrTqkPwrcVvo4eCF2K8/jAfJWJiSL37QRxtXvnMgEuaWJ1
jhMaLT2nANr7qWT4dqdzQatwCEHxkhZ8EbHN0ITP+1XG0o7MlS7qRUgm7WQIKdm/raKvgtOd3nlK
lEGJfWc6S0gxL4bCtDYwCKJwTr+F3roA0qfjwIHjn9+/vheBNL1M8WNc5/qeNp9z5I6T6596QRSQ
5zZPLGw8Rmb3uwi1vTXRbCb5QM0J+3IzDPEbRmc3fJ1BfNHmy4aU/bAi++vL47cBvPGvUDTmf3C3
oDfDaumSkalK53aCYANneISPr1boK3KBb2wVwvKvhnsc65cxWGnx8LFGHGEZgRUhr8o4RQ7lG9Kt
UVNgZUrgIPt1WQ9whej5rO4GM+3bEZ/uSdydZQY+kxfEH0IIliM/TyIn0QqVbzmbbblEpSqf07Rl
7KYwyyZhVSiy+TQarq4LMAJzgIZP7HKALrGUcaMBtGCl4j8DVGmVHc52MHnpqXKfSxr5IZ9ONYPJ
2CjBO423CHu0dBmesEw3r1tCMK0ACCxxLwmoSBkRZX9TLnicllDnKu9SnMv/WHBSnEGuUezjRNqG
9QE6NcVRgTMbVVWyzrxfCJQSNGbvaRAcvR3LPbqy+9tzjfKJwM3MNSJWyg/iwBxFd83r23uuhKq9
N+9F5682yG05Ql2RMCqQ5TbkwmAD/4TPBiipo9nma4b1dXWeHy3DiwjbCmZIaKaTO+VkMdMheyUs
Bm0tCpw6qaUZhXSDSnc4I/kVSo29s23kJItWOtrXw8ji0vB6OVnSkCBqYiFc6hyyLoJ3G7zjGh+t
TkNi2XgsKHWjlUHkCkYTBUpsyk3dLa2JHAmOGy87baj6PePq2PoQvmgRXrPrUGPWFRIAac8ZeTx/
9tYnVHfpFobGsbJvkU8SnR+OFgIvNPvOga5KooDwiQ6u6t9hHfd2gw+5dRg8wVMev8EJTmXjE98K
4IHJbUWb8qQSfBJIf2ob8czYxIPKPCbLlth5su0BPPPvaAZd9vKEAoenY0/OTnoW/BVLVAhWsidX
c9OHwnPfqbQah5oLgewuJXe1YxbNh53gJOC5cc1BAEqwUTHQe4RhsOdDD1kvnc1NngLWIzTyu47Y
GzzdS+z1sXE6NSg1aSM/sITSWy/hCiOY+OD5OMufj1Dj8O8eBNup/nl86m7yUw0m3GkcU0lUEGbm
BrAR57WvKcEB8FwkmZNUp8h1/4obdlQBsf9YRcLJ6tb9e7uaPlsg9nllQQnXifNfo8W8BgcjwAqe
sxF6GMVx6wb3gpRC+XVeG7bDiWbIUm2WMxXHeMauGrYsjUIWcb3ziI1gfX6c04qbtvJGIEwsvM2c
R8W3OX5za0UPmH3M0tzq81IHwYgKih1Hh4Ei31V92zJP5lOyQk1BbRYgpsTIjhSPOk+xhVE/Tq0e
mvpaFFfxkCs2ckW3GVpB9iVMFiz+AoHSkVFI4aKvbNXcaEE/QQe5iyHkGIvAl9tNTrD4lpe+3jZC
6NYMAbe9HzhFydoKoKpHZxWyGMNApEZ6g+xMkFxBaT3HRRGRYtH4iF+HGC710KnL6F5AgE0Y5HBR
0mPCmRK6vchwJDFrJMQEeicxgE1yuiPuKg5N2ucKa/Ck4UfGSs59pMBbPahkSIrHMCcLR9E14sgT
rEMTINVHOirrQHUJnc4Q6JsD/07Fp/SCewom8TO6q3nBq7uh64lW5TDBbgZoKej89kCD+LE4pwkC
R1+zNIjwF0JdLk3LBVYdWPpOj+Nzl2s6ALKJ2sNnCp6iVTTSgX8HcjJpRD3hEPYIwIG/NfesKQLm
W/HsurL68Sc9U09eYhh7UXJFOkd9QzQsnFFHylaQ9ioLX/MlGXh7S4MK1XDnT+U+Y8Rxm3WzmcUu
e21TlDNEhA0700QXJQ6FmE8oDZQGXp4hNk0i0s/3h6q4sJc6ovD5IO8qUlWLNaz8ETBgeLTEgW7f
Mk16PTks1PG8f2R9YvGysjWHlgE9Z4uXevQfrDO5wg2r1yJ94eOApn7+czf7rCbtSB8Zo3Oqg2EC
STb8rsLUuKvB10P6zeEcphJ2m78jJ5CwpqpK6tbpohJocwSGPg4dXNAPidKj50GjdYutkRZ+3/5R
RrDqLt/iDZwG8pAoHNBMXDEVXmu5FkRuUY9hmGazMHdQT7A5K3A3PqJdsw6IOr7OeBo/5OgYan/c
FUW2RJ7I5cOHQuOR023Dd4fsM5xF2rs43jPZjZ+cRX3IpyWK9kF2GsvYfh0VTBIJzXHL50oiAPCv
0trBWnLI2wlLtPQqhl5eaU40n2AGHgK7lUuz+x9hGjIIb7zQgsMJXsoG8Ve//8TNlcWEhu3Gl1MH
l9WrqLDNPBNcpFmqL32OQp28HdkwSVPhzeV0wsX5xxBrRtn5wgPudGXTWTg3b+igYpozfjpsJeqC
CdomBNHpJw0rXkZNASafRPksfAdQVzjAONTHChdEdhHzqD5jjBAG/DXBhOPyJsHp/dQ4P7rubrnW
svdKpe+YnkBtS6MCxNAZvHUabJOGY8Hx/ZJjUY9AQl069jGVu38lK/rxS8VZJ97xwx8zRGMHrzsJ
SY+uVmtu6xhSl+dj6sEgQsUJHXGCJ1oHJLycSEJ4bj8swqG1DAExxa0W1mKih1RVy54EmByJWlIV
a1RiBg3g1IiswTEls5EhOrg/YWR+hJfyUxvCt1VjmGrsyowfXLO1lVXJSfnyB9xZUGrwPq6lW8/2
q+ZSV7FT7xzt6Qw25fvnUIkZmVMWpn6inww4tPvJaZeIp6Tj8AoI5Zlb8KT/liAcu90RQ4Lhk/Q0
76vl8HT0JHMdbEbIUM+QEP8xcGznseE8K6YvKSJ20RzDDSoRoCZsaJtGfPWh5scEWgNXDU9Mf5kI
Wtr+TjmBblk3iGz69DF64RB0BxjyTpd46BRhWfarHbN+J5QJSgiDrgxkRKHSHKZB2do7FF//A46/
lREQgKHfK6rxkLDZVB1JEY8wlOKZDybsy8pD5B9kUxmcm3O++Di+MbE+UzP8u6lmaescKfmNi1eg
8v0MfsQLOvPwPANv5k5d20yNJjUGiqoTeD1O9TtIWemhjK+sUpy+4ihSCu/Rz8OJZ6r+sZu/gu+M
lOHdik72yaR0naMJSH7K9774nkEbmOrnzDPl+/H+wSl4ydmWRZ0L+lBHEKhNrcyU1x2sgNHsmHC8
8TZjPUlrbUAPOU/tFIPw5oJvCdpZgeqY5u3VDFAJjqB86LGYvRhgQ5tj64iHUD54Uatim60179qc
Y9mo7vZpX6FhPAsn2h4sI1qbbkgNPiFjyufZe36Zb5JdFJE6IBvuvkl+KPSd7yz8At7LZqD8YAoW
J2B3q9NtZZ6D8M2gix2VJKhetPmVsT0joBBNvVDnh2d5VfbRV/JoYyYe+hzNfzsfdGH+ZDBTBmmE
cEo0dmBXpH7x49vUVwyXo9CS0BbmaBsBZncRJzWfrlRjYJQ4fLr/GN3rJKXUVYes8UtsAF+Y4YO9
GwlSOV9ti16f6b8rALsFBRzXK3dTLMeinQJjIVgjQ3+sv+yuBs6TjNbzgwhxtJuoIAWowX/e6ncj
Zln/iZ51oWxGTheT8QFRKAx1kzNNCmDitA67SqSB/9XLKRDw+38Dgp4mhTL9Hbna6eE6+My/acQu
sSmc2+1Nk0ME+TQdlDNmnO+nvX7ZIchuEOPEiDhNIXW2DNY5M7J74bU8RNyZLMGv6MI7RRw3CLbd
qD0ShwxdiQWZz7iB5Gpk+INv5/3ho9xeo4sdqK7Cm5jWOstOtPBZAirkWeLIgVOE2wzvVGHfGEIl
u3uYwfl9BJOpLbkX+uXXo1F0ZUsIH27Y8/cblZ9g/sawKNfLCsgNmW/qMNq/w28e/toC4uhnsh69
D6CddHtKxmxE1aM/kCheiTGP/KIT8ajwSyeeDk7z61NtlDHMsWvLaQNPuLlbUsD23EDgokO01mtF
gBYaMOMVSvys4LT9tw1wUVFQDrEuFjJ9G7mvoRxmLWFSmKiu0xepwjcYstoA5IbJfLERXn1goEpF
h474TF069dMt0oaxVYOicgZPwxdZUltrVz9sEFnzZr3YYeq+KmE/ais6DqOlxYh7kzeMyPVA3QWM
tjDO70KMLxorCqydyhxRE+DWNHkE/9N8JO9jlWk6k3vDeN6SZvw5QaX8ABvL4sRY93qEnngZTdJf
Fx/5JkYGIo1PGZO/RgvtZ159Eu/kD0tPH6MJ4REWfaf1uaTDUySNbGAtfVmBLKTUawWiLy/MNBuI
8OicMxZuV8AQttAF2Q3Ena7i1pv+t+YHI62ElUjBIoQuiBAgLeP2dW3qg4B+INyuEX/ScVZeGNEr
5OPyMaos4+A5upsgqgy/SkEb3uWA/ip/DH9gGm/yLji0YHrIlj1FY25aWxG4hY6cmVNg5PYIiVv6
wjbPnEjwgKC+CqD/GeGtiqELKqPSSOEgoIPD9b7JYWw52QKI8BrxD1otGqWOqwqvMYqtu/yw3lua
c4XOwd+s3jbmQRJLuo1iwpgPTmqxZsgvRPZXcMP6mS89cXhFP3EBGFqhjeiVkdX8GDU23zCyZPci
E15DoWTkKo6ZwNBWakK9l6oS8T3V4eUCU2GILZBlUqRHonCwxHDUiYBN9c/clgO3Yb18n2/2AK35
H7mpg3CU5Wku6RQdPW1TbEuiJqaf41huamubTQlU9xZczUWXGB0+SH2C9/EqMwa0N36X3TFydMwd
Bi02SZPNyDvvHsfmFyGbCkspdps/rWZCu8zeJEJMfnaC1+t60qMryok5uv7IpnqNKN6ae5gqwbk7
i8WWpOFXZUl7s/hTwQmwQ8VeCV1C5S85wP+7hMiXR067fcH6AmO8PlP7IiMR29lTjQHnMh9SLqt6
GbWm/3pdB/MOiW6IqsSq/aOuP2d7EuG9wwdVgNsEAY3swPeKR3ILNdsW3IhLTkKdexEmBVs1jdpt
QFqy+KZanluPuJ+dzZR0x2tNVkWX7sorJLNWdS0D7Zko5krFSxiSMv1atE897hHG0LDkZyYGxX3v
UOLFHGecAjAR4t8xN6EHhwWE6ArxNQh4szr6KcoHpAIjSMoAA8V4msyhXcJV+UplEXWa9S4aSDVp
/uHHk2+PvR2L6olWK9wQbb5EdHcAeZc6092DQsN82AEvY56fxOT6CB9zO3QDZb3Ad9WdxRqBVCZM
Sjotr2/r+oygbryIAJpIIDrRahqpS1ChGxrfYWUP3MxxyKOsmf4+x44dNQauRuuQYIy50mBSUM24
AEnuqMxPaMlsOPRJupxk/rHBe5RBflCiFyMRtkLq3LXKESTGXAYxSrz+CzGc9kDRmKRjNfmxwol1
tlGJ1t4DGFI/FCppfW/zsRs5D/OT4STVPdI4H2kL++GNHUqr3DDkc9VcU9ZqnTfDlNSshuSJkB3H
ZN8EXmEL7cDrOL99emHPEGdeowS8VjYTs/KJkhrA5+M3ejfPJOAu0Vgjuett31JsSGNN1hIkWX6Y
Jnxl5uOccWZ278subc4Tw+MtMABPEWYZlBWlhIzGSFXi3znXneU6/OMgZflrUNRHe4Tl9tZ2HX4J
tt/t7eTqxueWJOM9sjnEnK1f5G3kdc3REfvoVCzMSr6HZGnvdZafazA88fFuX/mJrHwU5rH9YFa/
YnbfRPOHwqliHAT8c/ZLxaMAihr48HbcWKtrE+7gEZ6zFoVmREUK8SjQ5pCgC2jyS6ZzWfjmN/dM
c0/6HzyNqnYJp3xSFr7lCbR/bM/QFWzvkyxxoJwG0iodBlVVxBLqCdJKlGJRb5JDzwUpfdPtJA7I
i3L3yTm2Z4Ab/04EFWc0TjE08XpIC4iIMki2uQ/PsweJIG+FOrMXGqHV4pYuJ3mcc3SGX1SKNMog
xdLlKhktpFZfe2Yv/eMlSmZV7rIG3ajTD5c2B8AtHz6H+qX/VgyfClX2x4y+wvLTf3SQ+tlwmz7H
fvZ5qzLNVpRh5qmaShHJa1wxrJdSqMQxbimBtWriSw4dv75BlFXFCWjPhWa0vLjy081jF5dJYDAv
b/cR04nGWkQ5O8R54e5ysBsoZXBE9ysKga5f0HK90HhRqViv411DiKOaTlAI9OX7J8jHLjUN6zLk
laBseHtGQ0tIvu7gw5NEEtuhZRya9jb/GfzQpQOpMsNdw57Gp3z2MySeViEBCKeUDx+N59HYumcF
ZCHc0iJzDH6iz63xT6QMhvy7HCJCkWbpUhYqj3WMyh0KcO9Ca0jaaity3neZC5PU19JMIEIMxiwB
WM2Bex6nJpBNQ48PFkYol+YaZh31K3xcYHzu7jiZqReCwfTD6VXDJmFr0wIChBe8F/3lbdTB6a3l
Fm4eJ70RGCWFitRqW4Ynq2kpYG0eWSpO/Ye3TEqCGY6G0/YzpPSP0O4A4quP9WFA5uSYD6AeRCk4
nZ8owmMtNAWT8hdLfPwETa8GrSBryZMF+RxjrJaoYTFxkq2m6y1Lef/QSK1bWlXofh3YyJPz2qWX
fRfAZd7CC/l4PlcZnCEjLe1M6yI6OUstXnRcFjdvzHyn31udN2CyHf5BhpXAnDtEAqQ/whNBaFeW
RJIQTROissfzY0bWMuP58LmKDqyvtVi0olGg6kqAsT4+bQx3U3xYbmfA0aQYZGLjuwTW7o9f0SNV
7+DaW8GGffZ7uLILtga/WtPbBICt7+V93YAjZRY8UepXJye4sEaFwqB3jVwfYtpzhcJJ2f8sqJ8X
G0kXC+nd02XCjZTuMqhldRV0oqhHtYezj0lqKmNb6GhQXF5P+tWy1bzXi6MHTH9KwMTarjCqXVzc
66tn/kpXA9yX2bZOXfmSWU0gJALPYr171GyFyoK6BTFkT+Zs/TuQc8O7JFkOtBMNiFQpMJxqkudD
HeCZjypCzpWVXbEwqsygv2ow9xQ1kE5jkaHf9B6dtweKE1XU8Jile3U5WBTumxuyspV6f38ed+N2
IwOZyPb14iqR8CZxZkNOyfVqtdhBdcMlMdDTVwCROwN9poIf29kgud3oKQ9NUvRxX9agfgDJ6rOH
75VJxOzE1tvWGePf78x6lWL3XxdW6JtM52Kc5sNeeb33SIdebZP4xLUhJrgN57WaUtBfkbyUU//g
9RLVFOPubvyj/5SXQPIdYhxg9jPSPLgvSBJAKic5hUMFECCb79jZiOyKcBAm/n5uum19NJ5eFQYr
biquiEv+REGWJ0ytriKMB0lD7QejsTDY7hDmaGuRqyl423NOfHA8Rd1+hh+N8ySfo6oJLdpTUwOB
JU1eZ0QXSJQothP5p+DzJ19BDEEWjs8dRZr+7dWwVaeHQ5OKELFISCOs1Mxdbpm9yPz5n2ANiqqo
16TU1hegeO8Cy10msI6XirK3bscIbdF39ysBUK7ZOQIiMlR2vBGPY+UK5706W3h8FaT90UmM7ryv
9bDIIoQYee6sOR15mvzcZvNYgBXKacWR32yzE4o0YwD/z5cSP2v8TC8RScTbMx+Wr6OrVklRD1zA
mEFQHSsY5DbeR94XbR0CpYr5e8F/QBroYAdH+FTdfWoTZhxu1wJ4J3MNSwNXCQ8wQBCRBtwqpDCm
2jZXO6c9+juQ5yFySdGmye78+s0JbZcQTViSyu7Ccy1b0YdPbyx3XRYXNVDtFX8vTLC3OTR0jduR
e6WY/dwsIchS+WLAR1vGYHdRkZF62/LJSxJQNkeoj9qa3PXzWVjvLb+wOCx0sKqvLl870bFrNB+N
RZt654C0Q6go1f2y6p2OwqlrU56mkb3zpf5erBeJHg1Ah8HNZQjnKUc9mZsQqYscJW/8SrG68RTY
QVTaaXnMZ8DNfsgbm6ZLyHxMXcEt5lOd9UBTanE5y0i7AzRoaz/gk22meWV3Z1YSeCsFDJNT8x0s
7W/OtR9X8y9P5J9U6eUVkpuGPzkgKmW/1G4USab3vwZnCSUQooztkd5299i0iCHoAZbVSDqEj5aC
UIRUD9yZgiIpWcvfWQGLs4qxjw4yKMIvc/B+sFkNZFbYmNojOlU5rqufzBEYciIYFslvLMu5fXiV
zu7XHqcmMle38YAuo5B4FMsrI835/03jQzCWjdw42rWMDCVkpIoJAUnJKyvUY/mMvRQ9SEU8iIr5
qyo8mfYhG8Ffy849aLMGV8gJ0E0odK9WNHGsCM2fngB0uzj519QR1j4DRp5NivDNBXoacspT451q
Znnd/TgxyG9R6MxRakuakPTSoR3B/O3B2V+otRZ25UlRftkT8BtgLsMjIeaUib8MdsUVyZylnqA6
EUBW9TbysaB+J5zuRey/S3V3DVhHu8SocALrjjKaYwOJQ/WaNnazdWUML4zQNnWc9QSQJ47lWx3F
q6a1P7SnW9CakpSPYpO3zq0hprAynVQrAl8X3VavXJMPRV563GET987uOzvzPLBenr+mORrl9tKZ
2//cnyFj70eghQFIgJlBGxzT/QdgeQkgkgGW1mzkp1T7SrWb6FZrP/gKy6fOhB/fafUCVH1SZNTJ
hHrn/VhPrwr/+ezkvDLD9tcaJtrarWfXs5fQdMO4LVGFy/V187QNBe3cRYKbhZGLwapqSvPyT7I7
z4xZ5gUv+zFZhLbOKxWeIBZHm2IY8uun7MQLeQ6V/7v59q5g8CtSDAdEdwL3qm+aDpRA+bnsAnKG
7TNl74NcVvM5AaTSOgRkHPZZUfqWOzsLkdoPfDZWs5V7xIgv5TIil3ymSuhb1Ejkfcm34f+vLG7S
rTY034mc0IJTefkRpl3cyvAYwwk6oEpDtTYkvLW4JXBQM8QdvTyitbw+rI6ZCfX+Hk3tiuJBYD/+
wejYvdc4MtNX7nEfgsPCZ9V5qma4NJi6oA9kWtePGF+olfeiAtXjbnWU3G7sCyxjsrc9FKHexU9T
42o6/9aPUJwkQhZg0O/jH0ba4Nxdl6KEI+A9d0qj1O+oHfwm+Ioaw9OCUWTJrk5ASba5Z7SbzQwH
Bl7JVxoCBJoNZjP4z9iYU6AmdZ1Hpw2KKvEvWy4l/FpJdgzedHWHA0/h0ZG7Zdn7aeHgc0ce0uL+
wb3yNBrZ9LagXbUe/JtNBjIC9pHqYmUNcxDCpwePRCqo6Nq+6HOpNp6Honpdduie7rFpTMaBMfVa
X866o6AX6F3tJAqHapebY1dAmsRN9f8D91GK3Qd+scxhVhCEo9exXz4r+2MGR7m9qAIlMdIxs7bI
8nyYoXXjCviRwlHwwekdTcj98wh5IH95EpuIJbeSZE1WqgF33SqtEm9kCp+tqxUhw0fvJkX/cdRb
Z63XnFgJ4rHLI4sIFWWRx/gRKWZv99qTednbKFRhaG5wp4S4vrSMPmtSnEbYC6fF7LqqTw7TBCov
IGiiusKVck+Q7Sr3SCBhUaRK0ZLi2ST4QYZ6ebobhsKAdCpsPhz5HzF29Op4i9bcBWqfhF9MSfRU
XXlVArxOakNicORDFm7fItagBHC40ZIIbgQstZZAUlB7ZY3S+hkXJw1obxUmM/Z2nn+PcGo5fq9a
qTX7iSKbvuXlN8ZCUknEQgKbTm/0MIGxADcKTVV9gdH9ziuJe9gcerBx7093spT7qeE+fEvnQYIh
ttnSKapoSjPMDCqpvNc64fD5B7hsSVpWYDvsV/0KCoL6F4zOuWONjqLLvbLdZ//J3yN+RVq3PkCo
LpFG7KNTxl8ppK4g24PDzOyZI+aD17ZWI7R7Mxmpu2npj9r1BgQeSGoAaedB7AL8mJ6yvuIItpm8
3CO7CQpLQ4OulkSMhfE0cDO642OrPHZZsyM3godYK8iSkA0Zq6mAYqBeUjvZTvFdp7cNj3AE7xJq
IaIZ7YPv62+J8ddkjD0CqftEqumaINMlbIpIXvKQFrh9ayT+FBKJ/RLGcWXE5sTCkPhQGmawkqkH
M8PR6PUMIu/YyGioPHQvGy5RBUGYgIb8+Rdnr+ctXXp4Pg1QQYIpvubiPlG4ihnT7lr+SkKeeWhp
wcp8cDpPdZOeGK1OlU4/sn1qmtI4pJSAKiNJcboHKqPXgmJQyepJwyAgq8QE/D31XUj6vqrsaC0G
uTqZsU60SPG0UXmSn+HqXqbLMMRkRIIAjixaYdQkeGbWXoSfEOHDmAY5kN8o+FD0eOrWmTPr7dn4
v+pIjU+LSiYgxL24S0romCme186S6qjceVrXAhIi3ejSGRRoTFklq5lf8zueFx3pXesnIkAx1n1X
Jd61OeQX6YCJGDmQWhOMzzPvQjVSwa+XHVUWUiT/oQ4fJCk3V+TSqxDHS1oGopE0xzDXUFjqkWtA
fcDVXRQNIVJgYcnmFO2xtSA8JCCZrkaBle8LBXPCDyPmfZh03uRyw3P0mzqU1rSMVhgKu+gBTW8d
JY6zDRxQ27FrCpbYy5YpjkNODqQ2Ojp7h6olN/RtYdRSte3BSrHNDSi7kI/iC8zC3HdpsRt6h9Ia
UEBCOAZGTRPckAwfSsz02kp5JaaJrMH5e2urlc4H1ReHk7ORv2HbErkaYlyXDodp2FcC/tVQjjNa
J7+8haTVpl/R0EDOrTayWBs7ORS2N0FBjLukzcEXfjlbpCd3/1g/gOaCLUWLP6chTKSHgjP3a8du
H89EPVya/hs4zjFa7BgAY9qabeQ++JS1zSKm3Bz5C2oNBnGIk9v5yQJRr9DIYzPFdzXnVxjqEv79
M6KRkaxFm9joXa9aCh/NzQ36xzkx2jHXh32bvVDoxCwJCSOawb4XzW931ihN2idveVJEpkwRQEVG
OmMARI9bB5Lza0TW6hoCxY+Fy+mf/XfHGj7s1cbnxD1hFwf5Lsm9/h0SEOk+QxKo7cZx5C06uFcC
JPevwVqvUGkKg9lzk7diVdnKv8jGMWEREzwwiReau957L8byD4yp7Vhlb4aajQiX2RYMsGYigRC8
7vnoUTDCj6YOwSyH4YQ1Gk72PrJ1d0DtECuo/wZNVfeV6LL9vKElMWs3bcvZKQUIvg+TJRxMxNM1
xOZKg6n4xL2OynCABaClmd29XbgcxVf0hgYAdUQrORU6fz8c9qUndV+T1cFPgwIvQdZ9ocQEBk/x
IobKxVTh4xj+CHK6JKPwNbrQB2GStvmsvyOtlkV+xT546bp6wxsylQl/5By7XQ75NIwBHOUhupyU
41ECURAchLP73cTrtcuPHjC1y+ofoK8h1PuRYHgD1UNZPwjQwUtvjVIhAP27hVaeQTf/SS/xY+AK
E8rCfpXrBsaTzv2kDwbzhouAF8sKZ+rcWaU4qXvCLHYbGZK43k/r2BBG4nfSTe3Ri66zEts+pPLB
dBa79bi0/VSqhcyB5yOIEcdOzTTsMvhdTMKMv8pZSpswcPmlFp/Xg4hxKumI1Q/LPxqOGbNOxlhZ
Af+4ghws58QDF6qMhiJO2SgraL37mwQbz+LBfvYXnS4ShGBOf0O3tJt9WFiC0y2yR14nMMmFvKzE
0C25ylsIHTAGRGgPpk0OVIeJ1C8MnKCKbqmtaHpYtAKZqr7lwxqCjooAGQEXOQhRyB46Lwnlpd3g
I1WHmZGsORw74fIBjFHvWUXtoOo8xh88+E/w+kAHJrRe2TqiXEBzzoS2m5JDfQkRLkUJXcntvIPE
p94HPuj0+IG/dJLOJ5mkm9c4iag8I/NfJ88wl31Xji7s7H2wQkHOps186dUeqinL+XYfVtiKeTXu
1cUKkTREZ8nJ8yG/rPjPfzURj0o9KLSQetLnGCw628bCFbu651ti9RnGc+VyYR/y1UxXFmojjV8M
EM0NKD9+qkD2R/HZ+PBlIMAIzDrQhJUlHNnaTCgYaSQJDz5uLfjrnxWjWwSVRHzp3oUudhSVoF4g
e9Ohs/qvsgDposuEgqjFDe2xsCGjMKhCbavvUlYHrpz+rHTzNhsO2t+m9wTvIOsPtN91YF7elfw8
iYlv+Q3Cq8HhU+6Z7jZfFEQsMi+q5NVFLB0vmg3WVoDiuSRZmByPqy7bB3uLQtgwfEuiIeNEmUkF
ot7rKc/2tutkHXLYXMgNnMF8607hw6QoCiwJb5Sr02dpL36taUFdcl/gkqF5XpYC5OeHCF+Api2y
N5if8arRy5Rrsv5yTkP0Xp7I1oYVXJ++/w/GKAfRrjvQ4BDGgawtXCfDveMGyXGjnZ8l0d4hiQxW
53eFA87DucLEb/zL+BSQ7YJGMCZnrWa5vNmNQ2QXQM0pJ7AmKDBhgjrtttDycbv0hcnOYrR5x5ZA
l9ljNmGirPJkcY2+hDXDGtGzI+Anl1RDxNUiFVMAS9wuaJnWNuU2wscQ5Y21DbOlZpPpJWWWjHHd
dnW2NyKFV3vYlegEHj9y19QFC3sIEdMzRyBy4w1pRzevLE1L9Xut0qvYJbw2Ldb3ILqt1v7gqKka
m4mCM8VgviVnT10nOOxEYNIKmMqGynI4GLsrDP4GxGfktQLZ5Ablkz0nkUX+S9bG1niAlsNY9hQz
u1sNFZUxDmnXKkwDQduZb3TnjdQBIuUlyAy823NKDc0bhPAOqol3kE6gnRJkpB9UIE+TX/DsTmtY
FBDKEGHFJ8hPHZ3EVwkzfFLLdItlvNl5VHpylyGTdZsxlHq57JpIdb2+xrld3Zrfl6wfJ8GHZA9g
sDYGlunhCAN22pB/Nofoxhco2pm5fv4zH5KFx/TvQ8soDldWn/5ely3kprLni2uTwnXrXUFSyWIi
yFCjNrR26S4Z7SmO/6LI6/Aw9bYVwrChuajlhsdmy6HTNbSrgVf/nl48QQBUmpmryVh4etKutF4w
j8nIthAyHK2JciiKU9a6fZTnVAFMRncYZl3FdaHmdBmmlVKzFLY/Rpl2MBO5aQAhOs+bwbldgocp
Yb0UNuge+DQQEhkOMVxaRaOEUM3wOBzwqAFUzCDkGPMtnseOdO/X2VvpX5C7kEVz3Y3WZI6KlSyg
425pHWLZeNn6da0pfh5D/KrgH1095ReQGGxTj+XNDkDT1KRdPZ753LquP0czrTuWBgsLCNoX2aS6
OxXDzHbzfs4AMgK0hY1ylv41PIwU6lsS/nwEttJSfUCMsxkdb9RwKizaEBnetv7nQj1Ecp5tUW9Z
7RADKy4pJGZ+KFjOyX/tHPRN61N41uaa/K/gxBv6X6q2+9H7mT0SqCrAJWo4SVgsvwxR7tZJNJOu
RwcUzRcg7g4IJ8fIPKJPxrKe7X5C0C+fAVGpvSu0PnzyuJR0vJqnTN/kVA/7NfiiwJntnCCnKmn5
RVL4cRZt1ot+x+COR5L+74lhm46U7wtqe8Wyfx1VXn4S4nDgiB+mVtHl8TKK2aNUtW6Sgn8OkftF
sXklDqNP7X9e21k0PPmLVRCoJdt5T11S14FxR+6n/Mh2HOlHwEu8+NQq0DkhCWRBHamAbtPx645s
57v43pmv9ahQtO0m3HgnhfCZn6e6qs/NkVkQY4dX8vfo9A4UuL8lkAtHZ4i29cxZ3d6w2TAfUucb
UdD4ILJF+aK2+ME4dtMb3/bigESkOFfZGgXmD2Q4EISz/Pa9NzQW0QJ0nGeITW7rxqUeZSneQo39
iAW7NVQnlTZA0c7iirMA2HIwg3IaGWfztPVAj3scT3geSWZ7n6FojDUgX2IMBWLjSXgOtjuspHml
cwy+ZqM+10FCKxwtib7xezXxX5YxhW2da8y2z7h5oI37Thwj9M2vp3kcbfsICg6uXGHkE1ME1VBl
cb5QWwwRjFd4GFZKmsqfttdT0WI6TCw+UA4R5v83wnLSuG9Uctq7m/z1fk/1oPmtzgf5YCkezXdg
fVn6LEYOmIHM8b3O82EpIm4kJPmgP5N43+oSBgCAZWbBxC4rkv/DadSHdTUZ8KyU7dvF7I7fRrNK
xzv0j5Xyedc8GfUNY7d6KBYPFYQHk1NNayQHGWA1ws8tZmqtK5rZBoUosDEAZ3+2wVSuJKrFO/M+
j17kQrZgO2O2csEWKqb6Cp95dY7HS0ZVWQ13h0nnop5qILljg6PfVLOOGVOvfYcTxQZbbxMh222t
2Oznovh6vEKBjOMtreC+oOrL+Ovdl5weGtgA+8LaPeGhGQrjj3XxBUFdB0CyxXVt9C5M4qKqGawF
zrI9q7W5eLbwxUp8vRdCmd7OVmMpuVFNxcPbAuRT5h1rPUSK4KnbB8vopEGTgXTZaSXrYPh4K078
MPaNRkDUscV1KwJcHZTfUrTYttzHWkXQduaMT8Q3b5t/9Po8dWfseYRTA8YWnN3N6H99wlUw8hUb
TFpH+t8pqYw/hQY74/RRIV/QrzLLcrauCGP/JgSxt88/RaSNx3Y7hA15wLU7PeslodrBu4Ub2Z5J
3VhTGvp4y1gKj4UW4BQPNaUP/hJZv6RJ79Y4mlpU3ZT0GJTm+nLTFRFfYZIBcZjC052pgd8wGeHE
/yVoVuI/ysw9WpzbYH7wEGUknweivgeYEGbIcLDgUAswY2BaxA6m7Eap6fjIhkIeLfdDWQapLR8W
pu7RY293aivDxwzzOO3FxUxbH09deOrBiC/j3YVgg9LIwTtOVlBlIXDyGvicuj6sioR0VgHV3+Vs
GkHOhsupZBS3UDyJQxbRPoUL72eTmu0LElphEQUUjTuL19+qsvNwj7XUe30xvbuL6SgOrz8JLiDY
hGZ2NMjHcvLALXmGYEr3G2D7+rJ4f8FuWxxq9aED694H9W6bZ5c3nnFkdaArT706vWEc8WEfn/Qr
jaIMWfIhdQ8e68MX+Q6zbhBb80SP7TC5nnPkkIFoCBoFiSB0EH57fdm3PBmf8Wh5K656bfkYMJ52
hbXWnReLFGpd02Mem5fpF0L4r+elEYQnu8cCoOfIgZNLGWlEg0U51R2DWGEOIRSra6FE0BBa1go7
Qaxr8BVTTCxbblQEnCEdw6rLsDSpXsfKk5/H3cZtYbs/gUjlAt4w+pTQ9GvAD7zsYpL4XB2XuIUE
iGuIkSxQu0ljEl6MTSVLztpd6b1jDaUlJEX8KX6wGWbigWYWlm0ZYlrqNpAVw8NqL/pa8ZKQzpY2
E+ipZPrXxe5pZ93W0iqd71avGfYDlK1ScED3l5VJkb1iWCi9ncbr7JdXdcWkKmoQv+YIS28VVdaZ
/9IrjbS464rlRXk8/7L4SWU9u5aum9z8dIdW583p4y9QKBW2bvqLM8QB+oXORwJT80/GojI5B/FO
QnBVVPE+2Ip5hkKNsorX6vGbfjnzR5vTsdA/DPQfhYdNUieZ5KlvaTmRbuhPle3vuns1WTP3har4
eTNx99uiFMED7VagHh1x5+MqyKSIjChEZUVWlnDEYkIZL36WqrsUTdPiBXEgL/K7mtuiqnJ4L0hO
1FfuIcRq5fgH74wk//9Z9sYTX2hq8H9KNpXnLfHaTE4uOzl6+d6QVAFsyW4xU4uRzc7PL//mQa/9
nUpmp78rKCGbrVvKvlfyp6itjn+FxLF6EoTUdCawzwbu5pB2olKIlMI5SKxL/nWQ3IrWO7ra60px
6M94BvCtiOjI9KNl6JMSJDY+0bAPP447xTNBaW3Cv9bv5g8rD+zvcYAAmXLEptBPeKtZoLsgdXxR
QKtqVbuX7SnlkwaF05Wpgyg2Rv4nQSeXY2Rq4ZfmyjX4JKL1XSV25bZ3cNaSsim5UC7nqQL0Kig0
DaNWtQUHBuwB2Yovb4Y1L+43lHxoFpH+6I+40WSUtKC+HgkfAZuQvzXQv7tH9yPFo4KFpnhEBm11
YeoAVJVhj2NRXRPln9EkM7diH+r6wLrVX36zV+Kk0LLC3NonFKb4lB2WKyNT9jLKp83eI9z28Kk1
FQ2W3Fe4aYlxja+VFpMeliFhrnCZeUVfYnfBkQZMLup00iio9BHkdxGLF3IIEGlVZFr1CX+umwFT
tueJoSDObR3JqwkSsdqPiu/qdaHVjiIHNU47ONkWRv05eHyl2zl+q7pTeTb+Fo7yg27CvJn14gnq
q2AkaGJGvlQVxmxf6J7D5ZpuXdrmZrb09iA5s4y6lVL9MvGWsrtFzOCJm9JVvwZTCL4HkW0Iq6yR
XJ/6g3CzLnPRQp9E7q2ck2bGZQ6HwV0zDkbly6umFP5pEgjQjvUwj28C+kNB5boSSnK2F4+94BV4
RtqvnMtf418GBuAG14BTE+Y1ZV2G+GZCN3NyvX4GznWHU7yFtz9QtjUvfdWo9OPfUQcKaqbVkxSV
orDMvWxYgy26x6dHsV9PC9sE53i1oHXcFDnMNnBReJGz1txDu1CmBMekMhKWuq3itQIUI4Q4PhhC
x6illtpbSCebRzl7bkxdPLcqmNT1g9Do+ZUIhi/2TH5CzNQDtjkOV+OAWHV6teV4EGxnjfnlawHR
4fUGZp/oYlhYCGtMkWAne4QC3hzveBCQ/ZCFAs63AW3SlZI90b2f8Bk4YObesJxXqUlN7RbByLr2
qtwfUfmztPIU9/aAwlB5tH/yxNGdkIg5RLosSYUAxq0VBa1LuA7GENYLrAFEbLwjIPbp7X6Z09aH
wcHPiH7zoAXJ0ippwqno8PsIi3OaAbOejqdFqpIoEYUINDBdDnuyZExxgOXx2bMg4FnHLab4TtCU
KJhiF34tUCtuI/DA0RINFm/knNcZzT8Dnx6PjfTC/dnkpsexVgKbwuF90U1RTSR3x/QP8xc9H6RV
fytWgQ+zY2rPqMuGZY/KY9TiRrBYPnZgOLEeea3jPYJm2L5WZDwKiJJAqD7Hht12T1A6BFtUo865
AU2NaOxry+ZSnsasTP1nNH/qC2Brt7aCwuZDBVUyOfCUXkWqGYvmxl6wW9ELtxGatP6EQeTpKyxx
XwbvuLciFOgjzw+ft9VSRvRZZc2sAKP7n/HoIhxNQCunxbsnuoVUp2am2f0OvxbCJ/q2ilan7mOg
x/zIwjAu4QU6HfnPPO1gK5xHe/lr/I1GxqhC1gMpkMDjFOkcZcOR/fMeiCtL0eLf0SRL3blMNONq
MV9Vp1opXBin/cz+GNqJncqg9BeyAzpHe0R0hHssojzclqt/ik4C2UqFprhFkRhogSiK/gyR5I+q
RPN4U06eXFrBy60zrhoTJKdr8uJJxGC7QhmAMDYjBX5KVSAgi4nHN/mJLT8kuEiyF5uW94J5Rphq
BTKVM0ZJa6GBd0A54Hqn3loXPCWuClgB9VsAVSBafWrYv7ceFyLuEK2hakIjbg5BX2vxAB1/d4Pw
4hZWsaaI3A+DZUTlkztRZgOeBNa+FZ30kjinTerCwrthEt9GRiFLFzt2X9hXdmvlgbpe1bSZdEx1
2fucVotoStioyapBN7UBcO0XF5V3ZPEh8iW3VpSzzwdi8qGZ6DomK/sCG2zmsekuE/9IIvB6ID3q
vCGAPqdu5ykPnWqMzqG4NILneqMnM9vg2hvjScyk+h4Ygx3D/3V6Br/BtaPe1IjtlQpcrFb/jEea
RM24/8FB+PhZgZlOXUaznEpmPuAMrbCwF5NTaXlaoA0qQuLJHmYulBa4h3+KqnH4ZxIeuSJ9nSHF
DsG35PN+w5L/6e4rrpxSKDd8ZLfgZ3h+Gy+zLaY5O2VjgLe7Y1yY2+fYe7lKMu4wQLUCv+9C6iaW
zxmhT6Chk29QALVjcq7C2N5/CqiO708IfKvaUAhFIBvjkPhQNzLwKLlf/Eo9jYTcEwlS0ygJEBHu
Zmhs7DKA77ceJeFR7AWs08SZF29NOf1B6/YeFYcEpRcDReC7e2ArjiWWvJ5jDSbXjspfeL1h7Y7I
EevSKs16jtNYhuagEfjF24o8+ShUnRZfDbDIzxlkBisqnRYfsXCJjszYLteSpn5LJeG1pO3KFQ/N
Qg0Iz3Vwo8g01DGIROhDaqwnhONxqf5xl1n3dH6wQHkBwGVUl6irX2IPs7fm9Uv/bHo6efs1p9l9
ii9R94zBtWLG9IRZk6fvAJ6PzbzSvNImNbIR60nw/igTDu4Ta+qjry8RapdZJ/vuV+sigFNF/m9G
eYupMvKgn5n78VPzvipe2QC5ewJSEUXIP+IrFeuvpzrVmC02Mp/hCqjX239erMii7+K8mWJ2kPTk
0gdoYxFSzuCibj3kW67A7vVnuhiXCCbfVn+5TxvI97aWiZG9Xe61aQglAcnC2yjkY1lZ2phJuHOT
GSsqhDPXcuXSzvCJ3fcKt/ahPZ77jfPKKN0w8DqI5q11jTCjxpNV+Mk7mHrUmQzcbAE7jDsxFAui
y1GoZtOPRJDj5OgRRvMK0GSY0/1Rv+iiSEqDuSuAV/qX+fiO2KJtGSEP4lda9+iid9t1C4ADopLL
OFHsiSFDli0/PYOBW8kSlSQc3CdNgyqYbfEX5gapImmr39Zsfa6xNeixiSvrkujnw2jtNIpJTWXw
PtZXm5KyTvq50OA1v9W4Uxyo9MLM2lHz9BE62xmW2KBKwuROkYqX049o2spsmWU3W+21IZE9j9X0
mhCi8wT2AGlGhpJEoG4yj6/4H6T0lmiZZq/iMBO9xtBDerfEguh0Wku7tvs0mgmM67Q6+hP83Kgf
Pr3xQ1hODLeWmCDGbKmIiSe32X1vXkE94UuUBzDckQCBLZhuJtoINwNjForDVG1EmIdJ1foeajBu
5PjaL2OQPrFxxQ4XnXf8Y95M6UU2U95Te44kNu3or+aBOWV2SObeW7xfH0rA5+xBnzFfkBCi4+fN
HByjoGqym8kJrIIV//IEI2ug9N7XCAz29jmEdmhUcA1Zsd4sMJuiV4PkK/PA/jXBHvxRysJBr4Bp
+PyfljrGX4w7fgyjJX028ykBgs7Utp6X3tTh8VZ/hCrCqGxe6RzoODPu6FQOa1vFiwe7ITrOvnsQ
os/TFogOQ4Qe0vTSDXhf6VXfwuFPOZQ60To94aU3xCjnl8dU2DF1x+8GUfXjeYj3gNMQm7YXHmhx
wbNk4X/sDGWNealqGIhkWMYlhq8KrUQ6BGuPPcUkbbfdhGzq93f0Tnx3dfLaRB4pFxuLW7mECums
tYHeHjipbn8vDd8BLv6zTjEXsKeXyXLt4doVgwYR78FWrrOEwqs7KIl4ow7SpDdRhbAj2hhyynd5
n88HZNPZGZJ+b12UUqHd6Fcu4Bdpkm5RQZwWAaY1NXhlNzsbBZdRObA0U3M7DPwll4eE4s1SxScr
QujSOMAlhIAc6I56yX0427aQjYxpA5IE4T05tAaGYXWlGPa3oy+ZLJ3kDztGY7MQwl3GUcm1NAfY
Syen4zppM0HKg4Fexp9BI3fCkW+FoJEuW5T4lNLtBwHTshgL6TmexFlRtsGIsXpmpED+WJqryHGY
0fg6tg4UcCsJaQvuJKjHerZQ3XCP+DcEpsj94Nmfz3iZM9Bogyv2sk4X79VRlself0WYZr0uT3jz
83P37O35gK85MWSTkhwGRKxwtz3gtBXjKPCbntOQnvIsxRW+4rLlwiHv9c5rXm6yzVrNt3dfFcEx
hW9UO8BDrZ6JQRfi02rva9RR7qJzyXrQSnQBJka2gL28lT4UywAX5kLCqW39a34d6bBeCSaoW2Pc
6kEi7gLhTLLSJdvAEvytMA7tRc5CEVz0MrVxURq869jF1Iwk6TM6OyuRJqcPMsIymR6Y/iIZOc4s
so9GrMQaCazt9jSqc2IDFDt1MglVqPkuEOr+885ViharRpruWii/p1jKwFRfZkxBcziWZ1J4wtZd
C5qDeW/nkH1BVWsQgy0C7/SXkTFIUldTiyVzrzOikBJis+s9iEphW6NsPd8ecPTWynTrN2GVfaZQ
PUljC9NvpwgOetOeq8S7cPz5QL+w64TWpwWLPfGH7ndHVsjn8WAntrmD9T+tL5Om7vmyM0f+bI7F
YfyDIWdlhx3IrwAhxB7kUmQhlfEKORwGCQxTa0zjIe/WVPGuUxI+EuvnrRwZkGEZWdE8MnzaXOdu
qrrebTxukqHz7ULrIOGuFME/5dcnGg61VpfSsWUBoSbvF9ZT3RfUlq+5vsoBLpgHAngowmrFfJ4W
BojcO9bF6c4PhqaBF+BRi77GjPWSF6w73gqZw2fuMRIKQT50Rwe3JFpMFCVwzGm84Xh8tFAg2Bb9
imzbh9XLiQtPxAk0ml3MVmNiAYBhCraoZfuErUVPv8wZpaDOc0ydJlMlYUpzLQRHtW6eeHN/maqB
FOZ7sqLTbtkoO/rlTp1rwOtXS3tVV/WC60GCmR0QVv8Pz4nHV57I8l8aJdz3pujKcu2iVVu08XI+
M3KNPUmyOBm6jCbQ7sAi/V8jG8xIS2R+aeTIbYISyKEaJm4LiEu0Vce4/iaucb3If3NUweLCFCz6
qXMQxZXn7FnnYyg8txOlU99Wp0BiKiZS1NGcvEnt8MRNbQDIU8AVniXkeJaj4cZ6+upZwU1bB3Vn
z7w/XJiHo1drb7vA9zZKosk9tc0PMOEhUgt8tA4uqlH9ZInRAAoZ1d1SzFoZ/0jDLu1TD9LEzPEk
PTdNbJ87jCAmLvn6pdPrsrB3amkATVvkPIXn3Is++BNXUJdqr11InfxNVqzMyv4+0Qj+Tx2G86Lg
lJdjprQwgYd1CxX5nJlhdy4xWzUjtOwWm4E6Gi/RMG8fpKJtfcWHKA5yaMPrUs/NBcSQITI3nFw+
pAWSjOIVgwvZtdfspoQvOjXXWdEyJ9gO2JAluXO9QpaQa9K1guFh3o/zh2Kipu40Lik9BR4EMuj7
C5hKlDzugzSGwqDsIq1IUTnHegP0LtCPNFVTpd4ku/Z4NBynoLWKauU5KvzGFAV+YTqXqM3M5OwG
T8goxOfkyRvxokrpW7aDMXIrY4d3fnGEN/Gg7Ld57WcSUYNN7iUQ6PGC4Xz0rLaVLlyu2py4+FGl
V/bmNonWbJtuaihZxQNNI8fHZeET5q7nuTzeJ4vS2rYL4BvpWK3HtvX3xIaPERt0qeDdSvJU0eXm
JCtLpRm+WbI0jAzELFDd/3gTgCA7ufNkkNX17uhc9lDczZTaNleWZAnx6aW4/pKvpJ+XzkKxIgHQ
DDN73WjIVmZ6SpGyBiRdPWW12kKzxi0wx1G3hSHcCLadkXTXbp3J2PUdc8Vx9XafgfiPf8JjDuP+
IxTIyUzlwU/z/JTVhAC/6O6c9wc+DXfDjGB8b4OLuh4nv2D5IBxkm8lstwO9ZKSQsHCOuoc0t36b
d0RfO4c6KQY5TCx92cH5lZRJE6tqWKHvGsxYwGZgQlaKKr1A8rKv/sd8DUAP8MbGoUrFrd5XXaIT
sRzYN9vAXGmfA3PNqQrxaO5oM/wBtA4DaeGf7s9JRPoxCp2V3o52+J251v3/5Az5sIRGAARTZZBP
tcs3zz3NWq85oxnkicGSmBoHrkw0H635vHt29veK9kZVvP3IDbRz+NpE/qWFfAm2TGYXwLPWQ+y5
R29rpdOXzGeaHxPEQoog1bUXghf45mwE9RZJkY7U6Av+eT8q/owVlRR3yiNINVslLhADJ3utOJWo
2+nwukclpbWvWcSwOVWI/Q1UW/NOWSa8wpZw84vob15X4L5HZdkA1ZrmQmDyWbwwPZkbYUAA/AKV
WqYg5Q1xDaY82Fm4xdvIrNDqpgWv/tXP9qO8Uebl85OKYi6nlCnmjGKLyw1XzHKbQNyo9mRAHVRe
PpXdHDyt8zoH889lqc+clVy5kaARusfWi4NL4mcTfLfu7HuGrC2fbNKPLrUTDQvmN4RoIUuGgp+Z
CimdM3o1JE2RXFa8dQtBhGPT4lfvKGikG+S40fvP3Ju+WTRhx8bLaBKOkYO3Zf6rjCTe0lbgTj84
A9gae1tZty/FDm2TwG2a3nn93nMatsxK2CpX0AJRFSGSZrKYOYnXaxdRExCZddG/FmqrHgtqzySR
J/Pv+Ewxgdwf7uq7YfSglmcGTHP0dfZanBXuJ/MMDhaqkmZ82Ca9g5Hl+/H8+l+uObFg0pXVBL9z
ImYnLCg9JkHXvzck1YDD8oLvasTKXYvrZdGLtcJ7Vh3hQcr6jdyHGUNapjOB+/fR9eUoXT61Yf7J
lbbZOtySW8T+mgRpcade1BbXUPvago/+mTo6v3dMtauE/Vah9ooNX1WBG5cCf2cRRm6U5KTu4Tif
4soZnPlp8U5BeHh+4/55KOdjfOHtdWy+KCDZTD17rTsHFtxYuZoSDgUyZCP63DLPJzHQ0Xg3dKeF
0A93yJTbIjtGqrO4ttE3qMuc9uj9OCZvmmZ9eqB5jN3bHZqCobeDauYkcMCY6UDh3PCPtzekAzvX
kCyfC1RQDXtlvedz5IXIniSOWZpPrizPL/J2xREdQOQRJ+gSY+tL+HbgMVBkLuXgPmQ/KUfrukS4
N6FngagxN32Qx2HOYBr4HZfuKti1bIWpBdJt25m2K6GBbmNE/t6YXkAE0o6fcl3X4meXKBaSjL3T
U9iVEGPyTGff15DLZ1/9cZ1QjPP2Nri9sUHeAeClI5lKD7lv1PHrnq2Np7vAZZIDeDQ4p6feGdQj
D5o1oNNcW51oftoh51rC8EwgCfpeHljATL5bZSQY27p4Ctkarqgpjpz5xLHIV1MbPWDZ3TVXJcTL
SpotS8Hn8dieVPic7Wcsj4ghrF12v1b6jOOkGRHvcF5fnBKmCs10nJyytIEeHbTOmXiKiC2ud2h9
pmPX8W5RUifEqm1R0bG2R6ums2HhmocBoixR8cg7pe8quHcfSjpUrFivsZ66sW8uNYs3jFOAITkP
th9R0c3y1CCPTf6z1h8mmv68th3P8em0/p0BvlcM1Vr9Otrjky8mMJJDpdFbIa/HBMk5/gjr0Plt
FyQC4/XS8KOElWOT9Q4AbJQjicrc/nYjAwj30mL84ZkFwwAx6IMFv2Sv/jbjsIhLUZLe0zqY4ohg
8iIVwglillVTt8QTUaX1h7PYTd0Svk7vUYlhlGaJOE9pgQ5trZqmCUWjoXhJJlpnPJJAL96MDu97
EE5JPItrqRpk5earOv4zh8V+WCJ/pu1Un2uWrdLqM3a+Guuuh5KoHx2Ayxw16gGd43TxzH8E3qX8
a6vLdnrfQxxZxkAF+xXzK87eGpLT6ZbyNdHEjJ9Ct7lX33FAYnxrYDjuU45xP3rnv6pFrCg/5yaq
8mepcDtfiR9HwFhzrA3d+Cyp6PSK3wpNiE/NA3xi+xYI+rXfkP3gzrXR6qC8YqPl1nkweIT8fXif
zefUVAPdvi+qiDn4fBF87m28V8PqK0PtYe9mmKpoDlLO+GJF6DXXGY/WTUxHZFNcq+gvFdxZenGs
+nfpNDpSGKhGbrxaLiO1U3weFxBjhmmGNqESZ4X1adlUdgDOJr9UV5QRpuoVxBg3RLcNe+QTITer
75ML/4vOewYAS/rE/Jwg2sr6PNsJaO9Vu8f5X0CasCREYba/pQEADl6MTpMNa0fAjCqmdza+q/7o
eU0A+aYFb3L7mKWglJhEvEpWJCEamR/x0/sVhCTe2N3qs/dcTGPw0buAGSKSojbodibl/E3NfwqY
jQ3rH76D+ZPMdaX6EYoKkcOH4efhDBKNDow9qsbm5kKbO74JVa5nmZleEofNbTIGSEF0w2hbM/V8
WKXjb4I9x+twTw2Ll1BLo+5NgYhEMOcQktUwXTKM61je+IrAi3fhltV+YktnSRmLv7ZberTxPz1x
rlYkSE0NHN8JDcoCAjhXxL1ob2OFm24TmXse18r5peP1qq4JqcWkHe2xAK4PS8U7MtL2V6BLl5GM
hKaw1xY/gPDoymaxPHjk/NnfFTNIBv6UsPusAVfyLApN6+T5OYSVgaqi+8GwKQN8GQOrczOs30OI
RssNOqaWmSUOIwVIwEMLF/CnZlFiQjchodqaEpzNaTdh+YEAOtcCpj0scWASWTqz4f8lOqY/vNOV
/UDZKIbd4rL1PkxhAuMUm5+WSw9tkWTmsfWfLyb9qeFh4F0DRuRhVi8r2yO30pqQ2UCOmo/2K+nE
YRbF7zZHyWN+a/1Ae5QfqnSx/glQwAC4r7GYuNyv+D/OuBRs27Xu1bHnNPkwf0IHnmcnOfG4lnyO
nrb3o5YDtTR8penAoT6RP72yrb7J14OM3msb9LIKgKeqi37oyhX07RrrICurUqs3lML3JX6QDvpn
ITNzp2FJ4dRn6hxVlQaIqBqP9+dgIMADuRgFhwVm8HtUSc7xp03zfzvOoFP/ivsRmBZ7IB4/nz8+
pSvhXSGwzxMJdAGwVbgO9L6P81UMBMivDJsO9kHt4+7zapTe0UR51HFejeT3J/XPKS3QXuXm+aMA
BNf/dG6PTtLWSK+/ijngRnDBX84BRajYOfRERtitGiXtp3jhVOegornr0WsKv9uumnxTgTsmVzm9
RXarUQNpNYYz9DYXV1HI7bMHKZVao0Xv9QDIxHrve6pVIGglSsMNqy1vyeeW4wQQ23KeqoRS7s02
zU3tK7Ik/q7eXeTY2/L3xB06bP9VcNHiHpxZSo8illVX/R9cGLhyRLjoFwx5JLxGkMRss8cmaip4
+08VWA2mEbgeZELYct4XmYe3+KhIXOjdYXX9pJZj0/9G2rWLziyuFvd9pCzg9+r7Z0iRtrgDn2tm
pXM0zzIOjxzHTe9tIwBhvDNJUIpTbEt2klrkebxG7g9Tba33DRpZl+2jFxjl8z25bFwXI5xSY3pm
v0+nz+DOqT6d6ywiK17F8WHuFM6bQWIR7AGZO0tf3jiBp7cnwEFH+DsVzUdFBZlTBhJO5rIz4yAZ
H3Y8pw41b170VgXc+XJJ+w4VWY4Ud4sfwr4r9pPHe2j8yTBV4UErcEEkYzpAvA/Wn/LkHCBr0iEw
K62BP5W9bs1MG8SE8RjFeY9A3jRDXBYayCAQCjI1FTmuuOAHM1oJWn+jnBb1ExxY5nouH/oRxSCW
FPU0AYG3lB9rxRpaFkVWx/HLKJMi7IMuMcyJQYkA6pcL06LQGQX1BbD/rDD7S8BkdJYabsWr5/5c
dZA8PnbFU9/mvNbVpNaqWc6a9G+V+vNZodd0tXrxvnQr1kDN05sxIy4RAJembUEvuYTnJdON6Kp7
R+pHwlmsuXZXNoP467kJ3RpHz0rG4gE3OPB5UhGl/zOuq093DJsysvHW6KbFpWe5el5pZe6YXMmL
GoL4d+AbLWFFGt2fmogr2aaYJkHpCagrKdiqYOflciml7WlwL6UA20eWgXd4dq9/jLoLBzH3I6Wt
Pwz5lSm8o1KTmLxThnbW1iF/kpVZUotXoIR2Tgq1vcNRSa/mo+PR8/KRt2ALpnQ5FzN1Jcldfx2M
b1f/3EolAj8kEunanyd/XbCNXnyONeuHGvtoyzjDq3hrxyhYVshB6NR9RhJVZLkNHVFopRNF4th8
r0Ea/WON9KdiJtCAPGPmsuXH6J27VWvpNAAz+t81VDwNgaT8ctQSQPY0LREDU98+m9fpiL2MYm/X
7P3gBCDnOjM+G+yq+KK112ZrO8YMeCvcMkLRXxCdrv8Fawx40x9Mk/+HZ5ZLKHkbbcTeg9QTrRZo
lJWdVctLix+5gwpRIV6vGxwB03ykKRrD9Ex07YS7ruMMNrDHi5L0rjV4hTlXKDXgO25lHvFYGOfc
eYDCgFAKSHYqMuQL03n2WyIBPiPpDRTOSg/P4o+wFqRiWZNin+l0DNC+m6QiMc5wM7csxdyIa+DL
TtenKeYDlGDUMMJa+whix9M1gzxM0H+cuyZ8bUAEVstECslbFYXkm8zqKMFMxxqlGXUWzSUT9KiK
jB+n5GgVRy0ng2hGCBByEhMnjCCcgZbuIIiZzJA3j6eYz2uSDQjFURabl0VPU4knAKdn2+VPEHyd
nazg93ySaokaoMW32sLgTIXKkD85VDrtCf0CLyHI4rJHNHb3qnb2uxoqE68o8CiHqQLiDn3oVSXP
m5pVS+cpccHHc2dPNASj7yiUuaM7yhwWFvbpgmJMpvP5b4HTCLWiVaH8LTiIcEQLPVuAlSgITjXv
JheBb6qNcFAkCFOHFpFTGZYaYHwGt1/vrHnZEk5LUa0+De8Rsl+FE5zSZpXMyf5Ya604uIqn143k
cllpcDc7vqX9dVPwttXkUP0Q/VLVL2xp/kMeCzAtYBu/q0gfSn2wjbR3KQYLCImHKzaR2qHGqEAl
3vmabgZl7yQpok/8uz9GE49e8Qmx3FR5Egm/mfmXAOlmXwieIC7vZIVmHXp/0249WozUWK+M3AIx
XFXGwLcGLDKYb+WTCK0n5+3HClQEpFYFsJpJHVdtvoO8LN5JGrFDpKlcrB24A/B4Fb/mTy+TPdda
aLxEb9onzc+xE5B6PU/uVTVLcP8epzU/d+1t8mJJh/0NNpPlM0X9DUUlQtXBnY4kYHecBrzlZDKE
jUG8ayuqyoDevHju804HaKZzcDLtCBuJ1MerLR2gGvnJM0PFONotXl5SAk2R3zrl0FnfWlfZVTyX
y0fmxbrfGoqkfRkJsSEl2MRaOEDppxewMsQ6fMyT/YC3ruB89mflff5F0u4whMXi8Wo/9YFz5k+z
nkB3Xb3HlyWYgvQbe15LaqH6GlrFQ9ep+TK8vuXTxo4Dsgvp2/eDm0kkrEctwYDtrNq31jgM5LqX
XF/fLFsoUT3LppnFn4Cmgb5gISt1D/EDG/UwnCD68gEcAPem4HmAWXJDW8Zu3c7rztH6s0dl4Kwz
TcHDWsVGqnOFJWGKKY5KaPJdlQex+PiUyTso6xouoc5QFLyo90XJzoZnTeMGsZ3J2WZX2vdw8iJT
PvY69s5cqWfKICCtDKS2OwmWxc3BbR3sN9LEFWg+2RbiA9z5KGy3kGjk58MDchcHdXq1B8fc6Pf0
5dna5BW1B0/+6cxjmMqBxHcC+Uc/pltha1EBRL9QPi42l+SbnWG+q6m/rPCEgU8vnNNxgzRiEU3u
IKr4i0zdl0xmgLnnOa2poLpW33Jcu8tKv5x0IUqwBbFx1hWd+wnkGEblJaNhE5fAJBRl5ZJ2o0li
smEyw4ubHDURj+St8s71S/eLw8mS3UwD2A/0/kKHkdbv+EkfiRVkneRuAvhHHXVn95kZ7FyDNmwu
eYtagIJn/zNQ8LchrZIv2XMVZ+XZt+sylAtnSK3U8dO0z6vZ4mwhTrcBNz5oIhpOrxMjW1svTt5W
sJYdRUWU6qKJeKJ/A/satwmY204TNSmiWnA1bNZ1AcUJSpwmVJB0INgaC0baBKxibRlmBODCbfH1
81hrJ/a0qH313IsHZqwA3d7SpYg5YEphMr9J6yMKTcwZ4Gq7ykBzJmGIq8btaS+GGKxzE3OEkzSb
WGjAS95IA7n+eWMjGYkhNVrNAG0+8p7LmDLO7OxNlklEvM0GmkBrTiwfey+3NSlEKxIyMv73Fel8
93YdLi74rL37rhjerBYb9MhHmonl4HZ58AhTqeFJEiIPF1snCnV8ZHAhkyp5wMyeaWLFV98+QxuP
Y8BEymhMpRcC1uxNje30rXlfXOvvzgBbCg/Txdlun1rNViWh864mH4GvfiT4BaSmBZiTr/K+WBRm
B1Te7bAeTFL7l1cmRqLE8lgzPQmKEXQaxhRVgx6lcC3bRfJOn+hXfnkDgSz5XkIc4RKlbvwYYiMW
aa2xUVPa4kvUEWQOddDmsEp5C7D8PKRp6rZe2s+/+BiRkUjif6Y0lWskac3DtWfmoPMEO9mY+1kY
04Ubbyx570E0X8ByTGQy/o3khROtB36CZigF5RcltVhFGKlbf6v3vmStt2GOCKBr8NS1iFHj7l07
qDdDvSS+uUkT5A1/QDQA/JfHkcO3G+w+69+aSh2SZSO5xraA3SiYiGXLBEmypwoLPfFVMs1I/bDS
EpYIDXmJuNH8c1DRZB5eebVWWEDiNavCYnLB3hTPT1SL72AsCYpc8PtFu9D3kbosHwnwQHcm1EWj
pTOEdxQsyX/uSGxJKCRTLPZpeiBFujRm2v/FbPK3dBK34lAEQ+dF1jyyHsB9eGHVDPT/uLiThG7E
ctbjpFpvzX44wHNJenJ92fn5QG3jDDH+3ceqkJSrqizZ1KLKAfUSN4Px6KXjH6s3Sj4MEtzbj/O5
0LxWP0OJfOnLYbt5wkPbGzs8du3B8v3gw+5WxvBk/wdczKWjJtM3re10dK9PYoECWPNIXaLxH9Qd
DuYKgZZ3A8OL5KoGgR+7QRrKPcI3G8UbW+Qd1lTlVh0yLhFr3mfFrQDbY4KEXgVER+a06wLbdwpw
9a9HCmT3JPMVknm/k2HtvqNgvFKxbeJ4ZfvKT/aGv6dfYEhb6rbvoi6xTZO6tgtn4OmeBtK0lS/y
wwDhyIArjXbGPlFRLKN3CrYDKp/qtcHa1/I9hweAm7WhiW2J+lHIRxPwme4LGA8oZx+SUKSuSryz
xz/4iab3ruknmlBeCZHwFLbTJTOPQoQ1yQl97xv7gMl285cSViqjNgM+aY8wjIAKykxNfpYWqNrb
3iMorJoa2/toMPX5enRSuFDSoMxr5Uh/BVcS3IK4VV9svUH9iuYm+4/rBMJ7Il2Eh4NZdejYYlhf
bm9VKrPQZSsJjTYILpcIIq6/GVLgP08lG2ukCnL/vaIbBxYUrXf+29qmHK9B3y7IQ0Bb8sKALhAB
8I/u6bSzbV07JkvvkBIwX50UlTJjfQaaakRChKKXyUOnEH59zsObTuyL6UFqWWU+Ai69hYupOVkX
KJ9la0NHPTfcGuPYo8NgoA6/S2GUr3d6BJpGpWTvlNiUnNlOFovTHl5a9a7s+Qilt/rJoh7LzNA1
e+DDtVqm7nYKyf30A/Eh0PkMWrFRFaEvKIChZ4nU369RC9o5kNRlNJZQt8LF83wr+VqFtV4fPXiW
uGTpOT1vWMlVqnCQYkhxTGS4sXRrP2ZicjsWzzchH368/LLRITaPhCae4aX7k+cHUa9g2yrlRRX8
NLeniPAbwIUDSkXdQmDMnvGqV6fvV3m9zF5yPQr/a78mwJQE79zFx8HH5E9E1GoQPo9712U2CmEf
jQ+ADH1jmvrOWSa6+D70bnW+RKsOHucbyOePxYPw1offiHnIcB5qx9PKGXyig8KNgpxnOMb6DwTU
y8e5EXJVWEnhdUP9D/F8r3vQz67mqKZx0xfkXdFc4tIULkyxdpok9QM8SZSg499A1sKXf3Rp3XIm
ngMn+CALJYmLiSJSySPnbEyQCeIi3m8gJmK8lKuJ2bo30z5EFGlqOuVgVygFSJWz/nKshNUebTau
adU8tSlHWhojg4zzo5g7X1u1P8BS1QiVoeo1sH2wCVViJp79IfS+qXkewXq2A/HtuYHoBNdaZf5i
1KKu3G/iseKXK9NR+GEjilayJksznlaUqvPSxOiA4dnpGbyfVbuSj6GHIWM0Q6g8S4eTt/U/N/yV
UJnfVqVyw1BMtk0HVdbepfbPL1/io5Km1C5wPZou8FLWEi3f/z1HtvhG32Q4xZc1HZQkxBzYmw2v
DOa67C8QhT81V+vK4DWjzZ4A2qy7t1NVg8KTkUSSvo+0f3FKsO7/fbEEFYRU9qWF7ZSlSSXr8giI
3Uk8sRVSgUklBUxBTRzHsYtWZmzaNB1/d/15h2quep6l4fnySUH4BnXQJSBzeZnH5Px/QSarWvyC
3HjmuugVZYmOT+JovsT9hqozs2PXax4JvjoKSulzhKIWP/1n0hTbXKxwx+dMkHmYFz5ra3iv9YFy
h1KNqb2UPuQtO/UvVOMQJZkzLhUpcbyBHHrVD2sJrs5XWdVtBGteLBMCRvCe0g+SEu9j6SWV8hhH
xlAli0/GLCM6W9Zz6eQpDVIOSj4CGsBmqpD0wyL8D8R1cu9XrZlch+UcEL8nH+d4j9SmyB+myICT
LRrCwR/672l1xO6i7Q30blNfH90hiXGRGeMghpb3tsclbv3lBybqPXn6sorJVi/dCqBf8tpnyR5O
fiFGkQzh55Zf8jVv9Vq60FELibuSGljjHFZFAmZA6hFwFfS07yW+YQgOlFA84oXnYO7gl54iiPAC
ELmqalfa1aJWhVzTtGXmtmgtpEteYHoPzLHjanPau+oRApMrdJKvwDsH5aiQuLKNf51mXhUHzlwL
eNZqAgNDXGPSbwHh6aqfTki2RNsDGqd5ZnkXsRHo8dRZQF29P/xkww6TfcKKLEDxbjIAd0OQSGfm
P3DWaNPfqgypMjDYWfKB3YzeYLj7x/WM29p0/xeab7OVfdbj1eM0M0hfK4zRR6v3Uf1HXxsGKibQ
ALNTqr2AohLoEGQZEwdRbE6tx7yruH5Utp/xHRxju+6ppND8PUE6UmOgFI2j02LbtuhLAm59sDkC
D0gEOLDkgsf1AGe00dlTaUMIW4+qkicp0DN2nJqYbtZ3G+t5TNhBg1RwpEDT2faF29YzZuZf2wc/
igb7BtKECPx9bAVOoMnnVuQ4bCFoPLJRjcSFzAxAnaAnMJt+kkOBELV9BCnToxTmNtLDQXgS1FAp
1b2mt68Vkz8sJx76ihhqAbb42evwFhgAw3NPwkE6tp+WimdTm32DEZCWS9O7uDuUh3KZLkwsX97U
M/urg6UD5Xf7bjjcPOoL2Rx+UgbSXQkAeThGvpkninEYQ8molqyP4T4AQ2gRjlyGRim/oIEmsGf5
mT4FmWaqo5lU0a3kIY8Op9YsNdSTfr9e1nap+J2+u5D+1x9QWHmYkN5nSo4y3oA9i2OS8vwf2i5A
/In27kyoDLabAqZsm1jSK0TYj392XvGkUWiTQPPM1Ttn2IP/wtU3dgdG5VyJE4LXxn0NdiAHZBby
XrlMssyh2SKdjELU5bEjuZqn26bsgrq8HJzUINRBKnC7oAFhaP1SkeZJVLZ/jWYsSb/+cwh3Y2qw
IlPTCKzEljTmATMUvaJuuNWeQcyG7pbs1NQCGHs+cB63iBozvTpGuIYFUspYHOdG+MvLFFJGtfzV
7qwExKOmhpp4KBCSDpVXaDEdsNirXlfUWtXf9T5dXAvojZMq0XjdzsJ/Zl2yxE+8csSFy1IhFRx/
KoraKoLBWYxK0KzZRMSJ419OZZfBcxX6Cu4sbHCEfAm10L7mYIZuIitsuh3oP8WRcjiqMDoiQBIL
fMFNyK1mU53w5aM+hFM6EuUDUVAyj/2+ee99A19aEbCQAOfe4pXU1HCN9qREi92NT82xG4Q4G1mO
oKVG3SsDwdvZDcXx6Z1I+7/i2DuKOqyG+M8jTWoyttZUVh8WHXEPUHzVa0u27PoikdK8Jg9iVQ3s
v6gqDZyjrsuEgFY8yVdGN3KTkoWftjaqlvrxnAfD4ix0IlUqvL0wMypJMKaK8gbprdFtMTP48UZr
5kt79VVr4JhI1o+9ZkJITZfuMKwOrOJZxlJ5O7Y7I2FDMfrYT5UTAASw0A8WZRT0k7rgWUOUo4yx
jNs4Yr06G/1F1XZMX5/sVXss9lXCUp7GPNpr6rBNK4Zkem0WpIG/IMre0s7pA0Zj5ojVw4YeJZ+5
3alTM80Nhk8OU75G1612BBHzxusSfLwsfU1w1NK4h28iIdAQLj4j6cH8OM1CRl6MiOPp62nbjAZx
nhs9Qp0Em7Rwnjq9+7C5i0I1IRJuUDD+oOXOgF/e9lw7HEppZ0ww2kuShmifqqYJZB3A+FmWAxAa
vi2XaG6+0144I6CHWbkxOh5pgU7Sge1CXK6DPfh3CQj5maLAQAjXEy7FomNawSXZwK/pCXCd0H1a
E00y2tzO4A2ekY1j5B5JYeVirsmyqcuN4P44AztTL9zj3odGTHqSdhOWybddQf+gZYEVQMR+2nbb
n6wYTz06/29MV0ta3Pl5qB00xBdhJVrcQBA2KeYVfPxshAMx42cWPDvcsXX2nAwK9XBSCnlOuB9x
gAy1tGlmWaITfKeoljPYp10jS/qNuivbWT9vVQc7RrXVKL1kJVu5dAOf8hMCmaysm4UEsJ8NNooL
IhetKncDpFuOFdAhx1DDvrlpDASgeaS3n8486AIUnPHaO/JBO+Y52rjVFCvHhpg6ZCyQopRXfVW5
L4PzA6np6mmM6mH9+yRd2qUr/LgESQUXCdw1Sr5/ERvgkhnThuZx+8ujiaR2hnZSWAjcQxUySMGE
HbNha6JVr8a0dTiOiZjeFKXq+5JNHQnlsXOk26QpY/QWjP9Z4ADYFc+5WgonCb9O6V1PXKNrhOyX
HmCaBdo0g2SM9pxzAHSrEJu/KfLgdEpGuv5uxrtF2NwoPSMxnXEv0IZpvHXi+uCEsip1IYOuChsJ
atMxoqk+Uj7sGWlJqI14GazFNeEE09zkEoeb/Zo7gd5kTr7XcGPyov8rMHWFtf5L839DV07x43vh
2K73h2yc4069NvzZFSXA7PN+Dm7Wg72NQtqhHwpuKogTLTNzdJLRgO1gUkc/5aOcjzd2an3mRo34
B35N6Pfa3vcAKWf1c9kpnUYUkO6Web619+wmR/a8luKCC2BUB8RF07ijImkw6T51fNJ/myH5pTvo
VA1LDjtZnyiW6RnI016PuuDc/zAq8Iu0assajKy5gLy+tmDPFZa7lQMG/Utxq4dfB47MSkoMl6RX
M6rK1OChaja6kS7Zpzki3ugf+ZniKkaVXIyG4qmx9DhZSq99P4bencSUEEeUdfyICsEoNH2ILurt
uMu5Ko6jepdBlGKwW0OBEgxpoSf/yCEclPrOfkb1b4zG5RzUgK2wHo0kO69zoF8MPNJrchm4QX8v
S1nMpaVc6ZA6/SFu0oqALxVN10pLpf2zzPUa8K6QPzcnOTEoP7cjSjnksmG8yCG8T09l4fWeHX0m
vGqAGiu+2HNUrDQeIEMuvGTj7UxC49bt+vEs5gMo2HglYtkAnH2DmYWGOwB+Yg/NTTVbpMKPFAZk
Mf7cZygF7CWUkRrl2a/pXT/VUG+Ae9TZwDxMZWJtKssg/iEfO4tqm7qq4IIK/Ekp9bFwf8g7zK00
u0ccRIKdEmtBYd+Ex+PlamDyV0WcpQsf/UCbNcUgQswbQT9r9hjyA+izXLklykqnKu6ZhIdFGgPz
MzXIMXCK4dsaiKKatnjmwWhWnaev2hTC1Ov46Qh+ppClD7SFNFUMMG8rQGJRhiikWmmJKvK3GWxR
mIWAKz/tQXWeBMJo7my77A3J8++MRVO2KpIH56wz83Vg/l4/MfeweBSpPTTMNI1AzqPeYRp5xL5Y
HXAWigAjoASweVzclXCt0Y4Xf7x8r3ByZ+4b2CgYmp2MfAxVbBR/CB8BMHx9graIsYC+ertSz1tu
wxBeZHq/BBPIGpW/ei/YvgHGGC0onZQv/30EvpmMs4ouoRZGqtUFFMSEcWEyeIUQLMy5KpTfwC+l
C4oP/2N/j9nd7tE9RVTXvEnJKs/YmsZArycf84PHilqeiDZHfdARWlQaNWbf8RzfTSsy5963NXO7
SR9UT5DulQFu78KEblfKVVbVz14u8/e/EEDqm9lQtT7OMT5GEoVOTB73uhec7NDQoILhcoIkEizC
ZYBvqp3o7fMVW0BdIuYr7VgnfKThIBNx5qKTvsMnKdnB1EJTQ5zXpI6pHfDYSrDjDFQhHTkF/gaw
gjzm9gOjI5L+CpcBT3wjxH/bK2uU5c8AvrqmmZJWGoKOZnJpHJxZCQ42q50liFWbj3QcC/mEIfE6
39gldViyDupt2au7Tac85vJFdPSWRaXseMDaEetRHySEkKeulNGG3iEWWvh9XQD2Y97C+CnfwY8a
21tBThv4KxffrRWldLFkWt9aEyFQN39xSgaTE3o3n73un8LGm9p+s9QCnOFH9JGKVoNL51gHB0N0
bocY6RciT94op4TB0ENJwS3pZwgTdH86cTm/U8LL0IyK3+vQBGlojBEhnOxRg3W48A9WC6mytMJj
zY15Fia4NtcIe/Kwr74fsUgoujZgz6AP9WNkPqXbXEgcOAjPnhWVxa5KnD3oK1VzH7bW7sFDGUzL
pVqBohWpFeOkqrGHGTM0ehSI5/xZN7CWvIaB234Hv3q0hii6jBy5eX9WyTOHKzmqZqz2QtLPaEhs
+IafV1seIsr3bD8XYgd87/47/DW0pukBsXSBwGw/P95xgGeE4FKimVlSHvLp296fJR33OudRoovs
JMDDXJpH2LwnFJ/oEZPy06Sc5ZXx8IHpa5EbIw6IGqOsWE0aBeXXNqMAi7Et6cXOqKDS9UjhO5im
Ak0F5eHxxxNOvHOktY9oVwBqtK+vSD4nblzHHQOKg6ovRFdI3gZHr8hlp2jurrM9synFnPm8+QyO
gHNwd1rz2mjNIuh4K2Rnwim2Kfbuur0QwgyuGk4L01UJK1eyyK7YLhRXVLAfdJmTQeaRI3nDasT4
XQnJHdeJOLYdIrJ13ZWKNLxY/nxEFGFwSWgb2iv1dMlru4OyIvPQ3ue2rqWn984U5IJKOO48rFCu
/xV2BUE5ss8hQdqcF2Gnm02g2GipflsYnJGQMo710iRwDy2L+0CgQUU2LpdmWza93JhUNkOq9A3v
XD7DBST4sNL+L3fnqmCxUegRIaPwDhRljZWcYD7Bfvlz80G1vKX2WyhPPlH24KCb1JR1Vkl7pbnE
rZn5t61dbwwQhMYvNzR90h0MCEkrkDTNAnT3EIwGNyl2BS6Y8yPXcVeLAVrhOrIChDy8If9rkImv
rSiO0O+TafsejweMpK/AHFMrr+WmB0gZcC+9s9MK/qlcK1w8HNRHj+J3RkS8RTkgpsyUfrNsWhFl
N0VaZ3mM1GsJPLebNLXh+IFxkVqGK6ARPFUXhD8Epwh1+VJ10c2kfMFtEXrm9L0MXs+xMS5eXNow
ciu6uJKtlA1ItzD9YSzxVNwJcgAse03Vkf1pld13jY99HBn4+M891ohhhup9qKzP+w7ogUrjY/ml
zprCXF5htZoP0kQdvlNJJVFo9gYB6eZO2cU8xUvWnrDjMn7MHapKFAg+JKpo1OJOGN4nqcid0dIf
tyTOgrjhsjuYhtzqamgxMqzagmH2i5cymjE89YhfA6mLP6d8vdaW3wZQI4Yuh1Idb455vMrxmV9l
SK0t9qJLB80m1NoNYO75fh4g0W0N0fFxOBbyrxMRKcUGFB8sx0NDoG/S5EsOYPlhPjAwnbm6homq
VTX8LnDfsRvFsZYLT1eUV18/HhtHSpXI5WzOfKEgkXwKPpiTaANe/tnTt/JcG7hSEJUrT4HwlVZN
peDR7gsWEPSZxFwdSbnDjSB5OzLb3I3pU/yuyGD0XbBLuJu0m4mCvpOjvRDJrCA8UbRj/ApQmvyH
1XpX+F/NZVatjCgBRpWK1iBvMoJ1EUxXzRgu1accmqDnceIX4QR36kAbFCTpLxDa7z9aP/aYt0z4
OYjXgrIs61IeCOr0D+KvtV3Qju4B5iFDrVKAbToq0ywGsAPh5+6EDRDNCbozE+6KQ7J/51VcjQFC
ELrCipm2QJJ/D5aJ+PQoPLXizeCgm75/0Wmz3KpBlRvlTnxbqR74hjx3fXHJbFcQdTTqDiXCUO8B
E15TcjhVN0eZ85ZaXUEkwGDSDOZkuHKXCRste88QKhVTqCzjLyFJHNKU62ZbLfSBbOXT9AvFW4vs
/+SsgjiPI34cIe85pE0bdgE4nHzQy7ZOVr99wMkW0Gn63+NhcEUDmIdOTxkAihvYz9qOpLuV636Z
98GGWZTs2fTJnMs6hqiUvszzj6r3cgsnVx8SiCkBCUHmMckQIpOxYR2dpvK3AbH4nOmpEg9ZWk1B
PuKVWWDmQnW1dQLczoo52lqGWail6nMM091LBXWuEmUw6LtVLyKOHzOlunjt1EIJ6q3X5ScOuzJo
vrmrRcSrphiqHv083SsBQPlejrjyq2RWZTFiboxiVBkAtXIy4v1N5kEMwsR0xBXufLPnnfjTxNPs
D3ih/8h00zUplbY/bNaIMlbkvrt4x7LVOJ5jQqAYD1CBecxIPnMYQDWYDrdLlioNKHHuCD+F34hZ
ua8n+t/Kamu69EPTY6bdZ6+4Jp2SiuAyrvQrEVZcIKQ8yrxYUQB10TxJNtHD1jKe7Q9v831d2L5b
7rKAX6jv2e5621XhWA3PyIorxKixduwMFONS1KS3EzmINcbor3T+eVw5J3QqAlcQrNpJIWBW2dP6
sh8ZuhXBH0I2cXCkF1/+Ul1ifzKkDUI4pDovHNACI41rttjccDcQhClf0W+LjYRbxkRBFjtz5Z4g
QdazbY+nGNXJDnCyC2FyiqVUbHsnqof1d0+6pAEMPYQ8sHAjKNdcponudy8RSaaeq5idWnIRw4C0
PJvV54bwqvPGvV9JPna5HmQX+eO3fPohDvtYzegFLOWXcnjL/ddC15Be1Ta8AqThc3mDrjRILa9y
UlcmMxrBpimtnb73GkCIfzBq6RHQyiMNL3EvbSlqbYVwOcRMNsESTtId2IBNaw6JvO8i4Bi8fOZN
lWOVQYWVBiHXIgjzEEX0KhoNBuUqYLvcXPgMwR+huis2W5c/9sn1npzEXSseDxHryWPxSTOMaj+i
bngrDapZ25GdCzDX+Dzwbg62EIdXyPP0iwOJlHRoFxoPPyvl4e7P5pe+jlZf4yCK9x5O53V4w6yG
46aNQziJhZnPDfIRmCL9FV/3w+holHYVzq7KgkH/oFb+9Rjrih72obHnJnwip7hCFyNIftLiJRsk
l0ol6Z5V3x/u6AbAIO0/aYEJy56/gzK+2sq9Gj6wlqJKGQUUNllw/LXLWksIWvgbFGngtfOp72gW
aF/pA5J72tuDDvSYmH44AIu+YqCIQgNn8RKSqp1aXI5Pg2vOQ5dIuaQOOjsXMG5PQ+MDzrd12lF7
DzOc0ho8yiTyjaE7LZoV0z+k+EZxzt749jwVxTnHPoqfYnZ3L9Oh723ceTy5e/rEzaOYF5K2o0ZA
H6ImySUFlt7BpB6zlJYRE0dD3MbvlTwFGKByj5rJZJBgCCUqHa3+T9uWi2PcCMIRo41E9rstJNWH
9fBQzQ1mOCcMA4gIZw7HhHm9XbPxq5Vo2flRJsW7IlpngoyOjSr2ZNEkL1vxje76/2XMErg0eiv0
UFxCINMnmhz6aHNm+KXhTH14kzUCP3juck87FSJHfTrRDBNXegAaP7jOrrFkg7KVtOTOGoLZTesi
CJevcH31mPFg1EO1gQ/4koRDRgrvfDkqlwS1AdZFccycq616bUZbsCgYXiiz/QDjsGqTvXSHq21v
GGjmzyCqpRCf6L350FHIxuEwhBHYYDF54Jj3wMnzcT4KBQ8xx/3cZby8rxfuM9NPtSFqAfQ+8lrU
HN5I4oToSMV8L68am44TargsQP5KW/ZNW2r89f42fkn1XZCfCbn+xXPYIxEuyl/BuqKjPAS87G+e
/7Lj1rtElnf8R6nCq1QXvy7qMfPgLngB8M0hZIkjhpqr7rC97Hs9l7wzVEFvJslTyqCRJ8Uxd4FB
xI8HekBwpvrVsmXL/GkGYptO/C8xzLM9jifynfGTeKQ5pxzz9hWE3gAf2UdDfJfAOMutUpwrvk7h
m1tBLvqwx6vtK5KxLNdbtUAP2m6NYPoZtFznUtHUXaQ5jBj3BWwkYYbgk/+3b1XyxPwTlqXnfol9
MbJN+4v6+3t8YgduHgjqCqFbhxfU1NdPvsRASCmTpIpxlv1BebF6BSX9/zRlV6r4ruqi7hcxWbit
8NY39DPDZ9Ma/kKaLIc4QrY0UdJjERoqCzqvoKr4mJ/mM3zI4VGKnLVQlnksfcAewgGz4cPFc2bW
d0SVuslGPi0bXSpk2dBQAG4Bp6oSAAUhhfwYRslH0nwWnpXcqQMlo06gSXW2KSmDlZwjqHgtYfku
/b6Iadw0kXCaOyVdCJAMELlJcC4vm6TZWMpf9jIqejOPpAT9wCzM5HVyFaLXAAsKRQRwxlms7X7+
bVlkH/n1uyJ+ynW999iwb18lpEqsvIAwOgL2clFwV0V12SrrFcgZ13MXKH7+Tm7cGIQyxfOyaUY2
bMedhzUOxG2Acyr72GPBdkc/OtSc+SoJx77/S0EskB/f/rxEVrc9reKjvyWGWQnYsysN8BFDatCW
O+mBT8mVvUKWAP7CG8CezWcLj1kfmKVurePVS25zr95jRtHzykddFrlaMHwg3wmqCK55z+qiFOn4
HDs2OmugewIWxCE1DPRdJHRuHxWCwExXgMFMAGCBWBHJbauKjqHzfaEF6QsQ3CffV4BUujq6I1mI
xOlZb58Hk061ifVBH9CbHF7Am55JW/vjV4srFGejXJ0aj+wreKRUs/l0y5asaaTd+h68z7UU0feC
7QR3Toe5iGYemCrsuUsJFmIIeXGtyr6sgaM/8Im1rRgd5b/+LKTidJs9ST280XTicNAVUx3IdO6h
ZWomgi7V+m4l9myE/fny6Kv1x0qXuRqKrBu/pv2cemjyzQpP86Ped6KKLL2aGmpis/P7hcS0RFol
EJLro2RBwPKG0G+gc/ETEMlLNoDBtMzvlRQS8XgQsN8W24v9UVkn/tN8I0DGRLbWZd/5DqPcZ8Kw
dqNxPSWXP7GaoCszQ4Xa0nw4eoHCVg3hQFSOdZK2br4lLsdV2wQho+n16CASz0a2VPB8yUpLMitH
u0bGOSFmBDtXfHhOHgMC0rh3CZLUimGofXz4LFCnz/GtYkwSebrZpfn++hJ3kX//J+brVBS58dLq
n+2FpTlVAoJEFYuq/7xH/4fvhmkjwrO1UXx2LMEPvU6j74viNm4RND5XJzdOMUMeYaHJze5ZkYbU
54gwi54t5/9Le6bky5HRhQL7RNtGK08ct/GWJE4BPQ3BIE5LvRfsKfrLsrKHfKmVb5u8tSgil1/v
MA2I/4S8RxAJsZ6tc61HUiESktvbquHwsp7rU7VwkaqTW6xZLhT0nShcjfpgxRPgpLiqktuhgLgI
QTdfHO+T6ml6VBcRA8yOxV3GxC+SR4Z8Im05tdJahg2QGkJtyve+1y2YeRbu+FbYWrScwFNMfPaM
YGV7XsGaZTcr1pAQ7YSO5znB6pBpXEYD9jC1frj89LgOrOUvFkBORba1bJJ20uRZTKWrAYrFtR0F
qOzY1QHFskU5FZoP63Mts8FE/kRBlEPU69XPDl/bBSFn8YYbpfC633fAjcKrRgBAgzkhavmGYwjB
kLluuGYgUAruQivGfCoxyTSPEojgd5sRjyI3dIZuIAevZqxUUSmAw+yWKDTTZl8FPuklLVn3YoMo
IA+ZsjnK0q+rThs7+79pCfEVN6rFqheMAlo39WrCPkywHPbfewMpPo1FV/rZidhtDBipgyCujtD0
SkhULJvWbbO83YXLBmLk1axdYY1xBZ5UWgXC/NxmbbMnjQu+8ULCqtdWIsxVXN6/Jcu8mm34rdRi
5wrGCQ4ivRXuj0/8Aoxg/7vg0pcvisefkJb8NKOxnP9D0mXLN2B5i5eNUH6/iZxcptHlCwwdcw+C
UUvyblel2t3q9DPjukpGny3WwczSBZYmc3gLR7sV13mqjJjsnXChkyotugW//Z3dUru3AWApSDTT
KD8SNkR8/DjpcLZy3hPDdOzORu+rmsF4X3OOXnVbwp9g4f0qevYLCkavId/x025iDgajkMbsJaRV
2nh5dnmTVr7PunI5sARuAwUV+4Q+RIl2b4jDtcvPaGwCVkP58gD3w+0NNwCh22PLa+bzU13ysyp0
5IJh7/Ztr9WP7796bIblLZXIH0ju5CCyFPxOtslESoKI76Kre+cf6Icx3yJ6wTrN+hstYdKQKIQ3
FwpbHC9XzGCn/YqutOyJixLJcy4IrIKb4GVDhNLlUnBu6YgHHnKkE4NJ/oGiA9yyukZBE2gE3P93
4XRF2QBOnEl+2N0xmI7d7I1veHM9smgCZFBptJSzYKV2glvUO54zYgOT4Db0CIEcDrXEUOT1hrif
XCiGf4wC4PotzUONJRuMm5O8OgOdW+mPDuzbuzv38ei8lFRlYVt1sDnFFj2BHMXhTa6w7Rx2BtGG
dMxy9BuhskztJTnbEPHX2QWooxexXp28utSvoozPB2Xht08s9rd7meNPhFyFzwiEAv2U1JkBP43C
VDykB9D4HctKyzJ/jbclWslJUgLjNcpjClv7Mkowf9ZxwwcQdTqKpTX16+jzz2QeZtJS3OLgIwrO
1Uzeycn/N1IjF8rn0/NXrMckoytRyYQULspM8yfk56MzDnuFpqe7vP9CsOstvRv99DyKmXkUYMwi
EWqhyA/YcosNjBSnPWaUHb5z6BEiU0WOEJkHl8Js12sBNErbPXq7zg14f8qv5ydUs4UWXeNCeYFb
O9PM1nYoIEk4OzGgZnSuz5tEXqtKZgNpZLbv5m6r9JFGP6V/LzqRiYXRUzysUXhGQY0/tELOb39H
ng04K3n5FMGsGLPQL9O67XnKwy3DXzuvGGmnTAMmSvkK3Gvbrf8lfhST2bLL8Wl+yNb+Ky8ja476
A0+dWJsDkyxk8iiYZMm94rr1dZHwevrX3BBabV38aRjEwdonUnjhxG6S7GXR5ju9LddxyxLpwf4Q
R003aTy/zfaPRWOsG5zX1N5tGRRLLbqDhNjobqEKOR+v7rFGwSj4PW/VObkYfx/g+TDb2n5VPtse
QR5+c+sFW3lZmDx5kFxv7DFadz4kdKJ9JkCkkFbrpQ/hh0GALT7PApAqlUqmDcamUPzYVLLtyXS/
tW6u6PUhe5V4ChDjE4JZFf+bqekgp5O5YmZ19COh/Q5WmfqTDAsTI/GjN6GqBR/xTTM7YvoibKFF
5R4sLTFG1G6+Ijaf9/22fhmp+B3V9Pq72fBh8a+Dr0yBzwl2Mu4QzDGvAMhJ2N2UEI8cotNUay0S
QYTSK7fQr05cd+ZQ1te4GWAUjttx1SLYAfpkn84OMDuU6fm7l/NywHX3vNZh7eoy6064xRkusHeF
I2vhV7M/1FDkGDNPK5igrMdUHlZ6y0gD2HR+jI0n+q/3qq2guMD1klIjleNDsReDtdhQ/76mBXAK
mw9teRnJFxuddV7ZvH4dOV6lfZK+byy+d/3y/CoAl1PjgjDyEaUmIqX94nR7ujizNVuzNmZn7R9H
hELxNmJrA0I42K/2qifLSe7YrlotthiLQONTkwBV78/DTxzwYBnXFxAdJfbG0Yk26EdjCds/FcHN
aiP+OtV4wPurmz5/pEAFDeUEesIQnVNy4g2uduRxKIodlUSiyEGAf301LWD4g6BFH5+ILqpbxFmE
GFxsu+8sjCRX7/d6lg5lyzcEm557PsUWJWi4a8ksdw6R6ES0JEBCPkXJ8FMEeaxujOoos0a2xdG2
9cINjZkZH81sKoLo4Dy0yDKYBwLrMUOQi5cL+NdT5ZkXowyaOBrfbQcr4o++/t/294JA5uxxlH4a
QE/t8lPIXmiqCVHPY8OaQWX5xSJWTfpDdBa0NfSWdKF2XvvR7AfQUQqGLWa76qwEkIoERplgcweQ
7qeA8IbfzF8E2+feD2Hh8DT6/Kj/LolXRscY1voc2LVRW6/Wo+VZaPLXNwng9wh8xBDAMRpWZeLd
1kS9YfetTj41E1yDGwdfkNMPCcQv8oagVk7fJdpeOWrq34XFEbx5nAj+gQNonjSXkmc8wimCDt/T
LZBWlrMZPk9T1pzi5Epr4J5n+2HBy7zOgvXqaRn9FBvV1LQC4HZpIHzfSfmjweEZtWZKfU4F15qA
XTkvMY0zORCS0cOVT6EXo5qscHkFFu48mDBN8UmvNPs9K7VH3JXQJUzkTWggWJLUETZLC8RtmOeB
5vt2wunQl4LtZNdV0doZ1fsNlPPZD9D8UwEj2dkFFX5V+w0T1+SE4ofSEJW4SoBpJcwbzey6Zv84
EWSmAiFaGCpRbLaz9ST1prmg7qyzhlsfMc3LuBsmKf59GwbNPJvNFsjIjCmKf5QGq2BFLkz7RCcx
2ySShiQP8Eyy/LKf+VNNCgjCgW/lL74kklfPfFkulYomTL6R3MSyrGKg2Gp5PwrPnSYe0shEDKQl
H6ilT8Nj3hSpjh6o8e4RgNGom9MGR2wekckBDUHLknmUJKnH2a62esLDKqplXuOnCdZabXrhqHii
Uv4DWNFTD2e5dOL8BANaK1BNqFmyfZR5vTUCAyvYtRM8RD58pLR7r6y5W7FCp16+sg0BvOMryzcT
IRPlSeQ8Fot16FfU1w7BT718h/0fDvzKmtdPEp7fO1112Pxmbk3oqZ22ASQXcJzgMZuP/NQTWaSH
bpn0UQKYHIngikoM/7lIdVtIi/2B2NSarcUnX7QeVskvbm0tu9nBrrqvQIWdC9KSKjsc0fOLuZfq
cMl8WJhyyT54o8exyjdNeqe4aoKurHkuH8ptfoW7ktZ4sonGz5tE8k7nGlXCc0tBBejG4IY10A+5
45X2T5GetEyWbMHTFJ4Ykk2YoEmjV66FENTJomsrOiqrPL27vWm/QdxJgslNeGcVpJAwDkKqo+QE
I90+1EIFjNaLe9mzVkaeGxfB2P6PUhJL/aWLGNwgMcqZX17hHI+2lZKPTiLbnZPU2j6eBbAvg8Mn
deAOq+X/7o5mhujIzMqSiG8LnilzoMNnCmlak8hXyFXN9l+LDvJsOGXPqgangw6T8mKzNunGG2vK
Z8KA+FOYflggPLNM9SRucGNndycGH8EjtytRa1xqQfKcQzgQ5cqFjplSSDUyfj3boFHLnfhlotJd
20alFxQXtYuOJzGYLsslthnmoAJTpAQJEMnpc30jFq8Mh944UU5rQg54X0UyuUr4vfSjP1Qqa09A
GhpbBP/f51rxqKVw3szgS5v3h9HBQP9ZOXHYyxCiA7DqIQc0IO52yvt3HlPuLEWJPIW8jx+sr1Dg
ZhbdM9FU/d1KsEYLZI7xFSOSRcrV/fuZBSXktEydI/oti/v0OkSW0DVb7VQ9gCeixcRhJHY6rtta
6J1qZrQT3wot2AeGwZOk1GQ1aD/Lv5A44kVUeNX2Tc3UyGs6UALD4ewZaAvovkUNCCJSW8ExrQ/0
mseb5fCTfmZF/h9GoB6FRc82hWLbLO7aN+QVy+Hx8k6y07mQ0Op3AfmFgGwT5pRqO36amZmIWneb
yvWntlfs5Ae54NzMz1om0eksQgOLt0p99gDHvr7sBZ2WSucOsUlUmrrFz1ixJ0d7jH97kgkzBwww
uW6bwBnWISE7dNn2BMcWu090J8/ao4MkLtesEtGrU+GU7offG1DHJGBdGpEeHdJ9Ded39JWJW5Vy
ZErF9IGZcJl/scb1F09bpd1x16hc+F2ftAVg3bhGqpmyCFZkcuPWT4ZCIQlHHqisnmrHQ+Tmjso5
cIqNciklFVkSp0jVVVOX/gEIZEiwkV1ke6Ar3jQ6NaMrjclpFrrBSIaDTTk7kNIthbLiNNN8x7vv
G6OKhW+Nx62RJ9bD4/8tyP3fGBL3pUMNE/65pVgocc5Pgh0zkOveOoO3Ob/u3KBC4BBW+n1AmWT0
MCiC1nJMYuZvJJCbQ4bCrfgOCRCvpTYUOhJ7EFH4EohLTwSnqVkLoRdaTyGBhfzYoVCFfMkqawov
qO6N76E4z2DHjSWCvXwYgU3z+aEyWU/DCsbBre+OyPInbPPnTWneh48a6075yyHQTyHVGiy61cUg
P9pQWpgZWt2670epANjL27wHxI//b6AuqWxtwEZIFoN9k96oTS67kmwZRbsVxFB9RaSMgl4Fnfok
xK9vasWzzUiWW9TZuGnjvhHVSP4Zcrhwfo93gVuOukrxyqeSTHwqeYE33dIZ+V2lquI0k4FLhnc7
coxXlOoAejDq8bCtCQ1XcwWy5PrAzPNEQQ5PO2brNGW+H9pk6BRXvpW88vnVsLmiRxCMr99KjvAM
WusQIwZ7SJGPyefElmFoEpkNDpPL04SjvMT2APxLbHaJz30VPbgulwkgthtkd3zTNpPSWwOGR+/r
n7mJzywM0nwZr7hQACgaw6eHcnaFQcd8Cki0+9t4hTY3eAdfPAK2Sizdzyncfn1UwdTH4bvaGAz8
QOeAwoX++Rve6JmmdzevRtmk5jqJqiCK/EVs33UsL/U6MSbkgtXlGlDOq8sqoTBi29rNnTHJj1l8
FaGDN3abv8h639mX5sJM3oGPKrQZ2KtUVVqcx4WjLz/q8MbqUD3H2EZbQyX66ZFQeOdSmT39l4Op
k2lY2njKPqXWDUWyawBVYEavgGWrGmxjc5ZHFJOjVuX0AJDzCvsbzcHElO8ht1fPNwaNoD+pgeTa
7tlgTMc1caKyuoymiRNrLjsyTyn83R9TIRkLtKWl+NLpNMIJwCa33l1hlnTxRJFtBYqH1Xn7lkhX
ytyJq58fKOdAHJ9XlngTQv5TamStd2OKK3xzgFcdO5AGDz5ztaBgtMUUOKueU4Hh4ddjA4zHJBmW
GpslhG5RZVnZ391INXzhkR4zT0pVegR/D4sun0BphxbE8+PPeDRvKHqvVFgJGWSHHF9ILibW8IAB
ZCLRyt3GemLHA+Reqc58eNt3QLrOxRcNyAOKM53zgItVw6/AxYaLXYN4rjc72csAXaSA8CLJ3NHp
uEZpVzDcuR6yIf+tvnzm8KF+RQWovD7xqhvGXDs3yC0BkQ4EJfla2hQVqZ0VIDZEovlxfWVHCokg
kx+mi2aqJZdp/V0ZSieCYY8Z+h/EHH7tB6tT+zmg0FpEkHoTPv3bv2KBrX+i2/DVt/yK/SaVfit0
BR4PGvOxO01tjNXBdCCDTh/Fo8EF1xJyAHrsPkY5BF37bxBh69WtS952IR8eoSSUDijQe4h3Wexs
m5ZonPndj3OYhWQM7842WDarG4LDG0bCjK4L7YQoOZqOwqw+4dM/AJEds1qmt/jFcKF+bm2D4L7T
yG2qv3V1JCXUFcagvLR0uHL0ZazMZx2buw4Gk7WMHbMR6lewFSyz7e8zgbcd59uiGmydZyP1CF8H
Tl5kB3sedeTQFp1ROYt94kw1bSSBKWQaOPPyes+X2Jo2Jt++vnE9XjuI2UjRS/n8nrvXDB/FPs7e
I3iXy5UurYdzF7OvRUQLAbXL+iK3jF9hSTxiZgeV3ZEcXmeCO2DEQVQBhbQ15S41qZqFDlXf2jGb
vyV8YjXiDP+WoaY4SOmAcdjyX7fsOZ2rtptgQMkSoez0Jq/KgEUePiPAGlQ/D8qAtOGgzQSsXeJj
Vv0OqQcBdeCJXdsIZdgdhWupspDzxnhxX1h73tXjZ3ghR3GY2Vpb1j8cmb4r8XZevS9sIQuDDH3f
IICzpNXva/iRQEFgI1ZnwdIorO+Nj2HYcqZWwvL61kU+VMjAQlUQRxZY0fciLWvjXpfUtPaf4Dps
GE4j/v5qTXIpMS6by5H52kmNU18HirxHjlPgVrxTcdSsdpMr0nma0WbfwAuwyP2drEYNxJ8BoTGy
2mdXFCWWGHTsIC8MLW5syf16TLsXkfbSO84aD3Kc/7QSKykh4yZTRrpjIvtrN/Z9O+R79vpLQ1S+
iToUgGYv+KjTZvmeqASlacmk7VR7TP7mkr7mQlhBuriu/I/hDyf4zWHsVXNRDoiU5UgtiLXVrMh8
HeUGrZXE6I2pl9VqAxAsCd96deb30AsTd3wlo1XQ534Fl1T1A8tvUIpc4gmljBaEPrv5S1VKMuA5
xjsKMVTrHNmxNQx7FB02ooittGF6c6mDzvrnTvYf4V6fKoB4weS5Tas20Y+8aWEYCNLWJrM9UdDZ
WBsM5xXAvPgO0xGAZD3cEk6nQPxIS/sE5i9RmodOmOUCHoSIPqvYFesVdzlcdUznkY640OC16io2
QV7wn5yEqwFkOnxAJDnWKj5kYJA/Y5JX0XnYM1zPOeP77LkgkiaLiZdE0anf4QHEfnpgPDGwTeRt
ortpeR97jWB3XWL3Wwpp4Tr9n62wwaj/3lEoFdehc6zanXL8ITyywDUBbppdHS+NOyOa0jJcBNUg
Yd5gQ2X9imWYUvKXYmTX8v4Q7gzCTTbY+xXpHYo/pcnM90FqEOC8GWLxkM0H0ETgnukaXba4rcX4
faw5OnPcIj0bLnLPkfzvcehYssBmIXAzVJkrVBaUnuJz36MCBIjay6L4tSWt2QzR5D+Xqah08tSM
NDdNT8BQKJCh+eMf4lF4jks0iE80P8l0LQf21gu+ENa58t2PGyvXWdYutk3emSKu+lvfxZ3VfP3B
OXLdclQKVMtY3o4kgMmMHjhV+vxrrSoKxCC5xK8LxOKPa/aNflx7ddE/NtUyuMKM77jihpUqZP4U
uJb/3RY3ZHfrxf7HZVAATlE6moVhHORsT4I6MDxoHKWM8xXrmcUN9/roU7w0DC3eB64xFkq7s4nC
W6Dz7/TcJAKa2DlNcXRqbKfLmce+VGJZU+yxORYkhp7oN6xE8fbHgNgMTc5S+GtkY/9V7c5QJFlj
pDGklBvPuHjjAwBk0sZ8GBEALDFzdM152U5bQc2lmNl7PHcCUDYt/9KsSeTmuLaRnMlKSpsM0tvN
53QA+vFR42XYntB9NAdo44tOF5HLnL8C6jcuO3hFiAmHVz8+NW7b5v7MBtB/UKjBbmVU36c18jvA
K3283W2VNHrt1AzcV0DCzyRp1dvEK6DYevoIWgsHNXXAe+D6AtFe3rJ9vDDVdHYL5B65GOEj7Wal
mujMK58iJK1zyZfNpf3ATMLOoUN19jihqTbqeriq7hYS2ZlnjyMhFV9F6QiT8cH5OAVF7K5Y4YSB
Zu5W0hJlW6PgCC5DTtNAKdGA0JTkLh++TFELoXFiFJjSBXWHix4Bb6c6egRQ4FQ4PuRKrFPON0TL
Qwpp/tvRU0vErFiqAAgVOnCjVxSgUU/XxcJZm1hm52Te16wbAceVHhGiwVDD1gypEuNg7GGfo2JF
fcoe8Y4qz36P/7yMkTbR1pGJGiJy19OrkXx7AzoNvRCxDGKeXhpoOuyZXvRCHaQAJUMjHLosMr5z
1R5IXg9NvojyIKkX65CwJsnupzIxTaDCHFabzX+oOvEpfa3QMHiRxX5ToXxlpEvJ+m5P+LMBY2YK
rlZp+NtrShHMSGW4F4xm/2Dnu2M0NvalSERsIFR2Ve4DIxHXjYSpEnjcTAfC5edlklBR9iBM+RuD
AVYu10HviI3t6qmZrQ2wj6e0mjq/W0PDoo5I0TO3IoWymtdcqC8UwNZjBqRqo4ZyjeiYWaVptYsW
KW/fGzPzc6qkGiBys0gvRnUfl2nu8/Tz5sax2CRVJ+brAFHJvrL41xtMqxJuYM2dmWQXX3CsLWTe
aSdwXnqSC4h7/tUVoutHlmQToiO3OnO8w427C8DXOA3ZSEfHvh/uAsy/21PcGZ9n+QytCVVCFRDP
2rYZRcTKwIspBOGiNmtiri/HUlWgytM2D0ELN0A4QlfbMIkoMHIcJ3V8DD2OXhCp5oMjjF99Zqxl
QejxTga/hdX0AvnvFPgO9qC++Tf+GVtPrWuzK5gLAVV4tg3JbhCCC2E9JDydl1tg23rjtido+nQ0
wYrvfdib7KqTsvaEwCcwj6il8aTvFHkjYaoyoE19qLiCO/cCweSRkS0Bka61cMHJUk90tPznQ30y
gMmsCy+HZNo2rLYWHwqZ5jAaR7RwsXNy08BwbtoIKt7k5U7aAL56Wn2TtFEmyS3zgHDAtkhfeQqb
kQQ3mxAaI6JKZxgS4b8WDUHKOU11dgFqYsEHdhYU0pO19q8nREkPMqUQuXBYjT/FyK8440bex+DG
Uczyq779EVvuComkuD07KoUpOvKkxkSb1T+WW7HGIqyyclTV+ZM1QYW+i5fun+QL/10mHuexmkJ/
yrENBMbzH2V8cEue1Nsspikn+0e/AP4R1qso7EEQblZZSoneztAm4xG8mkAHjUQclRSnf4tX36xt
HO6L6DJtrowKY1WkqUlk5Z5PlTfLP0aGiKMV+p0RockoRnUO2u/384bmxNorfq4MFm5CE17pTBZn
DgW7JhTzL/7cCgwsf+7or/yeSw5Qly6UmldLC6h0p1Al58RyDSehxsA54gxPSKu/VduyBnOd2XCy
h/gf/MMbNfBKk4veyqQ3sy1m8bun6Q6sY81ZfMaZuNastFVlKUjT3hXVlPxyI8JynwSurNzH7zGR
6TPe2mIcuBrvFs6xbAMdz/CrXNRmyMVLwfttw5ekTyW89hvkZEwFZiPNWlVDgXZQgUz+Enwv8qp6
zL7/G31+a576+7uGLPVeYA8lry4q4rvr1OtXuOtuMKEHWqFDBECpicyMVGFkdyxWJG8aWRfkdUyM
q6a/PXAKL9G/kQe5zzSYYAdse1Lh7Wjhpg/Nc3dphmnfy1QATT5UHjUhtL7+C4+9CZiDvuxyyfvW
7RYlHYcFvfIFLGB18aRUcmoCssvu8h4hvdPCqt4TfxHZU7IHebWQHRvHYl70R0P1yNaBt9PCVtmC
jWjP6FUPncHjr5iokEpeUrVJSOKhIjEVbOixuKYt4psD4ihL6CGBGXN8/as8csmA40Kk8e0JuM3k
7PekEcGpYNJEWHVTHaScYBfP0lRc3C4hQ6rTWHyGZ7wRFLjSjk4QEz3f3IA3/EzmJmRm2nqo+dg0
hZPpBJlBJv5Z9Oqo8SiH6bUfHR94yiXg7fp7EQtcoG9hWwtqra/hh9y2LgtvnOkYHKf0mVxMr0eN
+yCG5qP5kOGP1U/HI4GQ/gPEdG6I2qopACSURPlMpmV1dKfLFtx+1uSFjlx2xJkuOkrCW9APuZxW
zPfblB1Ytuzde6W+JJX8Wxv2ahOaq/8nlQrC9cKcAdqm4FfOOq1ygkXw/zE9JqPSXLMn7FyLGRQK
qeBMNBqR45tPAFHNvnwUKWjsOCHRbKm4iABC24IYPLyrEZgxji7wtieI7T23XMHQgaptLcvJYdBK
Jp7FL0iGZNkPgXMiF2MkiQ3f8x0feuRHlDF9T5BDHf3pbfWdxTb/od+H3DfH9d9j19z7yueUqAwH
S9NFPKMY9akGWUzNJv5iJ6yOx5AsS19cww8yKNHucSFQw/J4Y2n0e+TpvDKq3FVkNvrWDYSMow+L
UpSxkKFGMLXuA/kcqGBho8EadBobeGpjWHvBSuzrFN1eFFpp4hWI9WwEQ5W9ffD1VPaCiLnhWWZT
AKviEvN/XULBb5E3qmzjtAAG//7prF/6phLOdCeioD7FfGujJGdul6Ep3DhgWeJlTOw+NXz+IA8i
93CBiRV+vjPkYrLeMuDnl6PLoVRU+thhYMJkvD/EjYTjmMsVubkxxLGMgaMgghhMKlEkrRdde0r6
WIQmrvT7bWo8ol16oEyi/oyLYnx2AdsJZlxze0vi/hTtca0kTR07PxB1ERPbKQ/wl8qcu5CaNHzS
svNjyocWQsCb5uCkPWwdgxz5t4Nrvcex2DM7BdB8nLV5wIZa+G+1fC0X0YezjjaD5xzRqZ8TMAgi
cbW2+kipLkllFZfHk/GRcsM5z3dfR9+7kClGshxPnPgXZ5vEgQt3f0XfLNL5JJDXKFPI2QFB5pcg
QZGNvoAbAics9HFYikz/HaxNgquvX8QsiA1LjxeKRmfGaPsYtholO+c/wJgyexRSD2QwIH3QXiCJ
fKxON7wMLflyXRcYDRIo1XaLbmcLH3iTOCtQT5CXLsEiiyWII+S34+fU5uqD/p+zwUEQC4Z2bIBJ
zuoSm2rrEsHCwXNHmB0+SHUwAuvRrrlZ/UK02TxFsAPROs3FIGQBR0BZjvN+J2pFqThw6bLUZTlx
PPajJFQRVqdmtu7n9puh5jRDT6MI/xDggsW0tzuPcoOct74jV1Q4Kbx5HJsgtcCUzpkr0XUryRsu
n8IjmJZGjb5k6v09kH6KhuJ5ltrzJZeZQP90YuqqrWwt8oFI49O3zzf2JqBsFPIlrDtWHaPqcdTJ
qM9TVPI+VACxyRv78QS9duho3M9nocROO0YdgH3xCJj4pCkwwm6m5Sxt0bAQMRIK8jfpQqAeGkDp
3TZxeGyOgPAfXzPSSG7ruSx5yT0yp6t+izC2JUhQXumWCqkkrvuUSrveV+3fLGbp+4VTywdJo7tC
q6L+kYe1l5lfZpQdN0akwhn9m5quccB7utklkW9Q78xgQXX2Pjl7DbsIMg3FoX11dGs2NFrvaRCJ
KxXZGDlVH9W+DdZey7ELxfR8903WwcQHVKBx/dlq7JkOL+VeU8kt2KkpFZF/fZxX8gCufpJoT/Bc
/0D1hgARyeSAE040xpqtXXVY+WVzXrRn+V6Y0kINtgrl7LwaaphFT+f5h6OcnmyRs8uaMp4Je7sA
xFk2WTjooU/2PkPy025x+ADh4zpVZix9QHhQpAl/zV85vxHLIzfd7bap05WazwIQP0SpVQ/JajR2
zlnGYL87ub9atNl2GXbihGOWxGjNQxgk5QIq4cG0PqKWuNcYeawVHoyJVwuZ0N6ACeFntfb4Wrqe
aRqSHol9l1BTGdyyg5+qMibwhlOGWt/pdDxNDi4qgvkqBehnkn77XxnS4TQp2nkA1cs+7B086CUt
aIaV3bRneU/shF+ehVRkxbNn8u2MEmb5YoEs2nIvaaK1GUOyxJJBmer4WZzWk4bl/7aGmKTTMoni
2BCBk37L7tETWYXcnrCmBCB/gTolxyxp+AASck/Yd4s4VbcqAm0HHKwP7aaeZCFk4t/OIfbncbiq
B3CFChUsbBmus1ybhlML7Swq4UwHy43Wg8Hmb+yRdkaqexSACYUWyleJcHs0a4HE+dhyEWUEkQSN
g0Dn01o0NJB/cDRCbY+5bH5v2+Pil4vx/dq2gNQWpr7r0+TTYtQkAFbwGBwSuo3gVFy5PrT2dk9t
8WAkjcVQ5aisXAc3GV1MvJ5dDoPpIr1fCtHp3NJBOsc8jq9t6RcpkV0Z0y/zoY29uTWcHMQa8T96
K0Yo+vRP9tLgnbkVTwqdQodBzRC53hRld8GiDrXzccG34nZy9yz2ZDY3/kvW914csDg/HrXuKHqJ
ctxKMd0o4lnO1pYqcuBDH13AKSag3onQR6X2LffJBshDfkEo1zeg3o9xnnOwZuTxwLx0gxx93hF+
EuYSMEu+4Ijl7uviZ+MDujdM/IrWCSPeu2xF2vbdazwtT0K9dPQbWnKZjC7stKI+QelDjLYjx7xe
HXlyP34Yre29mduSWcEwXVQ+DDklv61+HmxPwHBcQD9o6G0Ies3HbG5/hcOeUzMEoM65rtPlAvDG
LXLq0RjeZTn5ebk2E1hInuN+f9UZPAL0sZ+zfVtmbJAEs+x6MhA90sr/VkUh9wVfq3ymnlVmPNyb
BCUgETH8S6iBkcZ2F54+PYSzKtC/1P6gqjPSBonogvX3ORn7FcDBsHyIu5BJK8MkzEJGdBCvtZqU
v7w8aFYEeVz9bkEw78C9jvTyHh1X3hN0M2GmowTrcxXTA/ND5u+Ih9knnTA6h44p0QAl6L1OiAOf
dECHcpnt5V1fCfzFzZY0I8udjltKpBA/AqirtH/9KGspEcWqjlU/WzuYAGKHgSjl/BSxIoYcNl0i
sQ5hCG70W0gP+mGjq+fEMHYmXB3PhKDT5jhSwmrg+qiT2pNqcWpjsMG5KbVqwbmqQVehpY79dQc8
ak2ICB2iIhgMKpw4mpvOxo3YEmi+uIdGcsgAOaZTfzqouLSt788GTYypvN1/5EkxuH5lXrTdxnFm
AG2rstewpAR6rXV+TeKzAAVfi7UV1WwyLcP9+vlnmQsAUU20pA6hcrL/Y7yb3OsGdwApHNaOLr6z
yXch+WmUpz9Ik+BFyh+ePsEVKZ9nX6y7BjEynvdeAhFuTf0G6CkJymZcsKBU05J2IFqlWZN/CDL4
8gHGtHRJwpPm3OgUoV2SJQJ03CDbo+zSn6EMY2uQM09RRCasg9IPNcLDARewE3Y+RONpwe/q9bAi
46lB9ZuVIE7bUhvL5pO/Zkf9AYIXzdlb3D6TqW1shcvGNEiLebD1NUwcI6dUAyeL+vB4nhnzZGhT
5gVcYmoxkMt4QVM+voZvjajDp6Y3depN/sJqAF6dh8nwJEU7IMFTuWnvnRDHS+z85lEaxaDCkG+c
41pnv6vQU4rI0nzXRuouMVw8HSXmFl+zzmcGCPf+BLSnCNLjmXAKMkRPiWo/YQw6NinKvBOSBTHH
TIJ1IisXmasHkm8buJRICv/GdKjg1Mn+fR1BWPs8Twko1pCKNBvpR0fAtP8NyPvE8XZyt+rqMX2g
UqGuWOJj43npIOI7gHOiA+EE2A5T5IxFlWolkzmImtjP7/22kjI5PazBuD/gJEljZpsTD2RJDCWA
W16fvHYQsCWP1dkoFo6Hjj3A/sK8GjKb8CrhG2nf3UtTeTztdkdlAXGpP5iD1KjJZrN9hIIOf2GI
r7euF1I6oLOFNaVbC14XsF/ZeJWKeAdnfgQBWXFCVkpGxx4cj90qlIbF7Lbea52j5Iz0I/lOI9+l
9wx0Exzrh/wV8uzmvXdLPESIncSeElg02aDRmRjmIJgN7is3/GAkn+ktVJHO1omfNFA3VM1h320Q
yBBr+FJNZjlJ1Cd4GBeRfKk8iSAN2BdWthU/yZvbiMY9AormgrT+IwpGnylIE6iPRGRpSNNID5hI
C5MBMFRGA4tyVMi6IDke/6W5CYRI/yoVHGRRViuVs4YxZ0JSFjeKMlee+HCmFibvVkngVm5llq9X
xx2K8v1ho7ZUNoeHkERey+If+PO1jpM+jTWgn7vmVBC/pGSVN/nLXHvRaS98TuXnE+7BDS2hekf6
YunKeMnTxy3El16AbvgVzJzchWX6v0NDlvJr/Ec5gTCyAMuATmBHrAhCsDnMg88zeGoX8bN04GcD
13aCL1ZQC4srBzgcpo5L8xx51Xx2oPazSvwDFm2EEpkeExbzDc6oNgHBqKGhxEuYNamF45CJgUFt
bY9Z2lmPk/LK3dPPjeysog7YNCnzvwPQ4g8iU67r345rKqdZrznbw1lDtVHh8ht6wl99sNQUhXCe
/V4U/VSdmaJD2KkfIbLJeCMKb0kYxkeChubelLxJ4syc2UKCuNeGJYOuml9Q+6sv8GlRvDB5138D
rpT0rzbKvj/IePVBrt5A5K5BHj8m0Xpw2EnjTiLfn6V42whVGnBuErFN1VeCyQR3Kc8AIaU7/20k
Xl8EJsgIP3HNjZrW+tl+7gbV3Z/uwDaA/fj5idD1t5FzMekbi00XapeLD9hv1V1YFARIjpaSGsqs
Niw6ip+7qJ6UcnoFU4WuhV448xLcMQh90/fT0jqK6vjE5nIIaigxDWvmxEWP+4jwVa0yEQ/teH8B
pqXbljN5V3pZX75qwJMJ42eu/HaxylVuEM4dc2xkLJbU+i2A+jRvh1QLMo5zCsyhQKW7gaeFYQpL
JoINfmxBdYB9xQR3/EgarWQYINLKW9luU78/DQS+33wpb3Wk1h8ytxmBfrxbilfxMYjGJxo5XcUu
1gfSt4K5CKRiiw3+eOAp8S2JJgersYMPBPT4dRyonBnhouQVIc/zkfALByN1YArxjaWb6L7xqdBb
45twqUcxtibLgdD/z1sfX151gMOVqGCsX+W2TAO7lsLHSF+dJW7BvdDlvB16Isg5RdokAOjbIY5U
QLpWMig1jmascrbUlf8ybbsiGK615HJWAiQzrtwcMyd0ZeK2ubFdGpmIFqDD2YyM7t2Pn1tREhC3
K2v53x1NAoqKdqc6V7dJMH3vogC1laVzX5Ftd9NZHi68ddXt1d9Ldag+2ZVGwQk6VNZ/0Zyech1y
mKkC5m7DNgC/mfwkWmvq++mQ0+ncyJNEIaP2HkbwG3enEbxBIxYARbrPpV/dcfl0aYGGpMgP8hK/
gIlqd1tdZOFihfO2Kx2TR5FQeEvaOlwg04PYFvb+nhImjz7xQi9dVl9WGU7GJHty3RHeV9kGOIYw
5zJRg0qXgtFa60WobCUF90uaYpFnazRAfZJ9bkgZBYFs+oTyMRvUuNJv7GiQoB6E6Hovpt4s725P
iZEXj2Pbqo7OdC9DJ8I4t1zrIhF6cYtsZci9Q2TUoPp9HA4hZiqAd9Ab3y/BlJfFMVH6mck0Bu6x
BPzpVM0U1TCHNQm2575l6wkY1qU5PqNiELYv74EVPQQgmCJYV3dtIvUNoHp/KfwGMe8C3PNnbnLE
qJTjEwivjxRYIgffoeATu94GhrtFe/B8rR4FzNF8zr9bfnYFRT2UahqFNy+lZPydbwoh4a7a2LYT
f4DgrlEpUabgT7dHjZs24XfPXB9wztCR8UCEWdNsDDu1s9tBzD5IWsdd5YK/YovRvtqRSPeQB0SL
Bq2iRDIa1p95K3gAG1vLJ1BGRjN3+kHwS2BE7zgs5NQx7wMQdnIUqNPuBa2APIJu9igquehwYEMW
QvoZnXjrbBeCSfd1SczftfcClkHOWfSLdYKVLbmybD9rWd+9kZGFqFjgb9jzWXos/PIvd+gl3Brw
8cjrrftHkb8nE6ZkEAvU3foXAo6YlCUPEYtOOjIzS+JUCnlxX6lPpQCLX6xF/7ffRzFqfJ6tAtzh
j+82wJ6Wg+kpp36rUcgHLmUtifMtqdkZMrRH1dSAgMZDUbAlsZO9EGzO3vuhx6ZGbVJFrM9VAWas
KqImFs+8pxhd/+cHjJ1yN8/fOAyfoJveE7mI2mC7CVumjhxZVTQzxLv0+/opEakMjojMkFCM5EjR
p5tc6GdmAsA515x/vOANoDa73MzIP7Dr9yPLrtRTPCa66Wby4LnRaM/gStvD65fKzY/x9o6miANH
BvgJrEWwTgKQsBLYSuMoK7q2rlPjOY42KE1x9gGOSCCLaiy4Ac4D2GK8HFc6tv+VN+v4F/skThLc
wIxDgFk3R2RXPwnxLUnOx1RjvFn/oWgs0A9BfhDXVo+FoEmHug0jFguG4HKnciGDvGFiowWQUDFy
Q7Xu8XvS6tgTmQv4g/v4EYBa0VrpDdYAxGCYF6aLEQEzCVkuQkzIqn6d/8fFct8dd71nDAvF5UOI
+DipR+RB5mXKCCrXyp40wL34T7zhT4BGuV0Ac+8Dqe5ih/tmKbDgRpNL/VN4kW8CFvo/uv/uBC5S
EgA2xUSUwv/j5KC58DBU6Oewoo7PYiBLsk0jVdevL25bQMykTJ+7dWQsgfinZ3NqF+GHIQztMlTT
9rQFfV+CJZfTBf1V9JIp7AeoW8MXbW8o6YX/1xSs6tnehTfyFM9DE9rob7PVSVjO9jZfpRY3CD9h
uhIDJ2imlb3bBqmGqUDe+p4wTK344mgXoS1MWPhL83/Q5iEJXGrJ2ZWSJS93rbSm6gv/9r6+WZLm
jGM5BObTPRh9P1coNuCz+fcC/6YVcFjPQfmfrSp2l58MIwD/saG1nRZj+fTF18IWs3Q+u5F9BHrv
gN1xfSxAf7P4t8XRSiX0RORAo7zVR6JnHvn+fFCGwA87aRvVlbwFIxy8FM8nU4TJbpBMLX74Jryk
A8PLgC0NxdUl+ZRBwjoVeokeXiVKg1sl1riVtQaSD/rVhyaK7zRYX78R46+pazDJxolkwidnl3W1
4VFytd+gYBHF3uZjzTfXB97HVy0Um4dm/GVW/Yqu3SpgIT54pV9JLHrNqxVTLdvf7oGRecZ/Wn0T
yjVKXunalYOxZPY294yKZgkilxtf9XGhiXmLq1mdiNvoA/hmdl2Wnz0iFlPBqkJhy2222SCJ1OHl
3WJ6grYtMvFvfmzOEXI2MOrp3klghKQUm/zNo76zSWMD45JI+hWmT7DvkqHKzmAfj9ErLLPS8Zah
jr4Y2bm7XhvnN7p9aQ12xQUWSoptwe7f5mgOZyF8oo7I2ui5ll7fX3esH9F7dVo1BRp3Cgh5la0G
iZeXh4jzC/ZSvj7pa8G5p9AB5CFJG22/X1zrrpD++za+/EgtzfT3LuutiBswid36vM8DsQ/3vpuT
48UCoSy/bqyUnO5qT9cjtKPGnE7Dn0yeJwFsZS6eLANPVVrvYPAc9QrLpvV6JZX0lc5qXZl4iBZW
m7Ehh5GjP/O1ET1eSEqUp3wqaVOIfy3HHobNxrua4uvJcz7hyCVJrptO2oCtDKzAt+RqsIFeC5O3
8yoNBEcVrtSvxDPWSxB45ZyhoBNFswVbK46WXF2lydktzIBTDcDPpnQxBQO1hR1q4Xay43M67Gyf
vgnsE9X5rdqGQJR8IXhD0RpMinHamIPl/OK2gOqe6B4pZEM2cD9mNIk+wlMtnjTcwY/WB9KZ6E+0
pPL2tddOm4kv2/CvZ+ZmjQOrxeL2nJEeSF98HcfnzFAPwnjNHKZ0O+peogtXpO2+QARYlrq7y0b6
qDn9+Q4vKRaXIZYv+AkNfCmgeBePRBwq8ubDQ2J+KTDA7kvevmyhg+GR6wONoadyqviqHe+y4nLE
KkiFZclOYvcyuIJrRShecgrXZfmAWTCieI5Iv0u2B0Oz4m9xwz5zfT9ccLN/4Jh9mHiv7h00W9q3
NWVFkj3NLRvrSOxcpxdxjPvQvEuNP8XCIutwhQMZuL5mF7rDcxaHNxmgShljSq8HlTgg5xyvy++1
IXLCKlk8FDsEnkrE0rATtoHMthm9dDsYrQcw9xTCuXpyNx3Co40UU/15tdtJaUz9rJmUOToB9D1L
6lk7Z+mJx19lOTPgCnLa6nR9jtU2ksMYRxL7WiYia4jUB6T1/Uhv1ZyL1iNcQhhdICSbA6AQz4Nj
h+IN64q6ct4CRqJtZGlevxUwf5jGoJ1USICJIVJ8PIEjqdyMhPkL8rafyGcAHCZpEQcrvB1XIV5S
hGI5C+jaqQB+3gnxZErqmowDQDiBJQ78c6MefjWL8xtBb6W9uHLWbKaIab2JhOQ8Rc6rmzbgZK5u
twWjkTOfCPu83Xyr2sInUPGsl1Ujql6HidizEFC+KxxjELNPqJ8i9X7XwWS0XZKOKqfZI1YHQy3W
1PqzD7gDe9vwqJIuy/z8z1tJ/vYR8QOQYfQNphR9go5t+vlA+HAzAihuUXVfz7YD3LAkMKVRpErW
Kk0LPM3qgDTNJhxuWNWAUfa7wJ/ut8maC2wcJy90vcIbwUWbneCD8ItCVMyewwbwGIE10ePKwotl
hAa1ZeQwwuHxADt6+1iY/D/EG7vRZsfl+dS5OH6/YTequIGkAhY1aqimTS5OeFHqZ1BFu2BqcHuP
+N5qNCIhMrcWE3sVBeQDyyQhjdxwsbgOkzgc3uj82hgh9ewG5fJcBnaUSTnmydBaACMvK6xAMdRC
m0/Bn4x1hWhG0zsb5txUXKoWU24+GP6kpMBUmZMLKPK5dMFfkRaXXK08wXcGDr7LkrhMThEC2/08
7ObGWfcDZcaLhLgFxVTp/RAQR3P3y/bXVHHnMXDiafD15byG3TQa8b+BAR5DWV5+pEPUBqvO3MAX
5HWeQdi/2Q0YvYdIflQBQ7xsMFcOxGRLWGkfLaipNETuK7vsEKcIWroVLfSde6OMsIkGahhH1heM
zRTtoHGxYp8P0y1DC9w7Uv10o7cjfrOpsMzbJWdemcKNauixjHz9Kx0LhfZB6jK93K/sEdY9g06b
zbgLO3Y4m/iYI2+7jyaha61ksbnkpro0Ah+VGp5K2DkUMTVIpd+HqaNXuAiWlVtsQV3HS9VUuV7e
Mtls8VFNWh8S0P+SFkwrtx1Hf3sGW8Nwb5rGoSfxpoFqo03zRqoTfTbtj4UgXgMcV/GwMOA+VKSw
GGVI7jEQX8b4ZP8mQcbHdrF/maAiMiRZxwtkBz+YPsX+FgEgI5dNShHUIgcs9Otb8rOjh/5fYE0b
b8gf6q5SxtqDNmb/yJsNgJvltNHFTSIkXcfBCyhmLHFcvfRkdejgFn+m88lKVmQdBszVitJeeHiM
Nu9/KweJoRbXt76Pfd5BYsz5yjuogJLoSpdI0+Dp5r7YJ+BqXfOyBcJTg8vOTcLa30+mDtL/AnNt
oh0C9Q27G7mCQdiJyDndipZcLhP5ISxyOKiMFnjUnTGjDXTdKXzmceQypdWATmaUuRq7MujboN2Z
c2kduQr6WwIEfOCdO6kqClWz8Yecg6yzbMOAf1SI4lSD8BMhzE/k+ASE6j2uxDPa9/Wy7n+rUekx
aWL8GjB3iU+Z6H8HPtI6oYupyt/nR6TU0lJwHx1YiKBtWY+BOqtPCDIwCXOSbtofBNmwcIIHzXGG
k+Eaw/Qdf+Y0Yrtc2de/cE/OdrA1YvlNhOnqyZ/7DdD2RFpnDxvDPkXOpffwRl9UaBsvCWlozJDq
SOfOkFun62iRs+dDifT88Fy+JI3rTS/iCL31BHVVONRjbIbnH/PEB022zdIAB/9o0lZsKh+8RINz
4yG27FeZbNnzg4XXt+depJqlpBHOT2QSzZUm8VTIQCohW5SpO0/jCe+e3/8MefJhFKUXSkef+C+E
FLtR1wp856hEjhSIt+ctYsCJw250+QeWUu7bjlo5BKqKWj0VpliaTtdPU65blGhK6LHok3RQOEZT
2D/aqx+xMd1elbRfIbra9ci+Wvr9p3ys711uFL5JpbGre1j24ehEaDehbVlxzT/kFZDE1jKeW2dU
x1bUKKXRbjgKB8C3Cy4dvwqrXFTeFfNNaH6eIZ2eBDYEykufrXHRrbZd+BBzAue3J6A2cnMdWJKL
+EezaOJ+IA8fVQsZt2oUMbNB3JPCKBna4RRSO+w1vaicIIbH3IjdVjqK93c5dWBKncnC6TOB82Xf
3XFrwLgcZSP8lFc5YjKIZ8nVMuQ9oVSe14j/BMArmQTZJMyUsMLSndGhBLP+ZBpHhUdRz/aD36jI
N782S4bYl5bq8A7tgleEPFR4dxHuSAQDJ94x4jH55ARIq67efQsJ29w+FZzf+mqjpuS0zJldKuoT
gdR84b+RM1dfr4hZ6KVwoTbMrRsAPMWPykjkpDwNyFe47RTvCNtGA+2cmiNuaOTo3ev4yE14Zw6w
+pKGX7QxEvM008qixDoEpB28avyJN0XGV68MCSZNatZh4t3tS3L1FRzaqlVk25UH478rH6jPjvnm
j2n02JOcff+qWAAe7GzsARunNv2In/YaldlVHIOylNAFZwhMCyKCTIxhrgvAbdTY6OAWbvJ4qMy9
YEEQI8Th7RSBKbg02EhZKQXIx/ENDpjx9yG8A7Rq+473zuAy9HBIbHBqeriAX1VVj3QNtNiOqw5n
erLH0QSDtmEcTW4o85YUI57ERblQFUh/JjLSRv3RLmcVDNFh4sb2bV1LG7ulHK6f5GQByB9W2Cm6
lVRg4UuT4CKukulpUwUd+HbaXYn0evcgcYXG+q1Q7lPZaaKBhOflfEqYytF2D5p2aJ7oOpI8iQBA
EVGqpR4Sv1NnmuHusinGiqVkx9SyFAHVgUOhSET73oIGI0LxDGABN2N45nj1/fMp7apA2sy/Pb+8
4h+rQRmEliURRSl5E1M+rjn9bstF40ULRkUuKHrNjVMowZFvuAs2mOVb/GRInF2tQ0aOvjMLlmiY
96tJY2NKGeHp1WXLw8Pzyhf4aJ3QPH4zl6rvut/CqE12+QntZveJzzrQf2xgP2R44AXPY/Ldzsqo
S3IkMIngkWBUvJ81mBpka2ZeoDzj2NOc+ikkvmRjJGIpyRb+h+nmzr3j3gkUgnHFk82wEyuSZRv9
ZHY6/GN2Lm4rri0nejIrP3XTbC3gD0DY7GIp64qLQJCAq9qaDPhtWx9C8+Qsv2a+zMcBEXeKbAzj
4117/I1ZnP+rIZiDFDzPa3ImRernK6MGhtcexBQTd0ftDrt9d2lG5jtlT2mo19PP6TV+xKGJ1NdD
m1SC+ajAqs4ab2h5KUhU3YXa82o6YhiwWtI/Ny0+kM0KOfAHyYAgcS/Z7p5KB9AYUcbE1wbzNm4r
LAS3xH8aMfrDNI1Li39ctjOS6Erhv6Paln/eI/pQyJXEtVEfNZRhHb54J6mtnJVbIV2ao1G/t9pe
35qIVHhbVBqVN4RY90vYUo1boVN3C5S2rsJNMA9n2w8CqN5hHxMEV2uKNU4G3B77LBoP0pvE8sq5
mk+RvvhryplbiLKzLMH3pfB7eE577IQGesLQtZBatUnp1h8n5YxkiwhjPs0UPu0nnET+NRY1dncw
3pyxOO3IrypVpAru5tEW0DHIDyf6N08xCdTsaG9nPpi0Lge6zqhKkSWxyMEs4PEAIWcUwPq3VSdu
QOuB4ZDcBtNfnh3cqbXXOeYNpbmxbH4xnUv5U5yIe8S+yNqMz87aaw+NVOKqxnOkSk4KBXS1kzJN
ORBvjO5FC/yer+2uBtSF5zCxDVWFqY58twpzyTK9zIzZ/tMBN3l0i8X0nqesrBeVy24amkmPKDw8
RBV3PNOqm5mloNr6Y5Cg101aQHivHcieDRcytz1YRkB4vu2C0Kf1xDpOTyxHAv3YjnB0a2gYr0FD
4nxZet/HsTMzCWAlti5aykbvqsmLhQ2aCMQQUOL9PI3ms6Bx9MospMgXU007XqvZjotqbmcpwjcT
CeEtA/CmvOV7IEOEwCLNkHnixuE4Mjqkmjrp13F8kH13B1AMtrpHRXTGIpaRplw7JToL1KaYUpmF
MHCOTkg1R+1E9I6nU0pO8tFUiOSAi2uqazWbHjTiT1+uTaeQxIbOsO1NIWM9dhwiaaKYT8rAr9tV
J6RAoX8YFcQQYWSKsdofbzWQ5qI7pUoD0g3LXDvJwtaGALPMTfS9tTDJ2xNSO+FIV+OkV+fjYF7t
+ktf252I0MWmIzglN1gs5Oqbu3ZWOQjIbd/McA3/voVB3AjD8jrTtmueXbWEItR026OxYFTziL3l
NK4nOWKEbo1b2abJl69vfQ5u8I3JvG2itC5ch/qZDFtPGogZrw/5QUXTuUMCqO3g8SeXJvpz3HHC
oZUgQnRjrQuQAl9xU4oidZB1B5gTk0G4FeOw1ze6fn/vTlmo8sPkxlgrOkYsFXeUpTkEURoOzImf
kThL8aXeFeL3dYDlSEsu3lR0rGRuZ2swL26aAu0pYbVrxjGuksYqnuuL2rq/0baV3oCmC8zFv7GL
FwdGLLrnvc1PQdsiWexim9pueGh+egOyaiGAvpgL8k6QAvwQHVYXo3V8b0rOSk5UBcLO91qXjtr7
zPI0/02+h5Ap5Kh4SKHchP9DgPnJJymUk2KFD1A2Hs39HW1zH+mASPoC/pqtY1BN3hnYAFGUo38o
fr6CcfvsEaDelr+VDO1Y+rhFtRS96BVZJf+b8qK8s6VnRfUUjrsLm6AgCuAoIRFcJR3AURJD7j4J
Ci85IuZZ0YUYhlgQsI3yEm5GwbrmssvEwFiLMSAaCiNsUsw1I7zvUaWZ6uxfrmqOZ8SSlK1D1YAX
oV9+W6phAbGaNzgud4hJBTT499WwE/N5u2Gflx6jlD3+KlTkLv1w+FlI622bBRiTSW5FNUkTNc6c
Tt2cvJd8UgP6CTPNui8iW9mMqJi+lACqTcsDd1Z1k33mh6LKWly9NKlPTKYjPZ1i7WAkGvlBRkBX
4gfqHRl9PM8gJ4z7TPZnLqB9xP3D27IXfn+b445wMkGtFLLFBp6UgTheVuJdeNk5i4V7yckvXUpi
ESrAupUlfTvPdsQKYs+qbie6aYSouv7EC0N3IHr0vM96NPp1wJ5/tzsg4peoy5zDBfkoiKv+jB0c
zO+yrNC/WEFRvk+e26EWnE0hUO5sbgmOhvQgIR14ONA9AofpqnT5xTPz9ZTSS7IQmQ4DWSmVnwR5
487t3oaJOB2UOXXUrN8nLQ/U8jjX/UO/zXk2kg1oUIY1aO47Kfz3/l9u9Jcifo19jFMC5f9QfJTg
E7E5R3iyQ8MEhbh1/1WRS34ED9BovVQnc8II3wEg+l8zW1nRylj2AQbhVmJ1UXZXAyjXO8+AxYh0
jvrKN3uSKF69a6mbkQOdlSiBdahi+fgUrFwdh+DCYxjNCQbB9OqH1PXu4g3yuaa+eRQtSp4Oj/f2
Ann8VLVo8XHq7ZKJEsBbFpz69XXhSQ8RR4d8GcTmpfnTfybxHrx78XlE/gFW5DnUOBfTV84z19WU
4FiDSR2Gt72EV4B27xKjtkym/mMpHb5J5h5v7Fn5a+WB4UV3bgi+ZqIsuYeUtpD88GhUsWR9zjCc
HMO4Vp9mrBWHsMNETv14s6lmwGaKSrgSO9kWfwM+FXKN6N+gdqmIXDEhQR20siWpr/0Ap1+0QXGc
NfB5UFYNtNMWb49CZJu2WHpDzCzZ5/gbWEhWvska0rtU6Unf7Wn0hwfiHWwPv0ZrF+z0UJGMqwvo
Bivfk2XpTr5DQ2LSzND05oQ/cdKaCGpHWthvup3JvmqntdolHZKdASCGSsBBEpv0fp7GCqeqY0GU
PkQS1QWX937emhGTzzd03ypKL3HAyoDLD0o5wT8EFAEWcc1WCdHJd/9E930Nz6RDTV1aLrEHgURV
unuHeaLX/rdHRW7yp2r8sH98eFMMe4WGEbanAfUOvFDDgZjwsKFCpSbhe2GFal9M1rt8yta7/bTg
V3xpaRZVKeK1iGyqxz4xvpabkYuirEd6tu4Zobg4G97nyG6bJCMkWWnckMSqWTG+hqSd6dOwhji6
gWbT9Sy+IwhdyU/Ocd0pH+2OZeMEW+IUBk4MsemWDhzxeY15Hsq9Db49k1OOFcYAPOFCg2auTP9p
FKtunyvoaQiiyySuRe0OMyZooc46Ds45VqQFqClZ+QbhvYRoiW27hzcCfjMb8T9Ke0I0VBzUilim
t5wc0QriMd6SspKtx8l0WTdX3yHMVgpqoIgPMWcvvhVS4jKSgePuke/gEvYzt1HU2xH6M+h/dPO5
kzi5XEXk3l/xayrzZyiLcCMk+hGWGBl8o0FHhks01yrGFZ3Ojchl4GMti8TT9KBUZVvLz3BpiyTP
E4W2wpeCPsGKX9UGInf9w3eFCdAUxFhu78n7Y6QOVudfamdIDdDxt6zvsaIBZRS+0OiNJIgQ8Skf
MPLkvZqcZpqIdBWpTboc5twxgvmHAn0BbobkbdAn3QVgJZq2s00kSkqaoqlgSKm5WBB+TuY1r3z6
M8QMkdoiEFnEOCr1HyJVuC49VVbTUatesAEu7r0GbrbC3eLzj9Y1+liWkGxLVcYiLbDWnDupneci
MGWNW6pk5Dxbm1yjCEj01FknFniZtVAYvVhZR00X4fbrOEdUQpScxkJlh4aHJwE9Tc6dHb01/oxQ
ug9OtGnUyt5vnrkNbxHmxDKTs1Zo6bQXCNt+8oxpO0yv85zz9lKfb2TaFpHzpvRk2MW376D5eR5l
H6RCqCyWgyjGThi1I5sxU+/yCidn2nkczMG3B2L3VgqstD/5r04W+IxZae0srPi1jtksKduOsEAW
EfD9DbVPL4sY342TdKGft7FpGhOuX3h3Z0QBz20GdsaZMjZu2lBaA/Hm/ZWjtUeHwk3q5AAqzo4u
hoim3JFL13wuPUJkK7lQLX9XTkDh+c5PvsVpj7yNOaZhkcn9bjvgbUkSQYcgT+tXFvpHSjudx4u+
v5D0fM8asl/HzsiUk1PmLHUpgEoskzwXxvSrQalQ7GC5Ii6cl+jfbJTeXtfjwGfeBZA9YPyK1XoD
3fbS0HOiMJUkifMprlH4elWJNa1GI170dTM1WfMcA+mquclxtnjoTseA5ye4O4kjHNxZJkPTmBpJ
j5bnZOHbcF7LYCzfCTyhwPHkZdU6OTIFz+/S+1X1iGompqpJ0LepwnEmTfoSZ+NsSYXM5fhiSPcK
LAWnpwNgRWQRgguy92EMdQuebItv9PzRf+TGll0m4vwjNKoJCQeRvxxTQkNVgqJDCHolXxdERHgO
Npjs8WysSCQCMpcHO3sIj3SNSZeJFZJTqycuyHzErDsiLylMY7wXhgkAydGPuI/G3QT0BWAElx4O
nT6mVcY6jVizqwQ98TNGDXJyfKppOBrTlCtZ90VX0Wo19NVn1kM7PDBKA2I+VX/3///RTOYG9qGZ
ijt9UTlm/70K+DLntu5HC2nnQzH0DC+iBBGcMhYVK6lhkP6mFuVwosxOeozS7t8aqjUy53KEiNn/
0e9Bd2OgiPTcsFupCsv9DBLKeGzf/beOPNd/jk3E0sKGqGTUl8HjIoPw9DL32hm4PDGN7plFOXv8
ZtC3zic4eEBbRjxWbJFRiY+14fru3pYWutV3zBoMyfnmtqBGMiFXq/qNKjCXvbkoFr9gvdZNCB4m
kY7Tf4Nq9QMl1JRvWRFlgWUjKnh8AwAeiGLnFRdWs4g9a3WKJWOdQuyZRrRlDImqqYaKehuvsnEA
G7gsymY2tsrdvd/4yuvMiQNR9U18c2JQXi+ynVEw5jDd/33XLe9hdfNwVkNZaRZo+3gnScaLcXPq
MKHILmFhMmIwVQT2CtbqoWeY4ceYxuYA6CviXIzIwhJpoFmcteGECCAOP/zzCKIBWtT6qCPOmqWw
MqJt3vG9ZBYx3FmJ1EBzwYl8muOkQqcnxh/uMWUhMCy3y/2l7phxW4u6MreoWGpHpBpWDDJzFGKZ
88Fcmfejz3U+jFXkmeGusih3JWWCEb+A018pOGgJ/lUmsbKpkbNz3cRP4Xeot5HPRW1oHNxhjHvG
oYuGqz07/6kg9tRdimhLoegoMZaVmnYj24hwbhrf+deS8gNMRJrt1+c728p3bbYXl/AFzY+qLowF
6Q5lgJukAZM6144v5uIdsqWzt+Ih6xqlkIOm45X7OwBBM41Ma4VOt2FstYWpInBxaewjfkqqu1Y9
fUjvefk0yto7ptOylc79HwfLL6xAVzR+Pu1rE9NugErW7Dxm8NPK2CRpUrsUzPnSDPy44xK4rSvp
qq02AvkuCwNIDhAbdL7EdS2LsuhVaEoYWJhkNwcAWLExQZ9B+JhPr2SSZhYZhJaKKNOd5jcRjsP1
ye/FJmCpGm/LrZuNgcv9AhjL98ADIx5b+gZKNCheZ9vKO1Qxfg1b77ggyT1/FxCdM3z8O/jQoLDL
ogneQdZy/Nlye2t/j34Qt0slIYxidXzUnZbZ/zJEF5zRUXvB8fExfOA05OxikPe6fjWP1/yvKuYe
quidvBQD1VZ+y+mPkOWjgc399mvhJh7FooKIk4SFW3YoXOXKqk/vTniPOBrWU4srb1lOZTcj9VG7
HlR/osxY2Hn7QL/0UhY3gNQB5Ooa/gxoqg9DIwzuHLSE23oFoh4liJKULwnc4XgAE5IHzkV2UU4c
1v49ikJvUfDnBld7ZCe1EyEmSie6YM2SIdnrlRKQW8lCl12OddQDZLcpBq7gzxDInrBBg2NyhO8F
eJmZwtXryIIULB7hBSA3wD5rd8BykdA1ZzmI4N0l6TFglLjVULc+g93QWCwVfuGkLBg2zkQFJBol
PWvp/teycmCaST74PUNJqmBVcTAYc2nNEjNqenpCdJJPuF/kSPEG9yHmoh/w2aPO8qIzpR8TEyhz
aSs9ZKtFyWyHcpTQyjoGXBO+b9WBFJQLCfWIW6UOLEwSjyro036bdmwHyGEgVjeCW76GD8GItF30
N53SDtAYWFZXe9FIEpVU6GkC1ks2uxnONGqK5rRsmISs4n+H8wRdtv2aCo43jt9TIt+AODadF7ji
GGAy1vOJfaLVfAAxURzGQuuUeHMMV+XTFmcUWQchP4PbR9kD4qHKe7c7brSOd8FuYp1ULgYGPFy+
+gLhDmbq8h8dEkJwdTHQeSW637Ve/M9fY3AX7fNjb39L+BN8/337kK9BBOkCDrofjYQkH8aemqP8
mNwGy+A588qnP7gjEA6w2Tc1UeTQ74FA2Ijd+rbGIh0ZXd4FYddmpyevoD/DN49w0Pox3nWQUCed
wobKosmsKNBGEJmgkjoH3woi+o/k1H+a7iWXs/kBu6M5WDFGw8yLDQo4Yjd+MLEjwcSamwgRvUMm
y2kJEUKLbrwZ/Z5pHqU3RfsLMEM7r4eTKi2XQDiC1KGRkMcn//ha4h7lhs3uaWSfQTZlYdOpTnmn
Ppuz3yL/tVdhzpwu8pLtjfiQuD3FxGRljLGnh7pbHZ0Vk9ATAM64ZWIdAf2mEAABCp9RtrcYmEk/
eN2wUaS0mmQEob1gGpvL8RBSe8LlzB6ll4DParMIhhwPTkojP7uRK1YbbP2XZjJBvkNyWN2DkibE
yrQpcqVNW2m2ddc4dcarGmBNo6RTmETLwexXTZ/4FgJw9afqi5459Joh7O6ZBUmDWufCbecK1ETW
jlYgQrON7fWWU50sAgVNQ4NDW83ixwlJctZKgapBye8DLPhSWCR6BmIRaTSYze4lHdso5ySJ0ved
Lk+VGiA2PKX2dIKsmndWygfnK492zBPyyo0egZrnPtKWBzHc9oHxx+adSaaqjSm7ojSPOCCYZlX7
/cLn9kmeO4HEkGZXdbg0wGNCMhQnE5uixliIXjqHWumSAClRZZe2+hb35h2Tp4AcO8cI6Av+7VxI
OVAqrJpmuTyZW2r8AU3rDZmntgH443xWJAQvLMO9FYzYKrU9U2cKlmehn7xI0Q7Hf8fKIi+1436j
vN3tVlSKIeEd2FdmBXPpHNNwAQhAntNor2XDYG+CkMhljhjImJpK9PKpKyyhNAuWv1nFyWv6cKUV
Gla6GKAaBoUS+n8xVxjy6l6NbUI6zG0hpOvE37sanYVDY7DgNTZtsFQtQr6hEYm7noYHm5QBltnd
TicwEOyxSXvm++DZ9svsSxOgNE9SB9p0stdxcY+wjJk6BtWMxokH5ZkGPClx2kc99vNpl5SpSat+
0C1IIeosfE2U9oViwa+Hcgduk7ZN5HUL+d0fEev8CeZGUcSrnb/+PR5JDKrBNPywLOTQwTmRpXaR
k0dP/50Q3MjaCtLUgHW9IyEg1XJXZQf57VuR681Pm9aemHRRTUsdBddBx8NHXnIAmSib6TyYE9/v
Wzu1i7tCr7PT7q5XvSKVfHBZ2vAzZBNtriqLY0yHQXmYV5cNjaXBRcMoZcs/zqIhwoJFZVbOgQ//
HXY/EuqEBbXIhwhE/pGakREgTANzk8yHTXxX3/Hf4Pk3OvLnxM/h08w0pif17zUS7IXv0rX5R8nl
pMIEvrDR7anDo0weJhNkNeXNGyKXVdjtQALscAAPmA32ez443nETrLpsZ+MCEta0Aj5k0W2fCXYP
jNkxj6lQGKiP6wJh+wSoYoGpSZsqldoVeJ7gd6bs0cRkSN4pi0u5CX/9ZvKnpUDp23gv1dTnGsTH
53OUNC6of22aCorHpsQp3UnhNbczJisft3oCtWgYAUr3NH7J7NZcvV1X2MYTmigj/07EPNgzOKL5
yQt4+0RDp1gX1yOGMnHblhYWguQVnoN3Z1yP+UQuF5jLqfLxekoG4lGa+bb3r8FUJwwWHMLGX4yt
/YRjCLxVaq48cPD3XCR5ZPiWSVRI9V/yqRWYiXa88hPZ9MiHvXLH/4+RK0j3F7isqFmSiMZdB7jO
hCP1f8a0OJmfD+/p7jHG70NDtZNwa0Y2UG//ykTVCm+fJekMmtexiUC8jrWnQrcrmlv43LhBrxgh
aAsrAkyoeN+q6PBgHCKU0u7gdvub6VHpjMvhO5Y0Xt/gE1DIlzBvkKq2/VVB0RFO2gtLsay7PjRK
W+9BoxPUI1GoscBlMd83LTV9UAxCzP0PHhx9rawJt926+gJ0kvnWa85Gbq0h47HnNXfUzJmdSx+w
DQt6pkRIULqQw99bD4GyiV2R7U+3QVgXyo3kxEXd9VW4CceRxhn7jKfEnisXk5qxlqC90Jts/DQ/
KezwE8qy3K2oeDx/bnXYtaK/ujWWOLPnQdKHf3V/TDb4FO1QW3yzqQUZfkpKAnITc+z3JcRltVX8
WBKLBZDBu/p6/uax+dJdeeEloj/kWYMUU0YRhHd8Lkxw0I3YDGT3BKCD1Pmn2i0OhEaxINc5lLOW
kVfK5ClqPuOr3TEsZYgu/fUla0dqA18P6N+OkFPJxGFhrkMMrasaCKF0k9diKuIaldZwNqOYkifn
7pWf1sNpl9/tP2eYIWz+IXctLmeIZeN/joAfivilV1j4oJVkTgjrH9LdSYfIZR0NZNchg+dy8yEi
pGrAEeZ9CAGZyMRgag4NpHJ4F+qPutM3ME4QsP2vMX0t7clx5RnBx/4M/aUVxe4K9QszMh1a1SnX
jEiF24hap6GoI8p9U3dz6hvBZrqgTnOVURTbNQiIjzYYjOc7SRw6+kV6nu3iN8b+c0CJ1EnpKOEG
IAe0uaqT1E3KJx2B5VZAMmMFeg+s1PjVNpcUMbew97h+tnFnhh6KgCrJSo5eRQUPmv1J/WgQERUv
/yqAEwJphT7gcDF4vUGavljbKnU7QLLzrVDHX2ZRelFwYxlfaxWGWUYfW5XsvCCB6iGYu2AHV7FG
4TrsDspsmD2/y2FfQ+oLrs2O/+gPkeEA/8nPhXywvlHoLnVPC0ZcmlXm9973nrUVkkBnonTG4TtZ
K1iz1PiH/oe6krPOacR2nAlNrxyBKBT20NCBIPU5WBPl5hCYcySok21S4zYeeLD5HvhjjuwvQTK3
ouhLVC7pttNx3sf5LcPAoj9ahHKfE2ZLw/EJFfrtYbMbhoO0rwwxC0O1EaiBSRJVcoMRG1JGmjyP
+rHV9qkZCTVWjHVylBevt28rWbvLU8sWZ18W83Z34VaznXiFxEcQLeJOt3y49Jj3xdTuhTIm5M0g
jL20lXL/Qk31WEMzqLIuY9UpfpKwsZR1jnzWA4S35MNZVc7ZNxK16vNkQ4PDkuD/ohxeijO6/c9V
qSWDOZ9Rf4T0lA4PGG2+vkjE0zXWreadhuQpYstnMfZ7K/JxWHlsmXEqmIP47WY/w4C7GhBCjko6
W5hGeJmXXGqbJdyCxG5YIw3neEDPcFxpyPqOetDkWAx54dmgZMHgE6bUDBYnlyl15kQaqZBWZ6nH
xgFpjfXfSPbnRdrX7LNodjaavr7dQiryrzIJJU5UsfRKwYDXFQOsqG5Ci987Zza4G+uJJbjp6TqM
IV5GDCPaMua5PZ24YP3AdIpcKiRB+DYgOS4ObWYr5ECsX+Ay/cauKq2FT4JOH3jJsr9YqXzK7v7a
/J1c+8PtY4aOE8VV+uauPO3sGASuDYtJ53T9Z4aKKUGfGITVf1eGHtsZj4tYox2q0mJTRoVv2kQZ
SdE05Agrr1qes9vvYw9rWABy1vE7rpaGIZhfqRR/+9Ekr75pUDtK8R+8S1r1wTv/Y+X6fUpcnmke
lpOhKJrgYzvpCNuVS00S4f1b4hd4D4vwi+hijnXaRmJEkuPysa4QEOyCBF0Xs6ps5LjJK0Y2JnhC
6miNwjOxTtHx99qBosEnnLF4agsgHDstMcmPkE3BAhI9ZXUlB7IZ2D/5GzTFsLmZglYaXBaquURw
G2Im0bs91FNpRnIHHYg47NAnKOxbHryFhQV+IkTSXfKsJpKaJ/u2rDhTH0wxIXjfEMB2nZLjNAfj
t+EvFKaNIo7yk+TDeHajJZ55CnB2kQRTvr/Qopih53z4yzRkIJSJF8DRgbNEPbQuGgCNvM/nISk9
u56tj7VJmsvYPeqGvt+WWJTnZ7MWM9ZsPhkNOBfSNNeRZ0TyODOJJvvtxkLgTxta6eutTyBeJ4MA
1qB+3zL+mYfVWT7xuDovv+YFWREvlb/rfK1vyfu5ZnhpvXcfFxW95y9y4RlK4kDK4OFErmtFhZ/m
DkI/ghMQwTi32/1YlrsR67xySQmrq3TkDfVHOJG+4AV/1g6br8QMO/2UMB4kO6p1yM5Nc+NYSSMN
543hMeq60WfSZzX7yzJpnxUzwm/mYM+gCqgKrlh98BRGNIw5HyGN6HGNQ7v4Zo1yyXKIjJwnSxLr
B4BAre9wDOfgVV2P6jfyatVm6CJA2T27u3bo6Cucj0E1tLEv7cd+0wnDlug2dXiEZIe2kyyWIJHQ
PuofNv179ykxs73P9dqPPoQJ0KvPx/A3f7u8jqGw+LaPCNrz22qWQOUJhwE9yO/mkFEfYCu4aW7P
AmCKwVS7ZcUNpeB9EV5Exx/h3jnq/vFojKnHKwCT9HDDdVFq3LXBL/ME8QSJkbpGzQlCer0LDboi
HLieKPynVSI7QwvJyI63yI4qFx4KXvMNmZv6RuiloPNBDiVpxkH6VvbTotGvVNF5add/t9jtvYrA
dGlrjhku1LwNT6cy+hhCnNkxWu8H1SrBVymBbKtmwApCYWXvDD4mVYXRr4WE0d6vi7z6lEZGMSmv
zCZCrVKnpTEll9qiaPmNETLRKq5hZgnH04zfDKVI2Ozp+kOyT+obTq3aJzNNWU5NewlyFrO6qSjv
NIZWZmEDl2GgOhovhFQWE8h7d4rRtaTGOhunv/9h+5nxRmI6r2xKlxemTQPffUGo9qMceSH3iVqv
mW0m8BpGafZoAUzZ7nsTKue6tU93Vmj7j+lyoWlqAr6bUY+REpuj1F7f2Gv1rfyoiM/+/iVP58cj
xESv/DguZ9H9oAJFD8WeKpOcecggA9g5WSDgL3QYC6nUJXn7aU9QExAQtgunrb0wGRSxCsBUs6hO
zKUqoXm2cHijz6A5dWBD+yjjE3h/w9eM/BavCocDd9YzrMsM6/UHX0b0D31vko99FahvegbFyHFj
WUuEJBlS9gTxGH77YuhyNtwV0Z4FbATnElYDZ+sJuFBKExBtyjVrEXdPYSoa9nyXi4/ex8vBDtOU
jsupyKYlDBFxtr5TyyL0/K/M20AZODS4hMCEOINkwJ6dAp3sLbQ9undRduNUxEvGZ3I2WggxY6Qb
iIOhrSRfOpgy3sOOVGQJ02yzwnBlAH06NXjNA2IjT5fSePeipnX+53RNqxgsHvI6gdPGFqfGSLZA
eYu4/eyIo6JEkvFN4h+MGW9glzbqdLrx23B7lqSiV+RZWii79biSRvyyzt+QdbJtldGkAx3g/JCQ
CVNCnZvyXSLL/6t840DscCQpRSqgf83cnIZGROYnxbnLyiJY7UHOgjnyyGHNuew2nbJ97uP0d+R5
DZ80iX3xZjSPEnmTCCE+7yZuA/xKgdRkhX2ZId800m5I7iIC8st/63GkmUfI2703hzn3YsDpQbdu
x5RguIR6Vfr+MN12e0qIOhoyLTPyS1xDhewrBMGjuJDEnlnN+wQ368rbRfr+oT2XjWygd/T2IT/w
CB5IrkaBEi9CFHgRK9p0dgLOHQWRdJZw/20ykMlk1AQAtw7BpqeJzaltnAHiLbtWZPj4LqyzzzMm
/k6z1FOy2Zym8sS9wpj7e+0ixz3IGWX7VoZW2gV0Es3STLapXzDKl/awMFSq0kqPJ4JGFHxtlZrS
5NWwvCLqdOu2z4M30jZBkrKODvlv+Ji//+ontyEe+xhyALEhiM4ag7tVEDq1AlMr9jhoEVq42ax2
bRsb2XmK1ieMLJhYpNLF6fB4vVJT2f8LVsNGkJ0gdEpTMcY7kSXRcXJkWy0gjXzrsNB6VLp2n3S7
/0rj9/HYsfOUV9BpfNqgplz3kiXhbMVUrHu+f3F4EyQGyy5paVtwpWBrwFGkGJAkfHYP33LsVPU0
QndmoIic0AmUBNAr3napJ2Ad2jBUWN/KjtIIydD4TgSMXECmW2A5HcF/CnUwEGiX9jd+rlf3ytRw
CzRfZ9MHIDyqmeINFzDqKyFXhG6LWDEbTLFxjXXFh3Y/OMqgwCQX4PI1t1hWEXJQwJU4h8dDzv0A
mWJslReRHqNKQL3V+aYQ4TdqNZaVbCLZPf/HYsSlDmwopP/k4W8zgby75dWUODp+3aB2tF/KhouJ
nfCbF9UA2e5izlnwVOwwzsvzgYFAJu3bhJqQF2BuCHy19lzzpBzJby1asUoO7ChZ6VCbmwD41cbD
QZeT5caxjM7x3Tbs9WKLFuqoZF2jt8a2v3M8ZtUtvsZKmZzXm2VFdXSoX+kqqkdBmxBCjTO2tqFQ
pYJjb2xSznTOW+2fOEPGaSIjfJ8kKVW0rtxPmC2tdv/w97b4BP2rNyUCreQJBS8jytUatVTnWkmO
g+J104Kxevu1F/a7KTIf3S8u+uZdansldAkbitdIvr3wgC8W9UZf1QgA0elQ73gf0mPVwbknSLkY
lGh0lfPOtj0zpKLm4QrCMmWh35bV5T1hoN31v3kPyr8ZOFehPoEgC6/DGqf5ylNGakILovEWAbjG
QfSQtbVnlUaoUkbwlk46a00H5IbRTKlcnnZD2D4LAM8Zrp91EVC3tfoqpVIfKQkwrQ5jNq3nNqVU
petZCvgb1dlllvNxMhNTeqw8fJvh1HwiQafPooxb+4RC5vRZRfQWeEQSc/sKPybM2Xw7Cw/vRiuG
xdKEEzw28Hler0eAccjH6Hssj3qTDvXIDQyuLyVK53PZX1ait1ayu0Wp+HQvFjVi/LSQ4GqgIb7d
S24v/S83f7fN4vd7F3CStwKvY03EbwJhENQf2Gs5w8JCz3VV5aC4B+vfBE1YrQlCkXlgSTfHN4OH
/1SnSfJfIqAFjtcfb5wdg5nPkqjtodmeE1kMgboJB01Fj8wjc54vZuk7tFTUUjbaO6haI3XEB6vW
RZfjGP1SpxjlPO/TKHZ5sR9O6HJFVIu3Ic7myOhhrMnjF3S0WJuS5NbefPGf+aMVbS2/qYfBRlDm
6zyIIirTVJWPgGL7cakGxQ2oiMwhGjH3im577fTb02FGZ/EtH12o3FczJ23HEkZgLSI47ij45I/0
DmY/2HEEPq5lcDqfpjlWKmyA+wMwa8Adr/pqx1FyGJLY0A0fBzF3okmYTEOm+2aoqhIC9/oAmtsF
V1+ceOusOc8m8sUlRybv6JB/Ss2rIcJlYjBSwbtXuObg2yeN3Go9pjo+siR2sf+uHDCD7NtLHY8F
4hWob4JNEobaniUhdMklbmJt02XHQjxy/NiKxYJS3DIxBzuo7PV92hKnpNeCXBxcx9Rdbpqc94O0
RSHf5ySW/NC/eVV1OTm9Tc8aumZVi+JXOFicHKFW6beDMBHUrX0gDwKMtPivE+snC8PUFTir5hQF
Wm66ltcQkei/n78BYI/gwBfFz8AOUHv+fVq7cvu5gCDJwvjQ5Q5miFTG/v3bCL+5hka6UcKRozb+
6BiUsBedZ2q73ojLDgNL3M6ccGp/dsA0lwcxc15BV0XMRswu0vWTySAV0dSgDekckq84ekHLbDZ+
cVocey++LvyuzfUCsnB4SvhdXi+IC5sghP6Ig0o+MJOJmRhtV1hG2+KHYWx77gyM7IDQzHU/qa/I
CzxFp9gUszQxYbXrT3bqQHQeW6TP3+184pyvID87NSQ8W6EPNRBWDYK+uOtcosSvw/+8Hjg8CtPJ
VO6n+ufwJwxtAxhzp5Cvfvx0g1nxtiWy7DKTHHsYeb8LIhJ78hCjbLMSTia4YtkVzphFGpDzsdR2
SbdvbUtBH7LUc0fkLvfIju4WCU2xBJdaLQkIJhf/V01GRxj/qQcAhkB+lBHBgUvpWWQrSa+T2jqu
EoAwcnf10DEAGesOatcgMQLMAv8fmt5p52o0yKD2KhcVIL4zzqNKqPkE7wi0Y89Y/CqPiVcyUnVY
OTgWqgwelUWw9YBGDngUQW92LELje/BLHv/f7JNrKMr9LN+OJbS4hN40ZqrqIykKclgNMnovwNFh
NJHB6VrsLfluoRaMyTQgl2O1QoF9yz0rMwO1BLRJMZjeAYsSEiQt7MB6DmAYaIUCS91oIW7COmZn
2vixGVwj76LY6RT3Lc4hyjQYlQkoraD5GB46koY2f4IZmrxWhY4CGfU4JsgE/1wdoXA9q3RpaBPJ
Qj8Ae5hwHtMynqUlTR96flIkMnNzovn9mTCp5x3NgPSA2XPHZOCwMR2Z618pN8yFmTc1tww7GlVS
UaSpv7XC/hKVrjqfvQqMRCj9xszAwnvmuduH2oKXSgKf76Z2/+kE2mUKc2GROfB1ALsbdM41b8bi
TJCO3mHpUSYBMdTDnamZikhhp6kieCIXWSKOPYt+gjcBAd5KqErZY4VUC6nJrikc2NfN5YqvccAN
ukXGTR6eab9E47F06UB3z99gXE6JOKphBHv2ov7d+V0HBeEvpRWS6C/qzh2ntd7yQ/qxBCbLClFk
0HB6ZC1rZEbNyDIzNO/2kjTpuS2LZgbFQvVN7UeImZCsv1e+7BpvP2N0sPuIpbSS89giNCc/HyLP
VPNi4CrY/wKIu7Fuvr9nrxZcwKoiRxcb8XdKrPZ5Kb3+xb/7dLW4cjzOU4gxaOxTpe03jD9aXWn5
dB41CVgf7FHSG2go2IL9XFh7M3JUei6+yzYXxWWryf11TipXsb4Bh2XORe88lz+mVwf19KT3KIMm
yEGNXBpeAUuBCAJ8jXfDhhf3T/oehwnORU12H5gDGJAWzOrwxGwqZ5x3KLqhl5pdc6lzhfK/87TN
Of3Q1CBr7fVheL5LV8OdqBgk0USyL2psvkWRude4WBJIWI2uBF88DajxxJgZK6OccrFZs6mdMZ4r
1KVCcq7DYHpWx8AfSQxxjCwAdwuhJ+9jFaljfsVlwHeEn/+0+CTQA5omtScKWzf2Emb5NrGeKOA8
ZFed0v6YVJafBvAqYpa3YEJ+hhkpG0+aQHXsKZuEi9gGg5p2wOZeueofr/6AhNc8UIRmZXKyfhn4
yr90P0vd7w2loZOTreSdhrowbcyqWGnkHfRArPX1tzdHKPlS+KZ+6RESPv+4aZsrtb0cANow5vXJ
zFPbTR/nxE0/uz9aT1tYtxpE+J1i9FC4eNHNp98N5I0XYVLZVhrYBwGpbbJaMx0nul8pNQ7A0IO9
HKjPEr235SfbSbckZ8Q1KN5EaXkCrLrlTjlKMswwGgw8xtxb4wQST4/Hq/exLsXeDCTYr5WqlpUB
jKYx4zx7qdzgjM65+RzaQ6JMS/+7YUA3huq952ozT4mMpccZJMnf+ED59aGOTCNeshfCAGNMtErk
RF+XPS0sc0AQKPjPLuDSgePQvASVOis4e1nHKvsfofG8RxgBkO3WjOnKlzLe50ul/Zal/pqaLY7w
DdkRItVXkXQpuoN429uVk4MbWCeJ6/VQXrg1Zrhro+yt/+AqGdn39slEaNN3u1IOzHnM9ZP/DXiq
Kp4Vjq2BF07QIsc9hVMQ1MY6eHGbJSP8fYPAv9q95DiTk8J/M6uFekAAUXOXDLmaq1Zr0wUFU5RB
pHEA6Zv6VhK/o//cHBSBjyPvtNAnwhcH87dRi4TBo+whkEZTRd1ZypS5oS6y4y2jVZrLmc242Fi1
SV7LUs57ZkN2AqZxwI9YO4hz00h9/R6krl4/VFpXtMAKyxtIyHGYBpAqFTeDfAdVxHRrmFa5dila
qtL2b60qZW0m4q4IsfHBz6h7h7olWC1Oyn8/OuT3yBIsGrGAMhbH7rmDxhrzrLS3gdhk2oYin3Ih
FDaR7B+uSP/991ECnz7NAWfg0fSxYSQi0WF50Kx4sRHFctdu3kLN01zt9mtDWuKKCFcvEmV/iKT5
w/BcbINfOQWf0wG6EayaC44nAf6U46zmGzuok8Jur7lQmwl/gxn8bns1R1pniaTQxmm7pOdI8cO7
9qVV/Brfb6V366bJWg/+80oXyX3MzM7rI6Cxv9OvKeR9kBotX/HGiYwW+e8VPlmfV9Vbt3FgyZR4
K7Dm9reZo3cDVrrdIUcvWjnlerB5QmY4G745zfWkuay1ZS1v5B7IIVPB+OblapynCwyWb9oIbaFy
EwXOcAAhLhIwcrYDU9pY4C4jkqUcRE+lvqCe/WS8aV5HHaTEzvGXV8GBU+j8cZF78elsfP8dThMf
ELRIC1Fitwb7cpDl8DOtj28kiZ/yhKvzY5O3RFtfNS1QWTUVzErp89YkXfwKrr7uXh6GtizL47vI
rFND8ibG6X5vusVL98f5/WQktuy/q3tm1NeD+O5MjvgEJhXvj7NZqHmKeHceUYB2RsuV2vsTdidn
/Vk6dvpmzwGZTL+F0E1Q4IJ/sVeibofe5GP+TlEPKWsHCHjDlqza1ZKucav73lUb68Fxvmj723Om
rVAnhURiNPAo7qO27GoCkSzmIhmiSEQxxdYOGhXIvFsQZ4IMrQW2j6Dx2YmWnpdWekVpZhq/Hp6R
Ml5BsfKWrZGmXQvnyzRO181AXQ8+iSy9knamMrkO0QltDw/PJzLvzcjAYvzwssSd3pxDXcNG61zt
5mBbbbPPxx8jZd1z8MDaZtvnIhmSFJ2TE6R9V8KEHL0SMcbhWinK+6JSqYd01B2VGXIO34/vJYH6
bRxhp20S+aYB0KzFS7kZm/yOdvIqiwNvO/gYiHQbZaAagZNrv0XH02UA6+1oSHOi3oQ55pxdajw3
gw4HVuSwaFjwVqvAODyHyYpm+838ZkWB3qew743kChXMepLppmEPIAvsR/KDjarbRJzFXEGpeOI4
TGulyp7L7RP4rMu1KRuyRzQQZUzJ++1G3Bqthfl1qcLdwD/iudlPGzqmO1cyNkaJ5aVWX/RWwY8T
4o2CakMDioB1j0jAQelHKPD5eXSsb8ZBhtUxgITuJPBkQspmYurga+X7gMxMl9hUGHs5webzHP0T
whUmOb1OsshV1A6JUzotW2Q9u9oQx64QLUwy2oRfZVqJgVBGOmi92mRTehyVCgl9Wpvw2btoB+Fl
lOEFppyb4NBpzfBQFNAtMYtuVmRZxBt87kT51kIkaycTpRoI0Zn5GjL6fXh90BDum64Swv05U7Yv
LzrMNNyNKT/Hn2YFqp9Wegp5Xch1GuSHPKN/sdwFiF7IAtiyp+fqKELWMsyH9mhBnvffd8mTPVqn
yaBeWRR/V4QykRYh5Mh7BGCXStNMiJjNIh7uDu0ndVWWRASn6nAxrea2D65/NLHWpUt9oP/xMVM2
HW6/3Puey8yE7X0ootORie7Zw8n6jMaFma+lNGEcXtgkxOy6idCCuuzJ+RsXgpTRFb4g6F3YX4vM
aWiVakQkUvsUCD+iWpLFVEd7cp6JmktQXg04Bcr4G3P2UcBYKlytrk2+SvqW2QTdez9SoiGSV5HP
UlRSLGLF7cZLYmK50riSr9ofq6OnJz5EtnOkTSDAzvptRAryN8fJFp5v7T3j3U7m4oBIpyBvn8+3
OINryctd6Y/ozs8ckPt2HgNb8PBKK1tA5FWgxeFz8jZd+M4TF2T2ZDbdlDiGrDrkXYp5Gfoc6dor
rh0V5i6iNmRlE/PC1vEhyejjMOgVPkZ3/e515XF9ZUZCvwOnd5/+M62VoTLmD5yidf+DfTH9ZUnC
rgw7yfOxmv/JMaXcutbK7lwi9jC2jbOWJiorbfBUSVURCxtNARlLTX1kvyRxgsPD1wpqXWhmqTCX
bLiGx049BDOfzz9eZbUZ8kFFYJh3aDzAMPjssuQ0p01zPChw7n6/g3oJf1RbPq4sjTnmzKulcqEr
EzSIEfyD3Qx8u8U58oVusPTqGAOapcImbpq6XmWm5VYHHbdMfMPLlX9vhbKQ9hU4qVK0M0lDYp9U
jUDuO2Y/dTUYl+6KHiVdhqA9D+yt/LC6oJ1YZI89SUb/Cvcm88v/0qhs+hQA1+TvqgP8EDH3y3lV
zm3Aniq61D1Jjld0DAO8BGb2R0oj2j7I1pt7qhJecOHNdv9Q85zAig+maCYYYFr4NZp5Jrb9dfPX
DGx25NBJYHJViFi6lYQq6ABTWTz0E/2715pPYBLZQHWrY1W21kv/ynC7njwRwVaetifPxbCJNKPb
W0CqXs3RBl0/yj/JLnfmB2c6Q36RRhS7R6tewxlSQxvkMjYWhTIK4rw83TiKpDLr2jQucej7f8re
0/xbcyryxb9CJ0JJwmi5Ik37few88JMpEtcIet2+8bVKuEOArvQBvyKMdlhQdQK+SYqzMQAd9chL
Uq9zN3PH4WtvTNZZCjR8uDK2PCVV29GxcAEpnIamn6699VBCB4gywuI68ZEYD893mP3tNeGRiGKB
3abnrZgawcBupm2aAOJsgmFFeOG7hcE9sfEhB73U57cKdpC8IuebnUnEH7BQyIUEAvP5RhJ+htvt
Womek9LJWrLleLAHWGzNwsiDFz0VjFTSq9dvKVt2QIbXUVQRw9LGWHNvzrJRShUeoysMXXGXbpQH
JRN+yDZ26jzvat4igEE9v7IImk0XNwTMrpeIH+/K9n8ddiWLZ8EN+HEvOR3R9xLCAgRPyq78r88Z
p4/5BzHAHCM19PI3DFPxNKIfL4Zxusf/LTRCT7kZ5fC6UGnA1KjEQDBs1VxBwYui/LoEOCHwK0KS
Aplawu5ATjCpkMzrLtj44j3rSPMyL0NOjBOmI4RFvn62cp7mWm5jYVEBHmLu05T6OS6PXyMHHy+h
elLK4cSmO8cV1k3O/eIFs3envX9pncNmrcfBPvwZJ+jHewafuanaRw1h+pxuHm6F2PNpOiThKwRM
9pDjw39yrtQqU6ZhdDfY4x+n6sd71XB0hACMwFOu53RYwju5kV05MJoJbrATjgGZYbA8EohyAKdT
C7+FP/SDvfSyzfX5DDVcm0k/aLh0bt++I+GdOGlDUzQyMDatoq0/IWJrdxzB+JsRXFincv+E7nAV
5+Al1zE2dC8GxRN0xemvLWAQA6FgVo0G6zwpbPTQFGf6VS2pxkWfDxc/rKbqJPqP10x2s6YcY+y8
ARwIv4NNOyLDen3ElkteFOGNq08LYWaatkf4HPQcISCyCCgSYOVbwAXI9kCl/ianJJJdp+qY0XPW
ZTODjpEl2MxihhgCAhDLmkTvZewDcRxRcYCeTMdiEq8UFG6Vv4BMslKWfxNRTFHQVj0StxL8sZq5
kzw6Dzo5cQDLLcN2CB1vaesoAgSGCKNwSVUvCI5ypdd3E8dTNnA796KV9YtRQ61C25rrNSpEjgl/
gB+8vvEhqYkXFzIL39D4JNq2/yaadsuH6LtzddCO61TIfsyZsz2o3oV5FLbKCJkWLAXuy5joKzGB
1OArz6bXNzTuiVMNZs/lsf4iz8KMYhx3YA9jCkOhY3yE7icHjz4xKrvw0uRzPhR2Tkf1hnyZuaBx
woYIIhnwLP0/eBmYkjUj07gXTknvxC0rn5xNTvvrUB4TmSH2AIQTIbftFuu6a7cnKp0xtTemqP1m
PrSGHGNwgrYEUwNWdW4UwptP2V+Hew/5AfLi3MhZbKYDmKCrD+aTHEwmW472CJFeFjKhcKGhy9qk
YbzPwnPiPgp94BePziy+CErHOUy2qiWjupBqQYxBFzdrTqOVocMiEqQqKEHCoZJEJqJTAX8Wo4Oo
RFZhQ5LI9/hOgJB/Lm12TFVAyiQz61/zuJDUwrmxOxGPKGQ9Wt8VB80OTs+o+ZtXSWK3LjtaQEjd
+5gmU0AtbLrW+QcRsPXPaNEP/tprwB7ytkc0+6S4YOoQRgcMo29galm2hsMDEuvkgRQctyFoOhlk
2ekr+g20jH35uewLkHf+H9qa2uwbTu62/4WxGY4QQD4iNyUp1o6X716xnRGHYECpcN1gM+/itgLK
ogMTSWB0d+M3GfRe2lpJ41ftaGsnZ/qagMVYHAlg8DZDpMm8t3VpDWdg74qB+Hkjkd2QGv0xY8Hi
92qy/q7i8ASmxLNZqOAQU1sWIYshoe3lLUvnCesmv36HoXB7D7Rwl7uUgLlA7DU6xZu8mWUVNB/3
a57cqzFIzArO0LHVAm1CQI/yc+aE6kYP/hYmLcC3ohVLQzQjhXV/KCImhjyIPeLVH4VxfTLoEmtB
FKbXRtwTD1inXrrAh3urc+wp29TGbThKWLtHMYzVweggi9M5UEfKJArbJ2THzbHA+P48afnBXS5M
vxfosoTkFFJDIF9YScwKkDFsWJNSu3AvpxzspFzsNguwfN0z2jydb8B5tQgddPgX/PkkHmR7xCwp
8YhZ6iOyQW3vWiDC3Yz4oOqo0i0PP5AcedclOYpo0JMyF314RtRCGM2U+fqzUMTR7pqx33uSI62F
UZOMp6pmnEuZnYhUXmHxDFjKuBXu0bij5CFK5WsctAznOoY2fQ+lvi2jiyxG+OzXAqVJgTra35bE
OWLfGtwpnv/LuddEgeEhdba/WElDRZMQjw/Oun/3PmtBI2Ahu9hh2B6zqnAKlhbLcC00+e44kNaQ
XP2AZ+PlTibv/egWctBvrHEevTNYWUVJJGmPznz4m72PYNw9nMxQbD9DlzETNskAmD+tR+okvekn
tVGLwbDjnfFazEaZC+xo6gUSnvK4HgLz/iJvmENiZfmxeiZyWX83Bd1T4dVn8XQ77nnH6wi9H7C7
0u/dJvwBn1fOk4G1aLl3kIU6W3JMrZE53AfOHdy2MyP1hAOrufjomCsWsy5qLPrJeVP5M1YG8qLz
L8op/do2hOLdNPJtWWPPC+aNkMccZkCLehe+6YZY8tnPxzHHbkq7JQzBt/PBC+BCNgZpRyPdI+4X
cuh0kSOgb+TNPVO4pNsTIVnKIltC20W3qFBwHLJo7bUsV9Tvit5X/Stm9ACjU4mVKgc9oINw0TFX
7P7dinO7BSi551zT5JE3RgJofNLRvrZqq22hG2TgRNx49DpbdxOLLdfAKpt6vTrbxUkrhi/lULs+
moDYy+fmH+GYHgP7iYOMPHNokWWAtnn5kejYFBxCqKmmk+cJmo1hWS4iKZBY32Mj9+LYvTk2GH1h
5yCkzHHx9DPiieUGEDCwdeJ6uu6pd/5HwgMDfz5tlXEX3TRkvybXLKHS8pva9NCs3dxg3eyb4ons
g2WQPf3DhRszZ2o3kdungK6AES780Q6QcgKcZO71Dh5KetU77qoMJSn2ZpdATcN1aR7rW5AsZQxl
tfbW9/Kq2T40Qcfw+1HPcBa0LshqfKmUcDE1qEOaTxsE7dMz5C1SwspTXFD8v4wEyo7BFyg5DZUs
uAI/wMIL7MXG/d7cQNLff+Il6ZVClGpo2CPI2zuPk2u7irbXnYNa6nRLukuZDrGU91evXx3uygGW
1hMtNGpDEE+4M0OBZXLMFvzk8IiaxsJf/kfc8pA7/mYgLmr3OKUEoXBqOvTFHmzGXH5+H91VVxCK
1kFL+asXpCDcNqQyG2yvLUZ4hpb5dNwpin0ELWfJbySexInvtOmx938FqKgQQxsqgUwx1lCWK5Xr
bVfDsq32QHKquBld+1e6taW46qnyXEQKfDgyTP3lfoYwhDzFzng4XccL3GG7b3CthQreG7oxSYPB
bJmRrsP8/ghGPlYheV+g8nnSuKpG7590N1lq4GRsHA5qdNxFlc4ZR9wfMrCY1PApVfSjj3IZb4+v
jUCMftNJj2rXf/dQKNqXLr7XIrk4t4mFGwqKoZfXNEt+jHXGkecmWAVA1K6KFusqJqYIDug2XXST
IyQyLW95O8SSEkAyDOQfRt0TLs1CEuNyQiHDw8XMzJXiKEemAFgWsX+CX9K1zCRveq1wA/vv0biX
T4hJ5duYn/5bhYH1P8+bbMdYllQdKVCZ52dja2yDkrXQIeKaxhKyB6ESBFAmJQtQUFUEaEQELh/9
jok1eZfCcFBqUSyNfqWOVZWUKDKTXJB/37BYO8p0iwN1xUaWG2jv1vUBqADNT7eOafWvexZJIz39
pP4GQP42MEttMjKSzIPpniB7ntQH85sJbmDM9I8EBDFSzgWYxUCQW2xLFz2v7/t3nufqt0NMiLW6
xVLOkfSdHYi366NIzlzMCws1gPECsAnXZnT2p+Fpk2vWgL0icwqkNi9qypzdCIk5hxH2+VD67xhn
F6WtpLQ1SKnqWW++d2gsnD3/HZq10CZjr5S3cA46brhY7r/4VQvKNY+e0dOTbZvIOfcUuecD+6eN
gJaigiYlBZavD8j0kioJ5a4C/iRo0E9hMEEmVbQ51Tc4usez40tieyvngxGpiYsCL80fcFPjAHVt
niOskEKndNyGG34J1CMohqAde4FHyFvB0yk2VvWzuuCzNEUFwVv7tEcwNS2TUxv3aDLYnSB8bZya
9g9IZXPTm5Vunn03RRB6vIwfQYYVk6OItn0zytUeJkaNez1rB0pD0E07hLEkn/wmVzZGoljJL+ac
FdnwzqJB6uHjBTC1iutvUXJtAicee9rY/6uYg0KzivJvUMRv6beLnMXCA/isKm6qsIl3FH1VbgMG
VCH/FTkGlhYhG18h5HUu4cTLEBPq0zbfZHpRJGu8oEKMPwEAqsUBlMercAqHWhAYJ68j75PD8lkS
IdseTLxLDgbgC4uNOLrOuQvVA4to2KwyxdoKI/W9LTiy1Yui3PMSn5U9l5I+LQ7AqkvCrrHVBN4j
q19wNDgRznZiFiss5/2YrBr2DGdji88vCRAPiYzYbs5JT9Dz2AIts/UBMuiicfElPTYhZug6Mcn7
QIlNRecoKXT96d9L8T3ccc1h9s5rcCuNT2UzV6uiEf0ilV99z3Cql3Gs8iiO3dFmj+urLMwevZpP
DKnhBUs1ZSgI3J88opaZsDKHFrpYR8kHIrdXujlqe75Dq9DJmZzH66QzVjWV05FBsZnIUYWpEDP7
Rvvcu57Fhl9wbxlWkBmSsUzzo8cmiz7xt8n5ood98fh17b2m1YPXSQuUkJoYRott5AXVmewe7W5M
t+xaRwl8JV/w+LHFV6KXGGdDM159sAKVMWn38j1GcStEgRn6B9sOjQne/WYCgemdzLwGZH4Biu3k
6hRxOv9I+sflxW/a8wbXmy8tiFFO5MkuTqkQdxxtJow8vBVDPfhD8Sz8JeYqV45maeF8tJNMovbi
Ra0nIqY8AMQyMgHNpvjCgqRzz/xboqcjwZ97dx/GQPBZUA55uSAdv28+oXAxJUYovDPUODRqXFPH
QOcLOG0tN6FZUxt5Wkbz01Vy3ZK2jDpxpULBGMwFusxoBsNM62iIA+PF3eiCAlY8sf6xh9OPX5SU
QO8VoMuPQZvzmPx2qGb/F0Nn1qC0ZrAcWKwcFrrJAyrvd1QRPswl2sXQh3JyHK9iVKb+xD42DxoZ
WT1jY0+vZxWTPQVX42DzqPvelZltZ52TMT6Rse/uy/N/y3HuSfoAiiZoDiubNVEFCUW9tsfW8Wt7
FTl9IULfsAEDcWi2Q7riL8QXn8/7+znk5Z+taavnTCNMPbnmN8Du1/P7LeH3y5ttDhBftCVuksia
Lh9ng4BLI0akjNQ4PqYIRWq3OffHD+/stOQvduVMaH/gUVBH3Sez3byJOSPUaLudYniYXOxE82p+
S6hH4FheYt2mhB+Zh1Tm7Qbr0DjvhIwlzh5REbbnOHLXcD2aYpyG53FucmcTPtQsHNz6KgK4+eUc
1I8lkHY7LS+l3d8i8QjKtHbeNFayjFVimthrhKExgIMDGlpkFLsjSavGo9cQnujL1U4f1696iTWN
wlOHx9+9Q8B+kFDVaViF/LH800wQB8b897LoFvN8b0/FiDOwDudTPsWcw6Rpiatg3+aAbkusrD0X
PQMUafqUPxq152fyssTKLTWUlmxobGMOQVOKjCvcOtDcb3jzl2P42r/03OdHDSpYpmp4M3iOfynQ
FQtj9I/jQ8aTCEiyOOBC/iYZzSd9/p9a8c68lhL1IrW+f15oKrsl+TqXyZ7+GmTrs0ADM6gpfM0A
+D55O5SzbeAMFMRk22UEIN8P+Fw1GcxHH2vEgnlcSo8nTqBuQqO0u638+tgmgSfmrNHLTEp7N7lr
kNOQhHX2jvrOFGYxrIhAbXYrUtsYjYi3Jlwsh+Mr/tBBStJ64UBPgCDBMzKta6DYyXOFmgKerICy
xVvUL0nFhwk/+E78+uM16fgXMeRkfovsAhWRJs7vXKaa8qLE43P1tnEKP6Fj+lSc8XRm0rz8befL
HzY+5x8CZK1ICEZ+Q2cbJhLnCBaxd9EfJ+doqpqz2zFg3ZuTUYeuYC7LXTZ3PJ2hreALeafZV3QC
qw+y84Xldh1ydCFTXL2VA9OUjqDjik9Qs+5u4Uwtg5MSIi42QTEycdKtMUbOjqexwmL1If+2jSRT
QiQK7uYUohd3epo46aiIf36aMFGdBROSDJ2W0+VKFaqfSnVYj+w8VnkMth2uV6onJUuh/H1N24rC
/10+4USBgsAxS0Ru4egxfJhJBGrQrph9vNYNVpUuNRiZAH9QlUK/3HiPsboWh0bPaSX4VHKQ2N1I
fUAK9BLNQP+JQWAHndkdgg0QqNDibQoGl+XaRwAePkUz3UrzV7wjnWq1Sb2vLXE18qP9dKYfkDPc
a0n9v/U/Mv2ebA9EVT6NytnPegCtgqKx4AZPcipwQzPGw8uMYjtPf7dfzbj7+Y7oqdQZ3n7xKcSu
W6MwLd0ty4MF3FkIbqbxrA2eq9uD1N9kF5Ah9O+2Y7iFpG76AiqsEfZWX5MwCB4q9VO8Gige8OEn
eBBFjneL3VOGPrfzU1DSOM8oB4RZuohRKnED9u33WyDYVbxmxzArCGnPfyipFR8N41ncsvkbqCns
kMnDX/h/xNXo21S/4bpbfHfOFteR0wdeOXl6M5xh0MKluYIgaRM0Tnq0rZvsPjQLSLh2cjfrEbT/
Wa36DTzoR33m7Iqua54ZLv7NIWWU4LWSfFvXSvg6UmkAK4q6kFBgRrZsFX4i7zldJWsmwX/cCEaX
RI4L6yUT0cY/m9hNVbvydeQVA6ZCmuB6pGre64ZnGp/nHBfQBs6J5BRPhrCYO/ar6v5PJY8ELuuM
ycakNUGx80wTQ/aJ08YB4FworkJjdP2HA6y/3UMvngQ1s5FEy8O9wcWGyM14HcwY47wKvEHJcR2k
HCfaZAkrxFzk9hMvm9PreQH6IxvRGE6licHzm1Iut6xbJD9eg5Ksqs46XTl5DDtwprKyyv7SHZlf
AadP819uTQW1QuNsKBb49eqAN9/MsIWKqQU/nJfN4s3LgQsPeFPwZA5JihdZVeFUXX0ufVifC043
bNzudKInfydt7a1OLRBQ2ial4Dgdvo1alw2tlFe7FfcWSgd094kLgrv2EMbN0DrxzAs049NQJ1gP
2s2z3ZktdU1+FjnL8sOEaqIpsxcH+VoBMmSpkurkDpgbiGRleGWmcX12dlCO8+ihHJTHRaHrPE/b
E5rRpy1I8dJ253SIBsYhhcKKiPfzhRAM3Wj4afsQJ2/qBqsgm6+eClNKZFImQm/JZ233zbjQvuIO
kaIO/lHxEITSvHGbTqlza48xExRN+tWtD5tJJ9I/PVfCd2yU2qwZuNULrkR61K/Ey0BL5RrTuBg8
LiywBzdibqbg63586xundV1UXbIqg/vMZmi3JKWriwhD0KUNxJ2lt/DJ52Pb37ADHV3kcZZUL4tU
VgYdeDLnXw30bY8Pnkymh78OAU+xYEexMt8u66TbptJS0U21xASl89PfGslY2yGPUYOT0eFt1jNI
QTLxLaSsRNlmgrsuH2DHLQtn0txdFrriR5O5oECE7sE8mZjXJCLWrU/mtmTTkbYQWb77YWdDbiky
Qpoiw5mN4MB1T4QqzMtaXPVWrWxZdSOkiZBoQ60/ON5Gh3s6evhexpLM25X7b/7yiMQ8zBvQ1Tmf
mFgXNVKkcO+0M5fNnnlESbltc96O/ZfDGFLxtionM07si2mKuyOhiSWR3Kva/26NrpaUD2Bv0gQx
Cd9op3nCfeKqyWRNJd2J09CZEBeByFTO+oObzCyztyNcQh0aAtdGZoIc+ozHQwLiPjov7Xt6CUH4
zHc2K2Ts53o6ZWQ+eJI2BojgdGBlLWKvZEg8wMjEz8aSb83HHhg3l+lGklEI6dbza5GPVVz0Y6g7
e1C9u06AyRMXQUMsXYHzlO+/qxRogNBD0ha0rDRLg/vhwDlpRtHvwZ65tEnr7ZruwdQav04UM3SI
I+BM5AbaTlvZKfwoGbM0WJCAPtEaJSOlRrVegTL8J3FvK2n9C31yKMK+LjOiVFMVeNO9kutBfCB2
vUcw8YqmtUYPh4qJknyWPadLH7HPpOysbk4uTP6M2L4tIWAagXfzXo1MELltLUcGuhpWb7EVsefZ
QWQ5Z5hr0LTfPiI/IceCpsBUinKD1+SeAtcNqH+iY09iZPN4RjliGwY+P7P2cR618t7EUNYULLo7
x7p1k1FlcFti/HaKvw6hJKKzHGMC1oZpo0qFPZXSEiJvOtC7rnUKvGwHyI+ZE6mDC3lYjCeU0WMB
fTuqMz3vpnaM8/bL28vM/34sIShbHBCC6qaVjmgTX+faIQyPt1jc8+P+z1yINq9C+n0cvCSjfVVn
C1H4/2xWZsCbSWutixd42nTCrtneM6xaUcgEoKlkXyvo5lm/j7jXSfShzaCUwDxorvePHZObs/7X
kVh6JQx9LRiKZ1i8UnEGNBnci25gfPTv9mI0Xw8/Sfxrl45fakkE4ap2xdqIuKuaooiYczQfZPdT
+6k/Ck5E0KfNlUpj10pvLYYvQTwXh8hZD6tUHVoS4H6e+dYibMwOW124uHEXlJpbPJ6Li+NXEVqW
ivYhNaPEAjwSD/t27gi5o9+m57DZYrOr50Tzn6H20IrvQv98XXlurmJsnQI4hwZEcKINhOwsdkwl
XHsAOiXin9C08EhBomtl9Ghspg85ShhTD+DRdQ+oAEeO2CT3QmDDZwBS9DZBPOxKnd6XMTdX4hF/
NfkCr34uC/N8fzTNwEdoFKLLEgV0oSqyvijz3lgNpkY8fIS1q52Ld4FwQ5OhaBRRmFusZ3jHBJuo
XkGJrCjwSZ0KgC1IoGeWbk3lL+x+Vt/CyFgc28QjIXaEqQTP64lpwcPGgdGaUY+8WAm4ofy/p9L1
aGnB8x1HEvrY0NZq/zpG4OlToXhweOtQ1d7FzAUFFTbK5U7dY0cWowFV6A3mQwH/UxmmZGfVuEb0
Sl8DIIDahRc3MZKWT+avvdZ1QXtpjU24NB/LqNdxdZR75tjzaFjDDjtrKz6IFLFu3ZDV6j+ehkoC
Kcbu+GK2715cFY8dC5nuMEV4UXdJ2Z9flt8lWTbFrfrqtThdfhMHXwu7RBxR7hA6MCPzODrqX4cP
dw1LOSvb92F5p39annV4icSgnvuz4oxGPHosKY3vhTNzd947LBMzFiVi4844LYWM0WiTzvCx93Vy
YkR0vRgx8TOG0wfSqFwoR/g9ZmKcWEI6bC0gxHDs886XOIBzBfDsE88+M0dkVuiWjwHLTbnxAKuz
whGuHY42BFzA89/HXfz7Tc4emXsjkHDKXjgdodUfpBxDaYdAchP2/4sbGk7RwvAVa7s/whkyKsjV
T2OpyWyih7j9QXDxKF5IOF4kZc0GQq5rJQEnvCJkpTtb/gGAG++E0gGCsdDiIEUVIvjZtH4/76PS
FTOZ9QRTlvp7BBIbzXBU1eJj3XTV7QbGSvW/Dy5+DjJfXNDzL1FAtxGF7T9a6IcUTgmzn7M/PyDc
9lD/0hZvYnVDZ2+NyFWO99KnZoCY/PJFnFlgayZzS2wvOP9SfBrGUst/Gr5b1VQQlC84WtrgzxjU
1/8znOUPJOSgQF6DIDl03yio3LwOOrInSlYW0oGzxRkxxZCuOekebbTCBZjg6hIPkIvid1yhjvzP
aumrs/BS5q9/kWT2APk0SRdk375hN9g6jLNSKi8+5RkjWlCtW6ktGiHvlkp3EFCsmgIiS+4bp8kw
5TP79/udeIXPfORBGzwgkYq+cMo2rYBK67YpTDZmmIf2cIz56ElQFSDx59jgMSxwDh6+JoD87OCj
i0zNKc7977VYU0GdmQLvkwy91ubpoVOrnA01tZnWmyLmEv/f5jaxalPeQD1aBP8CXPTFRi0J4u9s
MM0hQ6t0q0T4MZQOnwrqPw62A4UANUraUlyod6m4dFFu5a13rDKHl77DjT+xy9WFM3r2kobvwSNZ
k/uPmQ8GaeJR6audhFgr2e/fLHLk1n08x2qKodv2L86tXeg/jUd1Bv5Q3q50j/uwVKJXCDhJmch0
qrcyzgCXQkzq120Ehgzlybf58C6Us6M4tn+j6zl4fIrNWsiGiAjEz5bULQtK7Za3rfcql7lDx/Ba
T7g6felVIXFSD8WDaRTrmLj07EuFvjnoJOc5K54WPHcOUI4ztdKOVK3ycqJ/jr9PNV37AD5+aAyG
XMD2aEgQY7dKHnIQhAVZuerdXjTlEjOE/bGWuj6v2XpwTnXjCA3Wp8TfKUjAsGaJewLIxrNWapy9
yYNJy2eV476MnwBI0UojItCo56hdOcWTPsg/NkoNWFHXmZtOSyUVzXTRhhkzJnDotbvNYIM2PHvN
EWgLtK8nRKcWMhLBKPU528PW2iWCu5/pYksLU8cPn41ESee5Vcq3chXzvV7ASPb5zpIDYqCYyt6X
JeZ76sDAbJeKDATb6YR/ykDs1baBL3Rf57Ay4oZ5NZLATx1pvFA8MZSi3jNAOHi51hcje8KxYZR5
LRKhk0uaK4KicgrcuEL0SIrmEHqIfLtg6SFYXWhsGi/NwblRjziI/FSPv8iSMLaXmktmOmAlNCv7
WwufMhm3jtRpMMi/Oo1NQ7f7oycqb3PzpponfXfsBnBSv0orSrWxtSANSmPRHkzlbFoWG4wwf94G
p+HQl/hSspqogXzlwWEwaF7yJ98buhO7YKe0HBoC47TbPuEMgk2lX5NLrkbHTzSTRJ31zYJ45PbD
A8SvAgRSt/7bB2gm1FveT2uLEQZLx4VPWMLUb/kHFxQKCcAcgNQbNU6oL7XSe97tSnx1AgRQhQ6r
wyKVL+TAxUy+bEC6LR56yjqdwwV091zVFtU6wqYRaha7edUUIiX3n5COThd/KvKB5dAKTim8Ifd/
OjlziNtEHxXWocDbDAETsTl/JvjmfhKZfrp0kdYNYfUOXa55O9z2hN6Bf6X4LURkmtiWcxpsYE44
bW6Go018IR9IAsLM1/hbUvjUYIEWFm6yUTEy4oaWwtnl0shKnzIH1Ms9mXF9XHCOsnW3lQ1fqJZv
SUlK/Pt0xk1y4X1TWW9kWWYEoEo1Ht12zDM7QZQ2lk+Q5AVJ6wth0Fx58+ANBHYyY/SKF3f2+M9l
8TnTDSh4Jkeppe9zzT0ymZQN8bndzLGr6wz+yfY2mdO9W/6IgYBbGmYIt/RQW+lJtFbKMxNBV7Hr
XHmGNkyCG+bYRitHjdzvBSZh8IbI7DttGBS4EzNzTObMX2mretWRRDboAYyCx110br6NG7a7lfWD
HSDqyGeMTl1YJOv5H+khFifrL2DxdLCctbJqWx2S/GgFooTgKmABld6Fa73WTx3yeLEb7O+fpzEv
aYSYnKzTHlOM7NofMr+2CnV+lCUHx/BHyImBjWLh4fl7/qSmDoqWRQAGjsdW4nxC9kV+QJ4sFo1U
IL17rBPgtcUAAlLD0qwlBz7FBmIO+wXiGsFkbQnOtGvHyd6P0WylrrfdE5RRxbqWdkMNNUfzpK0b
ADLCH88ixuMbLeKCcfXRuZ+t/thrHAkeF0IZaqb/0qfqFVERSfQwNbl8gK8Zhcpi0DEon7sy50tL
YmH4yGumf2lvfgzSAnKF3MFaQLTnEh+7ulvm1DyTd8W9OlX/P73rZU3P6ZnkrQ01YapHBeFHtGDf
EbvbnAxp8+gZc+PRwfphR8D7fZPj3In+fXtnx4qCVkyCq03UoW2yJLuRxE53EQgO3hYNHC2x+Gs4
NZQCYN86lN0n291dlPahUlD9BUkIpztGZV7OgnlZm9b3ox7V8KJO+bjjdbBSCEy6a52k7i12AZFL
4hkz6kZlYnhMFFmRXoJxPbMCovAP3LZ870zHOj9QExMKXSoswY1n6+dyzf/dMuaJtaGPKHPIckcv
JmW1EbMgJf4pGrzrqGmB49AAwMmXs4JdhqV4bpX8oFva6L9YXIrKAf/egMnXl9XAp5uCsAQK/k0G
jUz89v84Cc5qIT4fMtqkhkvn3m0Bp7DXaARCuhJh0xnhxn5KP2nLbLJlmZeS2/j7gvN4qNtHzW/Q
4yceEBFFrNrFE7BLai1GlnJA4Z6VYreEzLKus3IkaFDx+qTJopOdp9mf2d3Wcew3IuAIEVVzeNSp
tb3j7YRZcSXSgAifVRiM2B28lfhL92e6ceeM0skHPxeFlluzFAulOnUxaImqheKbtx0dTkAIGzWF
0FcY8DfIiKcO3jhqCBombNOEtIyj+1NvgQ4nALeW3ML4+GNwFh23ORMw9f9sFQGDdnZ+Iw27T/0l
rXO25eriDe082eEvXhBoR4Z8n74cATxA7sfr0khw4UzZ9UDAB0gJPSnttkeuZVGUagJoJQ3yxb41
U6ooefIMGTIhorTyOjW03/N6UhyW+xiDX5Da/F2VX8sF5wXFL53+Mu68kqFmn7FUiUKvZXNlGeoY
h98q4HpLdvQnG0Hg/fSU8pUpTK7Wiz0UpbKWko1PpWqbrBp/8cxFnnEgdLZldVyma5SYbwHyyA+A
mhOjPaWp0msG+ZkEAD/32IJsyd1JcRuRdZYQklubOqyiPYe874cx0tS9MOHStYD4n7U9HAVJ6m8c
/56BNwhQumXP6knG1SkoFbCJpt2x35EVbkBjgA7r+a3aoJvbyFw11bxFEOatDZDmj2J3CQGtgpEF
hdOW0nupbtP5Rzb57KEa9a4i6Y8ybndUhNLG2CV9oS7giTKTljCgmnDjzBxSEzS08lMEtwFPwOFw
7hu4aK2HOHhjMdCQiiFusBlr2kFPF916JqzOO8+jQKBbOFsWWvaL6z35OFoSJHWXIRXvognFSVgY
ZsMGg6Urw/ZNhFIlCKsI6rorBluUdh2bbto09cXZr7e5UK6qx+O4+18UDFeP4yQI6Z2g9C6DiKvA
lStgue8ElO0gwX5nI/iKakmKd4sByX34iezDo+tVW+EXOIN44HcNwl2KgjNKTmd9FRer3QgDoCO0
wGsYDOUWk6Pd9PvUX6fuGi9OZPEbpDu7WgPv8SKQ8P12z11Gv5ZBH+QSHq0kikr0FaIyqbgwpPyB
jK3VjxSg+vGXXeMv7991Ic6jptwC5rFSZP2UM/RD2DEPZ1j8ESbznMPrFJllbFJ0sbLJbkjylB8h
ZNnJSCREEKFwlrRZ5fGHgrtU0pdUa26Pywmt+LQ5EyE+u+fhdgzF9J0JFatq35mR/7Qzw7xRjb1q
y5/k72Tww0ixNeQnxVqWE8qNN5QbfaKOz4z1NuMqci962zWxUQUqWgyhxgYebVzdsOW387BJRP/K
MfVi4Vq7X9V3kCdC2gwrHyAhe051UGve6SD6I4Maska6PQT05siuBVsumKpEW+U3EB34VDoBDjbQ
LIc54cEMDyEQjniMaaqjCyklFU44F9Vflsf9XlfkIhArSH0FHRVxLSsUm5mZphPzfootbjLhfMMw
T6JQz2LiLCRpOjxblHJ+3Qr6irtK4mfsduqd8sHPF/We08aOmHWG+TOaQ820cElpgUBOJwTzN3Kc
DMLldEp8Ow3SLNTN8ayFfl+rPEmIOFAF8R+vF+Ze7+DyIcuTtmAVBH1W3A187GeI3J50xz/MjqjP
48JTzbi4eYDuj6mCoqSzrPW9YYXMopON163cLYBHAcfDri9cHco7OmrNliRWfZnu7PvWXXXF66YL
3CWhioPfvTNAwiAjTkVfjiRqvWbgYd3LGswm/i29azyMsAV2TkMFkc4GPYziQzk+0acsBsry7mgV
C8bAokmlE/BAtmo5A3dzZMuGmyaaPpxlM1SWDYHHHi+uJWJHnGvhsubl+sNY1cx5KzJTQdPYJUIc
EVSlE0zwJKLG/ADLkbXtslaPhIS/mEz9YiqiAiGvCD7CXQ0QpWZCD3+b7H2uIcE6xNUVj2Rihft9
7YvYk6HmFz9VGcrO2j5Pr85M4zCqKTsvw++8Y/ygfC44UlGK1V8xXImxLsBXJVxTPRc3OtNOxOJJ
GwEIOSDqWnAHDGBQsV8nnzXuS1KQs2kLOIMUrRuidG3M+sEuU5arptfKsE5tdKN873V+mC2+yQc0
sYyQqPgObtVn7pHi7ssHWLZtMxkAPHKK7RdyeY2vpTP1n7P4qs2M6KUN9iZXPoWDZbWnn7hfWGrN
Din1Db4R9BDz1WmUPWfkjcW5EOdtO9UcZiclgerTxmImVPEXM7YFrcNwdyFTByjs09bH6UUmVWFW
F8r19pfrSOEw0xMG/6XjHzpc13SAR6vGznfouDWBrpCjojKGivLb3JOkgc9Il2wcgvXySd7RHzXK
oNWSOlXcbHcQs/lVS+o4GAQsNx/KeDBA6/pTqLYkqgQD0MZFfOG4g9qBpf9zirlx7rl7gVclrfSy
Lws9yjlvuAN3LfAs8/+TuspjFmbzpDm6++3v46ljORiAx/pfi8Z+X+PPRxe8hPC6Bo5hEtFJCKL0
jKw3xLXli1fPTF8vMrbeLaPdPhk8uZHdigc0wjOs+reDURvzeTpxVeJ1M0OAf3NnNoSBPtFLZigz
2InHv0ECx8faWH6Tz57m+cpPD9WfLN2ntk9HXPxSdS5de1R8oDpVnC9DN1l1TxEbl+LQ6h88m14m
jiw3YfTwGIc8f1tvufWsHktBF6m3AwMTrViXGTRn6Ug0GscvaroOzq+3rIfNf6XpWnHG5bhUm7xe
XWiaogsA8KLNu2J+rrU0SMZtclbqCbUY2CwgKZFdsTnEzNdWQJMnsXlLggnK8oKURideGUWgaGYh
LQXF53/beKvxeMyCt4WgN7uZGmskl/uW0eCk+J83HSBd+lYOPQmUWqGgXMk8GE9PADdCK1M0GJ3l
aXmAmphnvXEpb8cGECvvKTTt4MBY+UYuhzYzIM/v5S0y2YokTskyDbeENmgTnmA/V1L+O8fG/vGa
KdmkXihC0wk2KngbnGo1xDpysBtBgGwXv+QO7U08UI9WRp1zqGuL5h9rCNkm7jfacXdP+Dpq7o0S
PhgZTaPmm7x5jS4s/JlbX8JCVypB14NTQagagqZ2xE1WpEYl6dHVfInYB4uLSm4vI5ByV/Mz6gjo
dJulOQWDkYVc0T+CDte+DCm0kOiHbAqoogE4S9bKctJGKZMM606GZytjGJvguqpnoc+1cENeEKgO
uM2ISZr96T9/4ROd7V6r+q7mwkR24E39PdF4BLCfhXLMrmwNEc2KN+Fh60GkUu8yR9y+wklOdlYd
5t/5dNq/dfcpcopjLo40uIGX0CplhpY/bEw0V94XuuIckkzic3gtsqTmZXbqyX+CKnnhZpGwU8pv
sb3ROK0pkhl1gKbHJg/Rpbh9aZ+WB8iGLxyVgwbtMoMjhJyTIyV94C5tJDnOaTYaMn6cYg6F9bE2
4oUY5YFgaKs49Q/+/7XzrcuzZqQDAA23ElgPv7uUUPWRatDibMuKpnub5Oj6iKEMzrYQO7ZWBXTx
V8DfXVw4vfKMBrdN0RA25aX7O0Bb7miRIMNOiAu7JrygQeuLp7B+cc3LrxZXxqshDmCVQk+BWSgS
2pqVjq+2YB5FB5Ab6aY6DDzPExC5ae+DrEyUs37X1Iai5vXfZ/hhoRPcKMXb6SUiDv9JgbsDGS6p
vJvnzgITjhKB9mUnhx7NqgwdN2YaMPHeio7BNHZ2+hPiKaYOoQ7/ynGv5ogrTcpDiekS4AMQE/U/
05kzuOcuXkozE7FFzKqCdQljZCDp7eq3XaTA8/4Sx+fW8rEnxlrdJuMV5lBwruL/TkgmJYoAlXUo
Ftux77u0Al56stInt1/aydq7njYy4x6w84dwD/98m8ZClRDZKv3/cC+4y6ZhJIudkE7sVnBOZhyK
E/fVQXmmU094aZ8Pg0QHBuDUZXmV7QP8JAvECr+sa38REJTc0dCMuRlh5QleL3ksRmCfD7QMt2//
vzUSxXCdfaHEOq51kUFe6vgSCBsruYcRV9Rjsy78B3qMZ52bTB4SnE30NBBAHyebjkZAmod96ak2
5rGwigwqtQOtgwtxoBu+Pqiwiiwl68zXR2JtM6niQtXmlGmQjXAC203VzWyzAsFAXGvf8nT9gH4J
hagM51Vbtqd21H46IJKg0Oo7Ogyu7s5oWiapP7ThnKkuHk0vauRsnnJ8V8OUnP4BoAdb0FgI1qHD
px7WMACv9Y9gJoLC2mZ00LzaPjBqxZCO51uCvNv1ITvPczaSYnjjOGwtFx0qNyWc9sbQxZfsMWf1
XWpMvDndHyGJ4qvJZrAxPUTUSWn9CqKpa5zqF2KR9hN9V+drRqdKOT8+SsJkdBxCyeQ+zkScaPrd
5fn16fiyL2sVHFTqGkGbTR+yBOouSF8AR/xH8xPdwANJAjn8yF44DlGcGvWsAu6pE1fvy1S2tP84
lZjXWmyPLGN+E0sUz+0YGv3GKJr98ngVLG5t8xtP0ypQEBp9qyYc1RVi9tBClrYQvNhJBnD+W4ge
c8yx/NECLhxsrh60YKjVM4b6vNHL1yTwW5MMHtunefIP+CxYd5HUt8C5LyROd2Qx/uBzDl/54Y+f
MdrJHOapJB/VQSeBhoWasMJ8x46bHvsevrG7XVxe1a+ZqTduRGlx4wyFIfrE4ic9eEqZe2sjQxCo
J3H27eYYhoF8OxXpxr/XZVsmPzhc2vBl+FKDeRmP/vMg97nySAShGh6cAuVeDLSGIxh8YdaRMbqQ
KsAohDYzKGgYj4cbU8yt9RjC3aEbC20zQPN77Q7FPUPNN1eFM50amSMAUANJ8S4gpKvzZgu1+OE7
p616KEDD8OQ342eKeMBIfA7N3Y+O7gfneaDt7jsVQI+TH9bszzHAwK703NtKiCmzH07535utScv2
GyTstm/aYx016V97DrewRAH0Y1mhbX8loa1P8++Iigp0EbMp/DMgEuNsJo2PYEYUchB2R40S3vbv
YbAaF21BGtR2eYvoMAU682IHc5fwXKTqJpoLzzEDzODI3NH3wibMKieSvGRF5CuBiZZ0vw+Sd0MQ
Ph7L/cISi5ATn8eCjeQmwmUddtkPSmhRaL0EeX2UkzTnZl6+gJa1Wec5cF/y5ZVCK0m3yacEpmXv
pkoZdFSZmUcT5BZCPAjiJO5JB06NoAzMkPotatZn2ZPyrgWPpzBfPDmsykmySkD4mhQrs+HobYyb
6xGERUwhUOg/ueJqQLXOJoYu7UDjHaLGwLlOwY8sDPMJHa8Zias7H2FHaAaNOerN65xgKViwuWrJ
obVhBEaScciF+4D8cSOFXRv0KjnEYs6ubKXhe0x8QgQeSmzxJAXhdwyMt5hpnmEfPn1reyUGWn3D
qc+zsH43pwqysLV6bHOl6sdD8EBT3WNcmbi3Rx+qGjhbNwIxjJbc5kbmHyyhmO30BbLir3q2hbxC
FxxXugcQHc9Q2+U6gs3cF9rq3LylCQMp6n8renMqyE98q/wk89iIJYmL9/+kQ/MBd31vwEQUouLe
l0ZK2mZ/VkrtnJFO8U7ByaPp3BBELopsyWo9IAmrVKjqZI+NGF25V4pdOwdVZscnQbfPltknX+zU
9pRaHb9eFJsjzp/Z0itz1wrqD3iFON1OMw3rpA5SM9zcgLCYtC0xR+KMXIG4tldXIKNPkbXCtilx
RNWM8U0hKsmPjLFlQ5aBRUJ6lmbQp8mt2BuiHclmUcSFY0Ki86CBJ28ttMbq+xwFfq23BSppXowz
O7XfcR9sx4qm5ofVkYdyhV1fWLkYJhQO1ZG+neqpzsHq4ZZxJPL1SSqAAINlKkM576KYcHrJShmc
2FfPAXjKXtMpRWbQhTVsxFCI5C8SKrCWjs2I2qocK1GG1B7cRKzwh1GzFAiKhB7jeEGeeCZag8ON
qfk4syZiiyL01h/+B6t3kfS89eNfBCbNFm+rFA0gdpSTtd1WkdAPr83N1Zm6LDC8dA5E5pOc8NCE
teCDshLe1OE3fqMPlI+Wc107fiJjzbnsEE+9q7Kg/ahTzcmiE5rYXU0qVSr4ApAVPBh1SYPUtQ8+
vpTNStWizYMeFr7S3fj/l/BPn1mzq20zz7LtpKHkmvaJ6gCMMMKGDCROf5rfYLErmVrHItMdCnp0
Ttfq2NqyXu7gNEKjEE0GU55Q0PT2LVm0J/MKJZ2KZMgfb9L61G4pmUYc8Gxcfm6m0+7UcfW27d3Y
C1eI+LMT8t8F8yH6UeR6hnjtHTjEU7zh9ycstZ4c7WpO3O2D6WVUYG3x0ACCIpqxPD+wjOgxGsa5
+fCS2lBsnqC1+xlZR77t5FnD0mg3LGfxiFqc1EIN8rwixg8SQVRRR0QJ7ftRM3/mKQM0b87xTG2y
3XOrmx69ofmx12cyr3HtuJOCwzmYFm5oEDZHogVFBJ4rYpkI8goDGpT5wNwSMS60SxvZZIM4PcT9
p/yCXed3v9O9Sf7g5uYKFFy+f+w3D9rFP37zyMe7gJx2ULy3aygi5JBEBfMngEVBSA5YOJ9V/vYI
E+PcdL5EWeZ6Bx2I9v5CizMQphineIG++JLXEuGlNHeAgMfVElkUWVHCs+BsBmJ8a3xskL8E2A1z
H2YnvklJlm6RY4rtAotAr/BKYVMly8QXuo339Xsm8nHyY4Df7IFhccAPDdUPCdXkAj5lZRK3CEq6
fLUeC9YR5ygjLTn6bMIeH5CwfSMMRsDxS+T0NDOpmNSSi7HSILhlC6/EPIzAxWzFMoiaahRGtg8z
JDfqzEJWrBegFRGWLNxpNwCCWQns6Uk+9G1rmaPixVievlaGwMlQ5Fd6nhA2AEs9+u5RlL8j0l9s
OCauBToU5RLwrOOizgVluuiRHfjLAwUOszlyJx06tXdfMeXRyOg3oz0H40++p/ennOTg+fQbc3zi
QtKwt0J+YU/D8GqkWeybfqQ4tze8R/Q2WGhW/sjRYtHcVBSM3u2eHHeFn0atJzyBt+l5JNiPUMKM
cOSh4sN7vaGowYKGS0xxOeX4hmCQaIFwn0MEb4ncgF6FukUOuN/nm4Y8Zli6Icym8KnIN5DUzFSK
fDxglZZUW1yLUXT/YQtfCMY+Bk6QjwK2H+l+KSJ1UhtXbhrgXxqQAYX5W7MSHHcZbjkyO4MAC9Op
F61zx4i9Wfpukw0YjACE+iInOPwodxzN6PF10Ng8sc7HxU2kEPkw1eVaCwo9+QssaRepIpHonvVC
4wbWO0ZeYMw6PaJAw4orHSIon/5DBHsquVim82RkiE+ECVJnnBLePmHuU8z+lri3DHE6BaKFlgqy
OZZVYVCr8RwiCcT68Piig31H+hmS8PAg76rAMhf5GdfgE3v0NKoEWjXC4CpjmCGWYRLs1A8sylRl
oBhOazglUGj82epLYbz0y8mmLMLu/mkk4pCxNODY52nIVhYCioBRZNCnWznYhE7NjoNnawdcF0WC
ADBn4m423dYuJlJcYnMpvfOsY900DcGS5nAjArBnTjwk8KLLp9dd+QgRen5ERrvKrgMKINF4DPdB
fl4pLekg8r9JpjKKluIBXWMApUO7UnFwrhKN/vUnUCOBje06Z7/bxSyOzZ9hL/+7PpKodKVGa+qM
J4sD5zeOlEBKTAE8lU/7MFQZQZ5sd2a9E8jWEbgyDywKXWrxNc8ztmcc25PX89yCPYFxUMOqpRUr
o/CbPsLzmBijeMmsWX1rBCrbSNSXVvl7Ynq3BrPqllM5PzmI3Nta/9NUI3aQ2PUgUqzkee6nXeCq
Ob8LMtkfh4FjQ6GZvnWktFQWiX1BZffqQ1Kuh7NJHKNzsR4+coFBCvhjVMqBzimsOC2P/vaOCwUp
m8RgAIKNZAmj6KvKC6u7AxzPNtNhLb6q5bMXYB32Jnpt91jUUIESCOcVJ4XL/HrrZxmMlscROIuq
plvL3bPrY6DojaS1UUzxS5X9QfncoAVuzCXJfm/TJy8p9W0LI84P7yYI3vCUvLtXXvCcARQ90Fwd
7C7zhh7AZrVdR+bYXEhgY2qX3Do7bbwFBpe8GgjwXyL+40q0e/4XEdCii7orIuR2NGiiOfT4BBLs
YMt/mGi3d8Gy2sXbsF3VDEptXVA7DSSI6baubxeqtkVTZWpTQptj14JsRHCCBNcInSVHEhZurt+g
NGLhqod/CsnDM73gz6WrYp5K/84uDg58P8XDqDZ0RoIITOsm9r0Cy+f7TBKZ8VmTj8lCeKw6m7Az
fW/uApOYdsTePzKO9DX49R1CQOLhMMr2HDOpcNFCJhOXvifDRzlRrU4xlkeDe4lRmKqsibNI1Cnh
XSaATa821r2Sx4zreIuSJIHV/7t/axD4yl/i5oTgphzSNq8QQARjOCNxvwjvDHEPgSBiJ6Z+9ugx
zGHVxuQ5AZAIPcMBT6DQZCrC6BhXYU9u8d0JhXK/LdsPCXz6+iJJmc7E2BX2ZyFmaNpokcFnAAu1
zpEvfWKeD+urEO93168i/ig3azUf2dag/sj3tfbMm54uc63Bk9Dke0fJAYSeKJIWDh1HulJ4RFVb
Z3wvb4lwRdiWPTEAkH15498Tf3wMlv8suEezdDmc2Bn+qDvFDsrqs4uZxSkPFi3m1HEIHuuD3jPh
siLD7K667VWDXaPCHd9/hmEcTbIeqlINT2Kjn0cySzIKTLTaItZ+IzjOJnw9N7O2qMh9bjzZeIzj
YzC+cVgEVxRsr6POAtkcQRJvePUwT4HfJE8HOY8CIJ6eWZO/RqBkOlwJbP7aJPORwOIQFGSXR08d
NuRmxEa5YareToNyUyHgF8NXbTFe5n5WhFOxBU5HHVKqMVM4rFNhi2epaPNvoECl12e62pFzdYl6
YvSdUDJ4iXqNvwTEx9jLXNgnmhmeqDhAWhJHWxINv+3LNVmbC1QJ3YBbmb7CjFcCQP+mW/ZSEOIj
f5geCNmv1PmgoowmvZQ1HM6sCZnYg0sqf84XZI20tS2PxHwuU6/zkcAVZsGAxVlWwFZO2BNZoxXT
n+wHEdvSyaO6g57zWPbaJzqke1+393qblRTiuLJhA2RIm0vxkyKc4n70+jx7YPkXaoaVCiz7NQ8C
NHwszPdLgVRxqsM8TKe+VodTLTasD5fgJEacbSmIxI9dUQYRvGoB8K2VlBTZ67krDrI+JpQsjCrb
rXuLE+nB3I6OclDPd669+1jJksQt2tAIpWxLrqiJhvX2sMw+4PS/k+Ik6G6CRnmILBLc7+qBC0D6
i0rsM26HAS3h7NadCLsPsYplO1O/07O/tTj9v8wrDEZdFJlOxi1c4uDYvUjWIpYtLEflAcirQmPd
s7AnjudF+n0d00lg/X16oROlwP+J6I49aqcokKqITU3DhooDRIKeciDivoZlGMykuFuOBlBrdUEs
FRFEtlheCGfk0JAeHxx8IdjsLQY6jGlTxUZUwokgyhIMc1hDCKuXezh9yNq/AtKqu9UabXIgaX0X
IlpvW0ycjH6vSRqMbdT8gIsAy1xnlPpPzfwF3NHoqTEAwPJ/hLSgNpYJJusalnli8YW686qHQB/A
w8bGLgeBi86a4ApOBcBG/wIQ3+WMeFYn6HvKBwcVvtmNToSadSj26RqYzyqw2ZMF3jPvRwADYHLW
U+tlvO+ZH27CUYFf/+IuEGizBIGGPqf6l+wpZULpWCbiW3unx1tzsYuzAhaS9vxORcMzpLjuxwbB
wnbViNLMBSW0ev6vq2B2ACYh3gkvBsY8jPXIG+kRjqpcnSbyFh65yMcoB/lk/hlQ63XK71EGwSOE
cBVOoroQ2bM+33ZpglZf8XO5+WHW3DqrEx0D2k/n5Tc8ywT3A5LaikqDmWjrSlDXeGNMTN3jiiT3
l0FLOXvDQECx4MdqcKAXaJerQSgWVBen4rVvP3javHhNsEKnbl7Bb0J0gOGAE6vxeLHUt0x4MHR1
A1QHlDk7W3+tVawA02FQOXlxI4KqumDGkTMdVB5Pan1TsopBL+262Nm4BqUOhSyc5wpjadLvUwq3
Jt1gBghzN/mZY7Ux4uHtaKPBuyUqjjo1tgmTl/5kpRp+dxhVVn14C79gMvOn/xUWHyB688RuBzyq
xUhSnUjVjEVRDXHwy7XrZdvYdnVz+1KKZ0Ji59HiMt3ZB8b7/huYACYp6+4fqVDkslRwKS6hexhN
WkJc31u+Sv3ZJoT0hyo2KpnqNKEdT6wXGROhkAGZkMaFG1uAh47jzdl7GW51UGO9W4yhZ945mFWT
T7YlnQGQuaF5XhBdlWeiH7ITeGGSyjm1VkCwWzDxs+4FdiBfyUjGqjq8ZpeADmcVkjSzB8HqDhmP
3v0LERjqv1lBYfymkLf6so5IS0lAwUhsulZ2qIIahTmfDd8psKVi+dDwgsOei48FnO2dFLj8HZpm
8uct6cAqdL9Iaidta96d4GserC1VWHQ8suO49LNsCngHwQBV77rrosgx32kUWNmVqdjYGWbJ/B7A
WAbck0NBGZxfc8vubYsB/YWAjiLPSgGiM+7affIwPaam/8/FQA6goxxAD1aTh24BBOsZp9wqqSVq
Pc0FRZNXKba9jonAZJjEoYlaEHK3cUUELHP/es7FTLZFTvSPaQIrCHW5+eL5/BQFXo9XbJmR8+IQ
YWwgzhr+YXKSg3x1jYGrjOtPGIwXmM5RwLC7gRGiYhAOCos28z2UMvPavdOJ99ZHQK6WbvD4LlFj
f1bgRL/cCPpPespDbN30pOJzYuszfuJNP2BE9FK6GOTOP3pW+1nRWcUCR7LuyKGZlP3VTlXkVTWK
OJtKCS8UsrDOYf214HVRw5QkygHAbHt51PjgJ3x4zttg2/K8jQ2Yyh+MrAYAyGy9YZoqpTfpmH8d
uhar1JakSA0m8n+orSpMJ2YiTV5AyoRcH7p3eFuIR8i/w19+1C9D2ZmLb2LzB9OhZUrLyvJxj1iK
TRotNpjNLFg8cn6sqsB/AFnShFVjH/N7KKVjAtMr/96mdCFmCe1sJ0WNltM+zJX5xOrU8IfFnxT6
8ZRxugq8Eg9+HdQ7rQYI3bNvWwKPHoaB+0NJHavBTnlm1MM/lEpOCamaO4vTXpvgVLb5XdAUsQLZ
wHQXstQLNihrq8sqyf+zYDS/3lu6vZbr5ZZ8pmsvkNChgux40JKsEEPGd1mI1vkMNJxrHuceRuih
eV3yszJsCW62pUoOI4+X7I+gpafNxISwE2A3RQAP0Rd1hUqIpTkY4Rq+iH0TeRujx/al1POFbyXb
hhXFk3NOeIlfIutR6CfyLeO3YI6Aaxypha1zHD58NV6zU5ReUh2ezQJjY4CW09wsJKZt0ZjTg/Ea
+YGvRv5N0B7jiHY00BieWgif3Vmt45+dyUgQG5uq+wrPKK1fIWotrd47wsiuWSq7cGndHz7LBXHY
cxsHu0Bns38CS7+rInQXRGEtChTCNNK1fLa0N/oeJtw8OaK95B69tBVLqwpu9/3qlihPEuRLr2fE
i528Q9nernuPzXzfXPF+Bvlw2ugzM5Rqd4OPxrm8ToZp5AV6i9De5M0dXPGzLZJkoR8RyRLj0h03
8QSQbGW4vwrUQ4UwT2UsvcepdPQTZW7dnxMXWFd2iEjxvR4SoKQkeiuzLSyog8SqNCkvwRwvBGDk
keBR0sk75sbW4SKx5l3n0WfPdBFiwQC/hIjMe3UGasau//5kKrPQGQGAC8WZXTHdrpM31lIoiU09
YSOOhgDMTSCNIYrkYwPLDa13xvHsOrCYPFJ+dJSeXIdfWZNsdfnAiNn6EdSS3WZN26Ul2/ae3vQM
cOyMGxyggvpbTpjBgUi3cWFRqmb9IqtegVE2pxOE/ghZW8XGaQwqnkmzLHRhw/umzJutsGLhePMT
22oaJf+SzR+X1JR472B8L4P8xNIuzPiBA5u1AdYNlOYG1bhPxobls42vWzBojS//r1OwxqyG297H
KoFw8nWJZd6YIYXckscXYofS2k1O86jKNIl9EURf8+7zteGscN2KwCYpv5KBnURtDLCHIIm+ncB8
mowSWt9sW+25SbbfL33Lc06F8wAk9o0bkszxGb73p2A3N8t4/itdMnZ9HXrPP2+XALmzGMYYpUHY
CKbXpgYVbWqzUp3u4qq7+AQTzGHurystxUKOOS3nIVnqW0OfxnCxkaLF+cBvbhGP0pAoXLZwy1ME
/RRuu3IUAYPz6Q/whNVMIJd3hb9ZOdONjhVSAhpdTnz4Or6HE0CXXUdtM6QNPZvhhRxNaXclr9S1
DMVQDUmOg/UEy2vcXc9/xcJ35kHnyE50tm/d1ROSkbQi09UyNdNZyC9hDhJjYfmMFehMnpwCtzRH
bnuYbf5+jWrwTjb+0Mc9ZOzzT3VqP4eeorys8yv+5WkuaCQQWp555bx95FJvflaw0nldj5JkYAa4
EVQ7kQYvE7zIYJvFjiRf+TfYz3OG8DekHrxqWOL0LRXgxB7nbtloMM7Wx2rrtwBQyECtaisEVhxx
TmOY9KtmzdLKh6ois+TaKdCTVR0SWx0hgXJYx33/dsYuBZf3zr4EQBLxWReKQfwvFrOCJcrt51bx
GdaRNrZSpZKfJeVAIDPq4AZWHjwy84zHxnVpbT3+4q+zdOO9AChDa+eKQWevTU659zTEpSoPfJm9
7FH0M9A2bG07utzzmRQuCBrplH/BeGjRYDew0sNl8aNjbhR2aWMv16zNtdy5etlhvUc89Sg9cBWH
lOkVDMbRAgPN7igTUY1NjdiTfqbbyn4/JZoFz95/zmOhyfu36nOJypObs5Sj73SPGq6Z9CS5jAWm
bgn49sLleD+ftoJwzjerl8Jm3fSeER/wL+i0pZ56ZVLCgMGlcYqOA9VzIqwzz4RG9ZnDy4c1AKoN
AmgyE7iGrrSOnoeryNxHbcfrQmoTP82f4t9NNhdOhaQUfw2bXzZySuWN3b3/DJTgnz0838JTIma1
dfM1YJ+QKQuYNbm50tIb+PuWCM8aMwTibncMnlhxlrTnyD9bqyqAupmoqU+w4+xntQI2rG5hqRZV
R5TpkTlkH0J0qrUdj6K/L1rHSYyb11zYx6Us+cfnIQ98M8jVi4ASxkxNHs+2ng8xShMjAO7z4oxE
6nTlkx/mN8eJ+Wr5PZ8emwM1vW3vx5+tPL6Wm/Z29D/NGMsIxV9ygQlq7Bf67KkXxKcpiaFnZmYx
k/FAfeVEtoZSwqyHc9J4O1EAdwi8kw5gPdeqBnqbsQsBSGxWF++LUziLBFKBnXm4KW8mR+UGDIGD
YsLnBKdyAQYAVfSUGgM1pIJvkDND+GN0uC8DWIRP4B+zm1YG4+eJefO7njzbGCDcp6MOqCYwNB99
jMATq/HCwh42DEFCBTvCXOZkqtkX+KjZmC46mH6rGoInwhMNtAYecx+gkhFSZ494mww/AhhBi3se
25j+knXgBLSAOv6R/sy7ii7iTEinF0fR6zqCGYlfGsI7hOolMve3MKneGBKhYrCsUDEaW6SUHP/J
CY03xSifQqH5yP79Tugnk2NJthrLjUOyFq3Ql2susGjDEdlu1yGe+1pM3KTMMcqkUvGvToPlGmb+
U4SjioJRWE5kb2ZOLyr9rfBcxY0tf7ZHQJnvBshvwa8qFVwH8zOw/jiv27AMZXdGuvphke1QNuHh
Ib9mckZSfPlxwH7glaYtatbnsTSUCEwhWk2PmMfyXaPEAu4aiPK0+t93uVHKIFygoDAXBqda3AWb
4Lwnj5zqP1d3Ll431CRgIaCY+sa640AnK04/j399/gc/RaaEDRn20Qm3d8qDuVLtC7FX3s8RkpeH
qEFFr7QVLGoii9GeDSbk/fhMJha82TqzCXSVi9l0CZZWXYS99DHj262xdcfPzaV+WBFH+5uQcASw
BF1mGO0AF+trsXbxYbMFMQb+bqc7gdOh+k36EP7CzpxvfL4hqmVX4bbHTu0sLY8ifL/9hVMoFMwX
pvhvNeULbo8Uh0djQa56Ze9SkbjgswmCBwq6gIaywZ9/InX+M49IE9lvDg/xWifB5rjVKVNDaVjr
Z8N8qXhQD0tyq+PnjlvVfe7Mr05aQG7wKrUhhu3QxV5ZhMo6zzbLTfd1GjEVEss8L87KIO8YhprT
7Ebd5OAGmxzd3mNxzBs0VibWzdChp1gv2Dg0JxVUCpz5nbdjA7ylLlJN0JdlK5fdDEWT413sPAr1
evSDZkceDABfBpqvNE9iIo/QLBihuUWSnoDsxBNE1Mb1Z2lG13mcILER+CdQJ/jNfxgVvrcbh38C
02tSN9de3eBmaPJ5rBUXZKk/svnE7Q+sFaYCeKYi/rqz/p58LZWexm2IQ4J6GDEfMeXlKtlUz5mv
aJJx3FABSDRB2WG/hLz+y3QX5eoKzh72NO2D/VlmIEfmhH0HaBRvY534D5v63BvCgyxGAazI52fc
gmZiqP/IhE+HhJAJ+7nja/vvNIMLu+5CjGEmuerxZUtjlZPrPKiAOdW9yineRqzVuFjjq2exQoZb
hAvSr5s2try7Shw41KcwnVSYY2O7WIVfmUHHj+2VcUN7v/i4yjEX1n72gFNvfycDl7W2Ockt8LBj
WOjGwoXyVgeO38DnGidUCnHJEQr+Ifh06fs+ZfkRRsGnYRD1jru8ZxmdJGR1rHREHqgSJEhlTVkN
pLJCrfguwprEx9IQEO0lDtZseYpzuGwJ16TfpwMm4VbnMfjfNMu9nEpt0L9d5yqQHXX7+Smkxc0w
ZJmQgTT2Mm4yMBf3vNF5tDWwC+Cdf5P7F7S5BpgFQGuGePTNaJoJT5QNGz4BeN8lvWh/YDIMXsWO
GvJr2EWBnYViIIIdwlBe0tBkpuw7R2lvlxZDzeo2lYKrIbRWhAWeZstlNIi3y/L5eKIAD0Ccrxgg
t/a6QeScbVavJv9EVsrA6WA2c8EMPpN9MDcIrtIc3RmoyT0X+pGY6qQqxH2dt/j4WBaCbdy0rfFy
pH6gtezrrI77ByUswWYD2+vyfaoDGVF9ua2JqEU2wi6DQRgOxUeEDcp6x9azrnaK1G5Cb4VsuYft
f9n3WmMLuMa2xmsDvPTl6JgVQ8woJ3+bd51sQp0LuzZop7s579dpn4HsDtN4axSjoSYDzMIhSdbX
LVsQjWyNbIB5S43i0DD/Fbp4kbSutml7Ziylmc7oDr9pJB/O3928CrhZFaqN8X8fiA8mB2iBMcuM
qE2N9O6OzuwT1krmfPsagcOW09Ue1Fn+E9VLZJ+V2QDoTR94jIh6gp3DEgIfK9CaX8l5KDlaoumC
kAMDl97OgB8NzkICJrNGl+2YM+1qTJSyUkwqFDGo5JYHIejvVJnW4vHA2GB5C7E0XEjiQb5L96Wm
IGWwgqYZKcFXYSqAd/xfWy7mu6Qn5X9FhBETwIpuOXIM1rzxeKet4VBZaCapsocb4fCq6t2w7sBC
9vL7roYRy4TRgEX/y2z50zsFSpHlNYeC2crqFnwrM81zydAna5wSiUGOAO5oOkuhfNOWgpWZ4gre
iWOLtmx2jJVax22dbvFy6g4ZJY0z/YfGi5pkgr9hjScN23rbFDvIwwm8NOuVU7eXOTqKkLN631u/
AR98Os+0cW1DV4fv0BUnsiealRRjsrjbuo1pu+HYQj3DsZ6pQ/hUQl8wH5cMbLNWa1smJH5KNx9a
BMrAuy9+Px5v5mO7iJTF9k4qKNzcL45kFCchHSJx4bntQwFnx24nICuwIvmAkmmeyElw+IgrjGNw
4zW4C58bscknPdC50BkbK28D0ufKeZ9l0KGsbiFnYpgn1E+c8u9LZ17nU9sFiAbDlCxls09EMEf/
hTEhbEFJ+5hknhLugwjI8M+2thbIysiOqyoIq08O1y5kiPSTNV/kMrIdQiL/IbJvIHvhCoV0dO3P
+/V6Y251wg8qciTTKGFa3qTHvaEvfZ6TSMN0GmFGcdpy8h+OP6MH3d+djS0nnROWvJUM+3CT5Teg
WyUXJSfA1m5QS8plQTCri074ibPDh+Rr8isqupfsB1WeNRpGPpZpQ+W3lPZUYdGSHZEZYqju4END
/eBYNi6+giMEfwSiaRiUTVHsEICpQlqngGhWybjU0JoexUwcBv4IChNO0u/i30GB+plz4Ah5ZkSz
B0dAtJkWmMNWLpMMoNa5oi65TWfu0kGdviWWSz2Oyr/ikZ0nwyobKHzXHHdcauSunvPuLhBcSF7O
g54t+PmtZHNqiAkIzTqSd4FennsBu3jaIvb+DeJSwyOp5z/qHSQEUVa/+s5VL9GgS3VAj8Dr7tie
29RHl5T87dp34sGWyNmcrrqeZPKGLSqd2DqzKS2VP+icMtDmDki+J35PxOpgSUGtFwtTHXENjdt7
bZK9+Wcmgl2dssgX2N2OQkyQiXZzSPJJNFX0EqUJNmGDuIpktHyUzIdrm6XrXXfWXT1Q7oledaAz
mPOmfc/Nn9jbaszzWFE9Z+cUbZF3o56DqBTP/m3x/7g7TKBOV2K9BwdE7hVamoGfzNnuKQuMulom
YfOvJX3qzZCJtR9c5ML+hUxjug0RozrUEcVdcAYLtJGvL3ljTfeSIf8AIcs6G3Ee8DZPPSDdhQ3O
xPSa5PoBRERAHRrJUO9AQR2dDfdSHIoOZCLCeHMPe8+C72kzeUBZp+5QWYiVsn1VX+/VTLEOhqzC
LXbAGdUDxwYttXenXiqKENiGoKsWORE2QSFCkO+VKVusEGUPb2Tgdy3mG2DyQYN/dGfWyEIXRBVg
OdqWtTL0xv/CI6rl5AxzSKkZ7ccmFofnWWin/nQ1aVjo9gz8UExSJavgIOnXwYJOLV2LA44iTrqT
Zzk3AP7nj54wxB+5izvwVArBcaRIbG8G5B4ECZBgiZ+/zuKZGy9RrqpBpS3LFCvhGnqWngevf0aO
NeMWsnca05y4iPFbSA8sijFwUpg3FszFlR6dC0848qRfhThmMJhqFZUEBMGWNj4RrJxresEA9CWS
h6FOJfiEIWNWjfMri/cWBU2uP9UKPS/ML8ci/cLhc9v2K//NzQwjRn1AmzhYFmkxcbn4fSDVVrup
bb65E/XGrJIbvSyn24kKW+367rr+GGLFiapyhoV69jtIT8OLSVeILVkqr8Oz8J71xjxNIr81voK+
wKetk0YoRpriKWKJcWzWt8sxQqLxJXfwt7uArPJMEwxszxhD3A+XVHIgMKNqpSZPwiQ2W9QeR7n6
UE/EJrfYAG7oOcckxX5YGXTl5+5ralsppQktSToUj87MLXiy9hTPRgdDTW5So/fa7q/T66m/7uhw
RAey3BqImxKysk89locEeBP8MCo+FX8IcVVxlLHjkE4B1Sloo1XbRpD4fKT152r5cDg+vevWq/rv
vIwqzwl9ciVu+wJa74rEJIB8ILRf43siyADt8zKC3mE/33FA+mWkcOBrY/bh60BDN49+c9f7xi/y
S5KJOk4ni/2X7AcxaGrdzztvrk3ngW0OkAX+GVowgzCWyuDCkYqL7UTNbetn+9kf+sUYhQffPtpV
UsF+cvccLYGZticLt7o2rQIsf3SrerYr0Y3krsixT+rbXiV9v95uaoM5fvp/50G1A8ahCCG+I6lL
CqOQCr2UwQdCMgU0PiOmYeQsc1dUTKkeRiUF/prCw0ud5sxljex8Pnn/W43Te1pBPc4XHrIL+itd
gNdFuQVELnuUUz2H/F9ngdCr0Yq2xbpAaodHU7KtzphGPU+xN1zNS2cJzjL4h86ZZlTD7NQPk4TK
gyAYz0EdLBLxN4DKoUWwQ508FHV5zqFJ5raLN5XHSvicSpe5l75fNyYZwxgsROkoibLy1bUYKezP
tPWZsOwZAUdgy835/jk/LK27JyJdPzguA7ApsYgnOSm9wIUDe58dMd2MWAdu0wt3G5Ltm7Hfu/tu
IM9vBhrn5ZFCJHUiXFHy/+QJB+uQdS9koJ19ko9IyvjndylSFnvWcV13aRSE3HdxzHRLecL53n9s
KkK1OG409lxrF0Rkgz5eR37mKxA9f72xpv+yVrQN8Ax3W74aK0MiQE3Vl/m3q74dD+be4wFkqVnY
118IW1l3NjhU00a9SN+1HI2vV3xNDyB8i9yoMBzUTor0fk+MFc+MIbN2vzPTFbdBJpsIrEcXGUUK
vL/KhRT7O2HAoeQjSbZqzTiP4Oz6B80ntuLUGY8vXYguGbs/Ha9SgmOkOPuosi+RnvX3JjuNPU5D
uc4PC7j+6TqPllLJZe/sHUp3/m+GSNsUBAksZ33m1HjModLqG+ZDpQW9nsxWCpH8f2iNZwdcTq7j
ysUQm9qzI2Y87Dwz2barYWTd0JA4Av1+SAARmRKajOv2WHvI6/IKtsPdZXLboZOqFODuFbSXFZxL
2yfrisu5SDteOVNn5e0n60CnnExdRQHoTyD1pO8ZlliLRg/bqxCb2Y1IjvtVyLpFm2lM0e8ycT00
qo5X/kiFCUF104eW0xLsQvrT6tm5ymARqRDIlmPqKn3caTzRGVL09LMAPPLhWw0DK0281Iu0SRbj
9M/M4ht0VJlBSQuNQxsy3s12+u2puFKbn2ktzjf8KNydWqIkX+iuNB1qaI4DbvwuExFIBQ0BpjHi
Ecz3cee6/oKolPBiwxtre+0DZAmf8NA0BW4FoucJxyVNREhzkQ3WlQ8X1aDsy7kCcGCjQ24ewVYH
iock9/0k5BBsWPDTDt4Mjbk6fD4zksZ+3qmpMT4PWUn9myn3euC1Q3YXBC70Bqe8kfukxQbGDdDm
YRytrcoiPcuwzizxAUnnk5Atg9KBtCDA4sEmTKhyhBj6Ir3yT99/KNj8oPO45E/czYkUGZNJnHtm
IpuN0q0QnuxAn7Q8okD/42MjKW6YFyyAFp4nKJQ0uTmCT0mrEowsRE2uRt9Sb6bTTmC6okz7WbNf
D2iQF9q6osTkf5Ju1cilI28u9MAJTUFpAsqn/rCavwPbS0Sr68nnpQCp93eI7IqeL/trjffzxNm+
P9C31ByHyZZZI2FxpXwLj8pfUva5OtEg5/OIfx5AwcjlEF8lZfej983vl60jN3LaDZ2+cf6qqM2t
OpGzRbBK8EfCfSFYM/ap3aF2yerA6FiRz+mmggl/FtSko6Ue9xcJUfpBe9ArG7Eafg5cMF041l2z
t9sgNdDaQAOeLVGiQW5YKKmgopttiGdupc+s75rhOXFMqyNKOzGHrW6at6sJDmw8u00PZ1MfQhaL
BUAuGsaa1YSrE8NpA8U+ikNbfW5IUpuwA9FjNEXmhiAudwi2yHil9uM+eDoZqSlY+mq0uvomXO76
XrjNb7wn3/ggDPwAz0e2ZCnodei10UlcIBUUvM7x6NUfhWzt8q7w1maNFgkwVFoaC3x0fQIB7Xep
uEdAPmsFxJ+Mrz7gxCiQqm/CWFhTBolHOgbbdiBL4lZgOqlVhiQQgTGikXoRp1FQftJxiLXjH53j
2+qlwI/3QF0oWza1A/Plm6tIlQgFVcNt239crobbzHZAIIiKJV//n82WQUyUTyVkN9kUS8dMsC+D
/fQ1dQ7j5mIi2x9X+LQaEvyBeZm+mHSsJmqO5/AfSsqlmOeigCY0ED+Y1iEUqf60VkoUbVhOHBQR
5WkjmF/k7n4VLIZMBNUtWXWf6RESNC+F7vHQF56TJQmgnhzpAhOzzejqkN1DFis2hq6e3aLiyKTa
yRDkG8CpsEP76wqHQ1s4k4ONvTYOeJGfDE6Vry0klW6GNgFtRdBBb0i9PQAckwvLs83oBKOkM6SK
K9nM4b5SiuUFJUlhNi6dEVyLq8g1U+EG1xQd4OkPzxdYKPp4/R3cg2D21QqkT9WcYMutK9F0tXXf
ofyRfxzOq76VupdxHqf+/qdzAUyKasQdGTRuLnHHAHZO5c2PeW+RKZd4XVJbcfmwMShyOIHKvr/Y
6N3hU/X9dwT4p+4RP3U/ZNxqNcW1tGiTjmf6c0FA9l6s/o1Ss5iD1o64DczWTJAAK+/ocSPOAoVV
r/7LYKVZYEQEsHKH4q5Moa0zbzyrRkquyc71gZAvv0n0/Lu3OpuxxN8IDujXMfHWCrAIm7BGXERA
SeYpcRgygDKoE9VljdsBcpnjYyLyGC6yuBpcQU/fizzv0cwq91M2mvl+c68Mch+EuOyDkrnkcbxF
8IsoYcnTSJIsWvBr5TF31RJEJydyP7gqrWC3a73xD0HpjcHSfTdPxtdexcUfCHEAcug2fxIjJXs2
DyeKNvj5LzngeZZSMgQMLMetqLQZ6+g9szitucWITFwEdZVckEPTAWYoAYpBEbV664fCWVTymQGF
A2+RyYLcaNFFVwxLfOdq8IDi57oiRpWDSuWJjhbvx/H6SNFay61oA9yuG+BnNo8lbJZm2HzEUqRJ
0efaCc6+xDEVjv2mreacCZaS1pYkr+CvCSzGhiR6QCRaD15Qf0DPHcvEnKcRamyXXLc7w+zbI+lJ
0dAVJfDEUYCb2/rDBYzmHzyiGJnemhxMuTO7FyUKuSzdDN5KQPYUp3n9cYSTvnx7072BzDcjHChc
kvOp2GhJNvCkdPXPQSP0UF9mxIbcAZB+c+XaDVgDGOgHo8bJ4cn5c2QiM0ufCjn7oS54YaNMXQDD
zz7x4ZKfLf4tGi524/TdSWD6A0uOHvBSeFBTbzIFtYxBGpec92QKqdbHSiNZJIRx2TK+SpRf7x1+
hhPOcie0KYdPNX4mOeZdfY/MOS3GFHJNcaUix+tJ1ufWAAhbanTfYEwtmCCWqwcqFOZBcwwPdxcg
XYy8Mb/TvEwA/AyDHz/gyyn0qhLniZrr+UPZWU/zQVuxaF7MDiILr87FWtMsREt84vaHEuRGO6Ug
eqrOLPT686gFviBhDs124JIpc9wfwzGd6uUfBjmbYG01w9mFsnMvlbWnpwMjk3Cfhrx6Lb/+Hc0R
bSZNkaZJlgmIplZMhtBUaFbG5FU8D6aTPiqniTzkVE/5ID0+8yV8l3RB3SzaiXwT3dkJn+5maiMI
qkb6hVFWpT9KgFl/Js60qXwDS1OMD1M0kQLekVcGiQ+o6FIauMX9XeMaR68IXJfEIQ86G2TCbKKF
/e2BlpEgJAxuvt5dwCsjNGbeoedpvtChiSwlINynyWFlx+KLSrpYt93i3yR6kGc2sSErfyTZ5E3C
7QTF6EcN/g0AXI9eNOCSRbwM3vQuhfsao/llRRqIwXYQVOPtUIdouDTnMoWw8BOUH4S9Pi2fz2u9
qBzK55n7VssGB2TiTZAtlDxoHjjpw6JQE6Q7p8vyqvQPCFHiFnjfPFIA27rfm90TR65BGm22BMM/
NuGS+eeoPEfocyDXvjxVIX1hJP+tm9fMDu7Km6R6KzlBAudX1Rz9KShj9UtzEvE9QXA1BM+EV05A
SAmcQ4u28OS7RSvlw7B+QC95b2Lekb9jukRCLOfhVqoirZB23X1rqL/jlCDV5pYhgEKklN8zYyD2
ATLdu2OQtNUim7WQxlewMzFEI6msBUgDKh4apwfBXs5+JBe7JrIzJNVuLjrppaXguJQ/V5PrASpW
JJxdhF1R6qUy49IK/kfEADLY6JE/3toMo6Z/15jQr5QMdvqXeRfku7z7Ibxi+3GaTz+s2KQC4eGM
jR7s9avanYEk4IQNcYEQAqIjLTjuSdDCTPYP81MncxKIvBAjKQ7ruk7Ry7ZtxoBGvw/xkzvXFbty
npvHvnjfrTkn2ypMRxUxwd/QtjodToRT76LPqJw4qj6msUrnZSoafpUwt4yr0YOkfNQkQ3gBwegs
Yct3z1s9tE5+0Sp7lE6xjeVi8w7+CxSF5/y1HuEbjPidcyjA0yIDhbl4LAXDr+6lokYg1MzPPsXd
QOfeWO5V2JHEWcWXOghcop8oVuiACFkNqBkjkrAhipllf3C6ZZDVcOB7Fbe06blzn7ypxKfvlPKh
N6xDm/TdxFI0YxOCJEXMsntz9qSbSSMYmloOpfJHVDilHebHyNrg/plEtg8/UxdE1P+R5W/9JnKE
Xe2QnrKvgzpP6Vbf0T6fk8T5fNPj7OCxbmXkR7u3R/s54/6vOwnhs/2ATiUwbR//HsHv9/aajCtk
ENUH0xbEBBhUd3rMuUxZ9eNTOYfQJt5wyetFjWZ7HdY2aD+l5IJlevIQtYFl0UeE3bw586qcs9hs
ecb3jxmSz0ulLPvLINtiv8InDiOUk+xdAFNb7p+UBRTXetCpg5IYjesEWilBk24fPThHOTejr82j
xlepMoCEvYibVQRUKKyERkI7AzOUsC5OaKhTFtcNuvBGKzhJge1I8G9Cavfz8oCOK7d7E+JYYsMw
hUL91hC8ufez7Tc5kt3ctH0pCE42MaMAo3UaOJGb5lR+zYMi/Rg83UHCFZv2shk0LxgqJ7ebvAC9
6dNAVuoHwkPClV2GHn5O+8oIN+GNdMnYD2YxTAqYIev/wPp/7tsiMqptTD1ghWykgcRbc6bXjz8A
t3/xatAa87+3r6HAMHH9voOoQuFjoCaq+sbRVSQ5jiyOyZZWq2LW1o0yvBDXXaXQywJRw+Am6WsZ
/WMw3QCzDkdsf/oFtp3NwG1X1OOLPNt3J07lqhHCwsQrRIjYKyvJxLa0hQVqK7gR5nX+isAT0FIH
evnL1MYo++qsE4WCIkj2JTOCPvMHL5YH6LGE9WDbvayidu2XABk43iaDf/yRimZLhN8ekBxpqjRY
JYeaQoVvgveUnRiuWRQ15tm3ZNIqUCO1WTto/Ozmk1TcTX2n2uIhcPaxZnztURqbrxiyOQ6Ee9aX
NFi8uKAuENhAXqDJtPBtMCf0LaXq10/JV+XS0GeEAiDixExvUbdnSj3hHd93KawP7Bn8BW2Djy7m
AuppiEnxefC/6Ku8NcbuVf2iJMmMSKyG975w704MTduXYggklk8WrbYm/U9sp7mvmGNsPjCM1EmM
EhYn+zVabadsg5mWY3m9PEeNOt8A2x1lvbLxagtXAxmbSHamDNnfWW4q62QAzccWzgHRKtZ1slTr
3p1UnDH1R239HHJPCr8ZfeCvaAHn83Hcxx/GdoKFaps3gELX/0rXC/rnjf1FVOOpaKMUfxjFUlZl
Niq+wSGLipKHClGIeyBxZmmk+pwbIL5hfIYbURIzJhjMwhy3r/9f1I5R9SG4ndyfF9/PFLEcOZ3H
lMCg8VdoRc4iPsXaGmU9X+OogrrLNdN+G8fp5pTrED1hh3K37XuOld1xcKt9F8rxbXQKzirN0Xvu
IZUYF05EMBLyFZnPqhHCfsNmfiMBjtFUjvwaTObedabn/X66y6toB7PloE5IRL9g5H0BI0jqS5fx
12K0WMOhEO0FUfW01wW/dSr7Nl5ZmXOTVToJGnGu5BmXLH16BwNuRyAnvbeK1NTEqttUAOMPwh7M
ysC6oBZqIZr3Q2uIqI76qHMI5NIxECtyRDUMgN/Nmqpj9xK5syEvMh//uR2W83BGeBImCMIHqsBf
zj2F7ybXRrOPiEhWFMW1VXjsj/+ptg7LTYIiempV91auygyMp0v/R3ErScUonH9UcIJhUnbFsUiT
A9h7YdVQhtKJdetqDXWuAB0Dzvcj6hCahGfX7W0luv/FvXm34SwJLZDQaEgk8pmr3vnIA1h6rWxL
j73ZSnw/JWR7et5Spf5TvsIyXGsiIWYlkK7K0cqf8fKQjdoTb5i/xk0b5vSCVPEho+aQyKk7i0Eq
6hBSE0oPEO3a9CWzDqsjC2gQLNKwy/cwC0WqHzXOdiiTTVqZmiR94mRVmhFNTh+ofTh8dRVwGm+H
Be+ZBNnml3NQSYdqN7NNWdbpCyxQWwMHv6NgDNVIKCZseYDycRPgLSGsZ2bMEdDUdLr8S0kMeDE8
+++xO9SSZSISwr+0vk47fDT2BCVurDbQWi8Eu4vw7CLQcVA+o2hyDN881CnU6nTrGSZDVtZQQZVD
lxW+Y6ppqWjJcUCX6tae+kDofdjRzAEiEBz8e2/GGfsl7nZ+e2QVngZaT5JLp3uFqXqC7+KJVCKP
1BzGu//6tne+95pgEpO5r7aMTeANTYUyXN8Fa1AirsxFwlQ4qVX++6LhWkJJc/sjmn34/oOI42pE
bp80WSXoy04wUFnN3Vwn4LjI0liqsc+tiBJ6Y/AvS1yswweYMKIZHPXiHbXZpYRbWX4t0qLiV+V9
L574HD8i91IF2qAJQog7qa3/hFZ6rdWowkU7CNAMBd1qod40jedgsAuT0g5avejAm+NoWLudSHiX
k6vcrp7tU5ELVmiWnXzkaoHHzAEXjsNxqRyPlNhuWv27rWGncQAN9JP+UxCn1eGLMYjab2HkicDo
HS7WlusmvV/mkt1pLw+gkl6ZALxAM4WifywTF/Hp+q4sJ11+d9w7b+LhqxW/j3Z8GWYkkLJ9Uq+N
Fgh/vDGRjMOjCltDxQ77rYVLW7hon0ph/DJgULTCMCJYs+103z//86BKItkDg0oRytyGlOD8dGU6
RFf9fBOGRNe7/ApbLpgbYXxqvgDr8sbP6RUQAwTWjCrOyUS11CtniHk40kT5RZrNX4OE/7sFtR7l
JFhrdoq/+RO4vTFl1v5eZPI8dCqXh+Hp3cCbux4/8GUlljqCRhRDkB4PhvL2dzlOa0vcjmXVVNnR
DmvV5jfAFIyheO6jE2CG7EJ6gdd8jCBi7HY7ccNXm++YaRaE8k3Jk2WFusHE/FiTTWSHOi6nH7xD
RPchclFITWofP4+z+Ag8kIUW2yjpIxmUON34BDi9NQHhfhWrn0CaYxjaw9h8Lvc3c07Qjkl9aCui
M+Jfm0Q1Poj3kn+o1ARPVnIE3R/YjzVW35m4JBqRdgpOZAe94Fyi4HHuTxBVXgb7tD4xylIQM7NT
vVToKSpU2F5rA8VewLlaMwADW8eHxjhZRGymKEmSBPZcfjPWyAE3RHWILF4SwuTDPcNRqpIMBwhE
xWFGoY3Q0OsGuTjOe+NJYemh/1MKJMN/vMZ378f5rhcdFCXsFy2TiZ4BEXxJpwEkS4YCm+6WT/Fs
rtMBFLMDbzzM0vfz+I4TN63gqA+ScnDJkEIjtNTHa/PdmnuhMHScmYVeDZD3+aNFAqDtU/BNiRpL
MCE7ZWxWXIPNHdcKnanOE03oAsN1KKuqkWUHe0hgbWOQ/ADkPeO6uliKuSddOrX0MZD0guXJpJEW
OhErNB0db/yCkdxKCo1Q1/6S7vO+O2onhSJqZrdz3laf7OBWyfyghVDM+JlzJGiIU7e2JFE1ygJB
o5IQbCDgGuSsaexfcNzLe/UvMi+TuRXxQ7j9ydPINHxQ/04ylG7yHNdxRgxrPYfAV5srqIUzpRLo
0Wdt3Q7xhwqZ3G0zRfQxVXsEPjdS1oWNKXz2q0WKS2usZpDPZOuIMP5bY1pwiFXHuypucs6q5TiM
6fV5Y4RS3YK7gY0k4ynNnlrhfcV49vuijq5Rp/RpgXcIWroceSFnfAoWYa48JoMhM60KyTpXOKDC
5fG/hE1udBMONassTGbzu5TIYyDL1GCm4jCeMmLlHHkZmINXiAEQgU0TclSDmjKHIY5FcwsR+pOv
gqHSR4+hPcLHlPdfVMJ46NTmRm3qw5EH28tTFjsGoKvd0kIPcTPj4P2o7g4+CEixE6KMmepri48s
m4QwBO2Ah5fAhMC2gqJs1APk8NkcacsgWK1u+uOEzUeMPEP/TvMFAoNbs/CHkdM94SPGEQU2Pi1S
p2fgW6ZPdcWS6dAJKc0M+5vvQjUhYxkvSKU41+0oX66XpTklKTjgPv1TMcq1DnSz+We2QPXb2CTD
wpTp29SdEMvhIvo7jZOLrZYBGEbvjBdwbpEk0zTKBx607lj7I8jD1uS7mu7ZGwRoBLmONPafLwWd
jWnT4kNsEDkXUbqfyW8waPXMQRofUsu6ZE+GmRORZT6PoP7o7WydnukR1uuqcM6xXA1od+3z2uHg
ime7FJr2i90DT182HKTaAd0YcWkY/UVSt5p/I9MA0zQm7Km9HWFFkkfUWK8T8YsfGwHqvksH/PVr
63ep+Ki/J+pJRh2mAIlGln+IECddyD2rWqp4s7mf7gW4Tai+Gz+GSjyvrYSKf4eKD6bFUwJ+pHQk
Z9IMoDTH78rtqqEovwejLrT4XWMoGv2WgQ2B+D6shrgJvGVQw4qr5QGbcpNc4MpUhSNm78Upjbgm
9gP9sFeQck0YjvfXZBuXd/1Ex/FA1RvgxEg917ehHW3GKD8hBZQtd4/pjLKAnads8YFT6v6R8HjV
uqBTnJQAf6WzXUEk2q3YsPdQBLVmyccXlNBvfMUbW+TtvwQEMsarHfjn7/BTz2RwewfLT2zxfXRs
CvJ+IU8+KyFXorh85Kn+1DqvyT0uB5VEqh3m4H0nOcA/A2I6iToJNew4TVGvJ0Ohm5GJyNAe/DHz
lM+Ype5k9UE0ZzQ62ZhPK8hPZmS7TzSHU6Ir+bJa+Rc0Qw/Ni/uDvRuZmh7m47LtVfrJmbL6dKwP
539TlkmclSZ+LjMLKzKbTdSmi9bvzmo4mVTrVBB8clnMx24zPzhrl+RE9yqMJn2CeqqP7g/iRZbF
prUKm/yR5ZopSTHHLj9O+LdcPbm7Rt6nm8Y17XcVytjXb5lybUln5d/Bycwx2nXjfJhJLm1ZF5MM
9zlKsm1eL1NWx1dRTr+baiJSdRIwJr++zmk7hoPlqAImb+vL7keXeby9Ic8KLTY+TwuwLsVdyr3k
QpridxFhSMgx0kXcqwO9rIw/IU5NhsD2xOBZ/RavpNHZ6DYptyXq6aE4xON8NMMrDjFqAB1bbIiU
g72OK8a9UIxSZwlUnkkA3e9MBOCEIhyUxKDOBzDFM+8hDHneQlhTDZUMzIozEA/znlX0Wl4HujKq
J9aeFHt7uPDSSl5I6TKTOu48poRqPyHDB0BXrRCPNz9/SEFu9hHFkcVQtCw0FJ4LsuY7B3r0JO8q
HZAQf0S1YvwV4rKkn1ESC8a+x63SQvcSLybTBCwhctCH9/r9Ww0KTPaxbOwaSKnG/vr18tj9Csw8
H/jeJT8x8e19jVCsBRpkRJbHhF+L7jFsAoepRTcbC30Mx/5xSeEUIyj3uiC3jhMbIkDCXJw2S3Nu
TWEOM1+B8tEIem9xlbNf//3Q8bCNq3yd81HTLYk3rk7YiXIkmqC5e9c+va8A1DFnmckkp/ikLlOe
WohWKtwFBMJYmNov4G6S2cFVIZj3n8CG5qGpZu7ww+WDzhCHhqd/hHNx364THdnfA9S6V/MsLi12
0M7xs3BAcvn+2IpaBjn1idyx4lkcBgXrLaxCaiqjaCB7nAbUcIEwEFOGaAUU/bGvHy/bRsBU6Y6V
BLATsFR6k0uTD1V9WVrTOb1b8EIGJiljtxJ/9wcWGTdykqswu3QQQuzdQiAqsElYMM4oob7O8vYb
4azHtzcQrKrpH3MutzoKh9rflGpS6C8KRuAZBH2wRQo/HTGEtinQLD+QWYSIubIq7+gfxESg1ewU
N4eAChKH0vLgvjYEd0DvkVXJUxqbXgfnkGGnC7N8PatJ0nLLlXMb/mPCQ0BkU9VJU03zvs2th8JA
83xbgdLy+XdK3/bDtptwoRlQRYLD3f0a+pn5osP8jJ6ku4SFeb7oCAmciGiH6xGwn9QYEKZeMGIo
cPB1QGivHxfiZsJxyKFdWlGPRTX18G8gh/03WdOAkZ/MsEXEsmFJS5aVMf6wFVjaQRDDOBz0B/4r
piCzweayci891L4f6QIvlVTWWM28WSlzYKZNTR7/wN+SNqKt0kjYxZ7qMMDVQ3fOxgOy52gjxMei
24xuEu7AjFIeyugTETobiuveiiyBw4qjoBUShqZ1SW3RV8HbnpsyInbYkMH0V7EbiBShUo2Ns252
EOawDtooZhQwi3jpsMJE7w+ofSwdU4c5NXHKiVFFi+xfy5d2u99KgcLZbcPClgl8EARFeGcxpCxQ
3yCnBWP6sI/IHUb7UZ83htIwqffG9q2ivRz3pZCZJmWt0eu6bPUGbHA8Y6CsBUKXYdmilnhx2Mgj
5pAr6LxQWVLvUMmc8iC8ou8vxlLa+XpfPdNN8ZysHGoaIoX2w5aZmA6TquDshqD6pgRZnUVJfhEP
Rh9WjUk8UVxeYdf/d/SuECNKmsGcaJHDt6+4H+qTMx/QqjqQziJOFw1d/9/0u8VYkKznz2Wju6qn
BpTte3lrHC6/wDc6azHeL8hZUcn3nisuBvdNOf6CvLuTRzTROYQ2q5K0+zAluQhb6B0cXOHaB5m2
hgnQiAYuawzpjEeFe40NQ9WV+RcUzt8CwiQmo6wjqL4vCB3KQfUxXPCU+/BZLpTn2aEL6vWrPHKo
Ts/Cj4g7zvG3TVle9LuImgGpJ4taagoYUw+baQSDc12OxCHqATDdTAHhv0IOKVpClk0UVGxn93kH
YGtrAOqRTOIPCSnrfjMpIl5iN247+i/VMKhmpHabBkXd0iL5mb108UFAlYgp1p98s9FMn3hodsrq
3M6VqGaEPaMWKqRgoDUEzsfpyFup02WZ2u8rA0i42sqvzGmh/1gm2pzqx+B4KeoMPBwSvzLFuKjo
34+Xq+ZGJOtVEZICyyIZASOyeHo3dKQ73fDyA0gcZTF2AEu5a2QFPbjQ3syntoUMm0ejdtCctAk4
MrhgT+6/Dxf5n+EpG7XFDIVvTcGqvgTaEDHRB6R6isWrveKtUxBjXy8FuYn962yb/x48BaU9z920
ilo983YpGtSK70Qb4DFS06IAjb+JbLOT8cPlYHkCjloj+OEa0o8hp7AshqJxa1pYoqbOPrEiSKPz
eMlMRLJsj6wOjw/UIR6iyH8zzV4cWTnAHU8qpsavCgRYJ5RQ7YJ8nw92yItCSleIEMhv6iO71Hzr
3AXFjR4CLopHGERVVLbiTbbDqgMrO6a52P73Fq92lqhi6TK6nRpI9tGE3LhUEjIvOC4GHl+84wwT
nJS/KDmvxhCYNMXw8NX13T9H7JfrTgrpNjQmgbb3mEdIfnby5r/NEFxUMuuhAUE1mFzXEaRSMN/O
XIdb/uJveamZJVpZlqWKxIWCcHlWu6tAR3nFXXZn8B6iTfa64hrmAzM3LaWyU+AmHn68Xd/urcYs
FucVZ62Cyy1kwVQDU0HrjurkEe3W3ExwcDzOXpKzwX+FDUBZgLxqgFofDyUKedAu523rikFH1F1b
6pKrHXdoNw1k5XxnMIIw3bOFUnHBNEFDYmJ1ylkQywH9jdlscgy8TTtX3iy3JOWmVmG9dp2WjHT3
qFQKG7iOCBHSN/l+0GeogXHaGZ0o531SIhHHkTNxTGHr9jSpfsHhrdRVcHCjzG6GTqihfjaG17BD
Hwr06Da6/cvQfgYdUKBOb8vYit/NIhk5D5QT1yqOdkfhnk2j9YvrIMeo6KVOelqiO1/MTWUoUNTp
JkFzBNdS0orVTb2Lu6FnktvuSNOYxVvw8NOGNVMlK7v2s5xry1Vj9U+Qk7fFP7DhCn5FhVmQcaRt
ijKqvLNDpgP1/4g3cW+JIFNhSLqFCdPrtDUJ40B2bvqDBYcDJ1/Sk+H8IZTp7nobNttJvvGY4NBq
I2wbimnAADoGNj6tWrLNRSfESaWU8WNu1Z7GUdlcAsm44jTBenrgL9jIxpGjhtyoJWkYHv1pPHIt
RAl7C+fa9/PThK7z4eIkG6t8KRU8n6HgkLH9u7ZZ5xWAC18y/CPcGh3gjYFcFhTza2mMMeH9wnq/
EUB9cSgJmHZp9+e5I2C/1bt9gM5gZFBOeTykFcNAhuNQhh7dHSzThwPyg6lk6ZZTv2ILld1PpeRK
lAqTP8fL2Z5dMLsLhnl1yZoxq4c27n9uC7VPQ5tYKbahXmMejJraOTjLKbaXc0PBvsmT7N3k7iKJ
E/4QrU5K9ahvyPxworJt81nk0CA24ph22ANbAJv6TCNdAGMj9uXJI0TUHRoyZjfKFDA5IcO073M7
DbQF4rGTfa4pykgz+52fJ/jlYi5PXxgCeJRp1bQKGb8C6ttaaQWo/UywY01OCTpP069wOIhonkgL
Jz39NRsWIFQxpi50W/Q58Wmb+MFehYL+uC6O7RqY0oyJYqd45J9FMjNz5vvqccURAnu2G8852gN6
OKnuTC3wWKSz28FzJr1MRlvKcspDfP52XjFoMTHf3zPEnhC6PzFwK8disiwdsDNwJfq4stSMzR9v
DVPk1V5m4paFmG0GO9QzzAoSY4Cz5D6o4BsDbcHH4OD/hxPVQ+itFfGfR2bDITtsG2HBZKizIS7D
5WCAeOUZT6RspfrrNMc+QBussCFFZXWk+RFIyznJQJbk4knUFSO/2rz5oTXuFMCRb06e2HPl3PrU
+h1/8OL5yWXkDMAYDurB2NH8eV3BV31cvtD2XE5/RjlQfrY/IEJRM/qGlldcJpDj2qYdslXx+LpE
w5pe2qct0R2wdbDGzdBfr7UWnG72Kbin923BvL4bQdr1n5oT7gBMjsII0ivM9bxzn23eE+L06WbL
zt13jKBtqH2PyZlaSwp6ooJ5S7vZcwgrWJv498+VmsSUxazH9O80jYppLDIaa8OXLkidCU45Ky2y
mv/23lvq/deMifOWROWCUJwGP1ZITaFtjqqGwX8TbrUtVWtWINaE+7AaXdUv9+8Oqd04tNPa5rw9
VnRqJve1Aia1Vt2vLNmRZOhjdDKWWEiWAoCj8kOE7jJfYrwITWz7tiZhqnvmVF3OMXIlAPKi+Ihp
tpNXHv/NJfzvqrZ6eJZUcMb1YXoNU0N3dGi0aQIxWqAnA06WpKkolMBsAIE/OfHyIuszoTdggYKR
KdENEeL0ETS03GsKP+aNKxGnLa3j0q0dnhIbOZu/hwT+t2tlBnM57yotwVIUPmNwgd5Xq/ROAski
MMj3s1WH7+n0hy7aYc8ZZkqX/TCwtLyFK0K8FWKo4rxDrSkyU5k7FGdmyELoX/tmc5Fy7N5sjD5t
xLE1+156dfLVo8W9ukmdeW9IcdhE+9lPCxdFMRmjPRRBRVZspBojJsMy2eBYe+r9NNvnW/LRaELV
7n+f7y5cR8X6yAq7EJ9x68k04tuUklqpY7VKAHPPUF7eJ2H8We6hE9z65JFx2VHwRH1P9mIEXo6m
zsmkf84c52MK0GHE20IvMc1zfIQzhMdKSHG6qsGdK4RCnCrOPWzHRvVRFnXS9crQqb0vqFAkDjMo
qofIxQYE9fs/WBrauxD+HLaF94n6X+3vRRnipQFz7pGG1VX85PzMaNo2c/twF69OdLFjqh1utxYT
qNqg7Ztl9QQ0qRn/goT/D/yza3BvCxMLT9dwvrAVMayOjf0HQ1n7KwFJ3kGUwnjcd+Bk3nhicBRL
YSPK+4j0xufKXNPmnak9D/OYRwY00UcZqHYTSC3kNhC98fsm06E1SSbGJnsIOk7Wfj/de4rgP3on
bXdGbp1fJ0EsStWjGwummRAw1KoIJXVg3tOMT1PYYgfuR1q2FXFtHRvu5jkwmpStlc1X3utqEx2z
3LVB1tz31SPenV8JuFtThgzgW7EP34XVNoN1UrKGumW4A3AwwO3uBHD5ydmKM5pvRA/jABnYkOU7
NW8KI02QUP9rNzvQxxYpRf6CzsVflbifcPrKeM+u8u1TupsFWUDH3ErRf70uoOCrxCctrjTJN++w
YcPNGluCQZBVmvr/J5tdjoURuK4nVvnyLGvBsaHmX9HzbzyHy4UgNr1smDlUtsvqvYKHTpMyjPPu
tuVpXvH80yw9Uy0D2xyIuySXOzlEg8ncGe8rGAY59EW/U8/8iODPxiNkGOOcGj9JDjR5wzYdgUcG
t0tSCo7te6c5KYllb5CPySk5nzz20YzOY+80RQUZkh/nCXlWiY2PFvW2yyG1xqyfowvknChFussK
D2IRzG/Vd0I1KauHATnL2TfH+7c+aHjIJGXCZAqdrJttBCZTBbnUXnP6D7Bcuf6Dlxzhm48r1Wka
NKVUp9h7qr5rvCKQ+wsROPBXx0jZsvX93cjPcMJ2GaQvxNhXCXti03/5kUPba0SebfMTh3bSvtfv
2cJ38oMOaRXD6NNEmubWnpHaaq+MD/6nkMfMM3r6M3NzEhFvLMF1uRkvWP7q4SXyyqZ8j1RjMcWc
uiYayuG3qqtjPlJGkJ7PfAZf65RZ4hv6hZOhlvgJd9Hp3ERlj0zXR6w7KgMVu05elGdxcp3mtrSI
qoGhY7BQUv42kFBy50lPKdIbIR506mT3hcTl4ruypqXghLuwUw4jCOMEzWPckVuakdpLvxToLGS5
ldVyHeAHo1zzGjXCBKLyl+eByqk4E9fqjyW5eUQudEyNQtBwTg0mq9lTIxxkbGBn7cv3q5C3OQGn
9kI0gxEtFyTJ52DQSMcwmBE/vEj5c3DejsUHEOqZLgucqxC4lUqz8hRhX61eBEtuUS+tRTfRuPUx
BzMu5vXGUrsy6wZpSqYnTESlD3Fz9ERIa1FfFvc1oKTyqdKJX85lNymIF27ojvlbnwwjJE52nB/q
Peqm05qoj2gvAk6QjZitwEvEOWVg2VwUNXJd8L2MIMhca/Vlrw+44mJp7dS2XKQ2+DO5yOHroyEB
XTETj0uT6UsXnPuR6cyYTROyf6f0xPwS+dTo2lAGSOvBI23IQDEZmfu78ST8SULSDRGS3OzCvTp8
oY8apqXJnB1sYhDsUaFed266gPd0bws06tCBOwg39GURXObvuAnFzrGeVFlghTYW1d9pRHyrBach
NyWGHaRngbai9aHEjroqM2jBOW0hVkgAFkUURTnHKqWjfwk3eoMxTmqj0z2D3sd1x8eSUcql5gXP
pU8J2/5rUHADg2sxUbhe1vDFdsI9JeD4ZvEdTRRdTddSluLGHMwm0vW6c3Ab9u2pDERlv2cXpLrf
NZ1lin+8Y4Fz21jI7yPoFfUR4UXxZ8AsgS1HJoBO7V9IDnUD9m9+lomNIyY4Ha+LPd3gjemdnLuU
ElYg5aKNY5xqYnaSimVj8WNaF8+TVt/VxTZ1uUe8voptDQS3ic5Wbk1dW/iVuAy3w+g+rTTJ7tLL
widf/c/m5xCuVnrHcMHnFbXKdyZbB7+UjT82O/IxxjiJp3CjoJZMm3RaiOAlfAqKOWy2uUfoK+Pk
aZMP6X/uI7MRVnglAXwnyokBnRqpUsc7qKQ7sqW+om1MjrrdIRqDz7T0tIhR+v8QnXv49yW4/uVq
DesPD68cfyr8iYPQtS7ZPGIimFPxKN7ZtP5WjghHdChDHeqOY/f4XtpFSTPOYUCyIVACucsyBnyY
SLbkR0rBCMDzzX+05yP9VIMtSb7uCqsML8pweqEVWkrnbaGpiXTvs3sPkyUl5YZw4lS6Q719FvSd
6cCbd0J+uLU3i48ygm07sGFnrNwjLJLoNyimy9Ei/Y0Ch7qiR1jFD1IVid6go9Jv0K5LFHfGhENw
uX0sEuwQngM89J5V3K2dVEr8usDuXUnQSmBMGQcK1G9ZprmZ61kIRGLIxt5i6m9mAJwZIudMFFnW
SVhQDVfeqZaTJhlQNs+szLbY6/rNI0bfg5GskJ8ye9lIB/cWq0o4qx/5gLv8reM1+m8hnm0dHCdr
CNdsdSnT4EVn3FSLHgsoE3TTKd6oh63OlBFxLCofU8HcPnXzSrXwnxRG5aJ+LY1HCwUbyc4ig2QP
+DOcM4JyEiNjC+ajSWjbga2bvBOIGxvH2JXOJNbgElnK/utLCHZjDsfICGQ8cjTWUbFFKtV3NqcG
0DYaQ3UHCrILfsIu2Jy6YZTvaWq4QgUQVCenf9j+UXxnJMHOaldv+eHUb82QH1L/dhz8fwDvqhJ5
Bf23XolXLsm2yNRLhBEJdhGXi36lFgUu8j5FNuhfjNdYQBa6Hg7a1FKrVujNTeE6QBRRoPnHeJ1B
Ilq1teWPDHWuu1bR0EOA8gfOlAYb8nHzFDJUJRwLerIn87jnKhYSStGJUg1StcwDDAkW3KWERg7J
sevC+I1/Y5/eLunS7SVhP8JtAHtz/QUchGJKDI8JcU1Fxw0UorR0BIEyh8v+et25PcIKZaFKz42k
o3dutaMShygAvtihQ0Hy0JRdRb0cEfS0Jh1hBaVwDilgo5SRe8fGhGk6qWfLCFKTWLqWqEwSKOVr
jPYOOmYI6jhyERqTiJtDuZAd4XjENhBwy6Mj7eYDlF4/k6JXUaUcMPRl90M1qPK77bp+gM07iBmW
7AvzjOKKx8jjuv+dnXgsa3ARiVcaSZ+6PYyMSKQOJJ/JyvMD5Q0pcJPkBiOC4VqIeUJcIvlKmjP0
x0GY0+YPZlGaJZbRGCpNGXMtTWurBnKD0QwWAhCcYkoQXSbnQyHTBUeZgZDPGiGmMRX2eHS8q067
M8scX8D+jyUhssfbCN4xTEzFO3haLR0XmU1PLF1rJr18Or6DWMTT8pRO133qDa7X920v/ONhhDgz
8lJ0cPsPiOCvmXzpgyTwvDYyqF4BozkOJcs5cIb7wmZXt6uIJDJCJRMDVwpt6BMmcuuA/lJsGwjS
/09RkVEGw95tw+93NPr+pUXNP04OaNd85+nwoiU+R0WO3k6XQhn+DY4aZtdGAr9ZWC2DdNlZykDW
lgzySqwYuS5YHaJIt5gXjrBVbzqsTkB6S02TtBt+ytTy3zgP1/Es/mhZBQWH/VqnzeSaDTSy3TYW
s/uLQ4VyCUToV4uUc/oGErpAFznXk2wrdpZ9QnyYgmrmhiDYK+g6WUxcWxBTUB52T3hBg9bkf2zg
SCQqT0PutbNA66myozgZkLu74WtwHW3pV8aGdJcPo5EznyeLvzBNIFy1LnHi8MUN9imzmKkCua9n
8q6K+ADWcmdA0edIG1XJDlt6XiTrQTMpJGaRA0xFSwvTBWbXycfmUxluW5IoTkgjTXyMWlw1jlR3
6i7XpnFv8L0PFGyCu4j6wxKa1bFB+iKbcPQrrGZMU+tme0FU+gwdIsO0GMkCxin1a0D5LNywMuD4
VHeMnVdUSZd41tAACQgsNPcPJ4t8fG1gSfcudyJUTyeJdfbrGLOXZcWNEQTvfdzpwmfxGidlouCG
rKfPeQffJrjMMtJi1CPJyhKxnesr/ZGK49v+YTvYbIi1t+M3j676JWnvYkrM2a8YKXM557trwE8B
5vvmV+KXtK53TOGgrYbTBNKVYF2C12ByswlEIy9MTvVWiXage3NDYZfMdLWd0BcTd5x7BtA3mD00
LC43X+gUhXkgKvt4owDGbEuJYgXJYFYwH4NjBhDqLqqa7MbTZ0TDBBa7Vsup0rvgTZFdpt4SoM2m
vA6B/f42+HlOicWFayR896IhNi72GH3nkaIHuCr5VWJlAED9u7yFVBUZYEhxtZy+Ub9adGqbxX5s
9w35XpfjYQZzt0wlWLovmua6HHt26R1zrH+WSDhlaV/3x9Z6/WDXzd07kZA17wdXB90rQatVqIi8
UBePuedZZLw74IXxiCI99YNY6Hekr6KKdUyaWGFZ+jHv5F9YrEy72vtWbIfM3CM5Qinp1FfIx8vD
b7G7GRc9CJhds09Ke2g+7LuOAtmtBVigulm8o6VDGe2XHf3ARF459Bc86Z7LkzEXUYKsppUo+sbH
EK+9b5bp15QJmAXeV0x2p5lpgoaH0+QUdFTXNXGu1cus7sLRNKTHXJfi90b7dbGJr6qp/J4bNrm9
1XwHr0M+rV1Sh89vMtQT+7XpxMD9Ev7tLo05SNBLm3myJoahSOY+wTNlW5PMTB3DYQUz7/ht1pFQ
qOCcNNLMzaCtGf8l5Zby+GY8NqHisvo7meJlAdSJn1ywC77oNfh9GLB/JXDuWTXa+DO7VG8lSGas
5jQbaQgKJpUm837Wb1/18y+3kEJGQ0PDTXJtCckAPrErFXkliZCZEhtG1lYa3Zlxd5e1HIzhQWg9
wZ4ChwOShlH8i8CBS2QcMZFq+fAQ68QuPmG8QuQePnnB/dae13pTHonWPudzT2kA3U3SC6b8SOvk
733z9FXoPeuqO3Tnd7Dic47P61I1wZjpbUa2euERteHupIF0FecAqXSyJ/ScI16gkkuSk1BYCyHI
218O6H0Fp4ZXSMmJa9pnJKpC1APIp/Un6kuS/E14dkz4HbfmUC09DdGEtwS0Jue5CPoKg/75hUd8
poaliuhiFIMbUs1mnf6yTkci2LE/mBGuS+N0PXnU+laIQ2v5mjtM3sxi+GB9802KChQCN8fLYU5S
c4YxamURT/tPiN1WSFSjXrtEtpjPuq8VOfXFEcfLoReaEi5Au2qa+SF+2/EuxprHoNTnjZki3a2T
Kr33dyRBvtRz9wCQjFs3VTGiRlcjaVtP7C2TARDcNMZRsZ6uqxcn/3wkj/u4OhYWuvBs659m6Nlk
p1QouRwXN4UZLbjlLZK/50GhTpl8DaD5Vskp/jrjEn6MbNgD2QX8ZgPf9Sf/pwJ6tRYFAoBiIgNf
BLnZ6Qq4v250bFBDbaGjnz/RJWd0OQl8l8LLIZdmXFXl77gnG53jj8lDsWPJTMejGFCdwncmLKr4
4h/TAFdDwYd8NXar+WnWSCQkoA7wfaM4OzTiH5J8xm9SUdXXZe9X63dWz+qZL7oxLpZ+BfMC3kM9
wp2yKjpqJGlLHKMttXSypkt1UckOdO+Q9Ep60WIr+gWX5LPpYRe1twIec9KlHuGgW+TV+xTNRdE3
GEhS7n39WBigSqxyhcV8VgSMl7AH9z/oJ3a9156YnwvQxkB6peblNZioX8UtGnvm99diQp9439dG
IUz2BSKAvkMVWyhNWJ5SFiA8OaGFrxtafjIGbpBiH7TsSteZ0x4JwAwvDjsRG5MxD4UbOUKPAPTI
ge7qExvn1+H8n/Wr3PuEZ6bwlXAWCnulaRRGl//5wRLndrQYMVYUCYyas+7LS8PoXSHR8pvRcyQv
iSmeYAQOQ8wg9WFQfqxWL6WeLT5FT4IrPhxpXrucjo3rflzpNBsn5qY+zNAOCN8+BcX1eDQgAxsZ
fy9T/LuijkwL9yf0Yh/SBrHj8zTaba9z6h3tM3/Upa3djRnBSozkVXeBRXbDX4UZ9JHodIk1j/bR
OBy1SB5irFcjkSlpCvxioBwrZUjq3DQvyUdujhA6wsQB0HO2T3tGznVLnNDScXPp8kqjxBhajzYi
pj/LFxDv7QKz7aoFE8rthMEO7eNN3/R+str+S+nqr7aSCO4mZg2G+FQGMjtdwCpN4D/y20Jy7DEQ
LnlDUU9k4Lms9Wmgtu1R4loggcDG4i89x6HofqSfZA1X9+bUTgQYLvwT5m2tPF884QC2sF0dXu9+
HyWSP++4CWZQY0xEaVhQkewW+NpD6MGLYO5s1tLT6sg+mG3lhKY7om0Zcawv0PPib+pDbC3RD83R
ypD2SYVyR+ZS77KQzusAGKXXHHnDWyCT1bJb8UuPxcFwFXCw6hx/uxMum+JhbVGa9KQ0Y2zk5nv+
VHNPGfX0JcYimiRoHmZ4ih0Er9m4khcUau4OYWdRZN1z1KsE8P5mJL/bJDG1gNQke2qQlEs7Srdp
QfmxW5WbVPTfTCEtHEWChKYEo5fKI3b5gnfbI5OtfH+6daAbI3XhXUVQUTq+5sId66hYkgR+6+nu
nk2FDL6YDy7TKRLCj0MTflY/nQleYptq4sA6kFW8jvWqlMzYVYAyziPPmgTDxSHBcrIAGAz8CxC6
DbgJyuOb0QO3lhySG7Q5CK5sygoi/JpS6TAlyea4TfZlu/xeQqVwXFE/8rlv76gESblWVM6Izcvu
ZL5e5Ltru4+0fdVdAMRl4oBRoe+bV6vGeIu/Dsdbc71HFVKAcBb0WNXLeBk3XWsj6KeYeDwztk/Y
LMv/tRjGSubK4LLyp4aBHRCOq0h4L0K6iHqNOSjhlQsw1MDVQe2Wcvm55hAvVQyEN1JElS7PLV0X
ABsKisStgObm75WeGwVqRN/2hl+fmeLUKNorDz1QAyzHR77s0sv6uxXeFQRyI6ikGvwKTmwP9Plv
ztY2Y+Y0ruvFjOu66xsomA/jtN5AWDAgNuAABJYBf4SCfO8vSqho42M/34eABbHwVJVH/Jz3qopf
QI9Of0KoXc4X+DjbIO8BsPBJN41dSCl2mSsHmcTy8DOKP7KoPfwSsZo0SvGcQjEHQ+FHr0HxTLdx
YP4YWVfRsElnnegsWKzdZDREZPLxVtA6HqokVMCconxXwQTznc87XIA0/vjv+RfqUkA0iyh/+tmV
UAH86E0WF5MgvgyIVa+KqFB5hRFnZkcGR48boVabBx9QM3ZfFr0MKf82EBJFx6DvePXXLFSccQTX
6/BWLMPgloh6CdwdWgbVTozDFtqhYcrUSHV/s2xYRoypc+RGFh2iy+TDKc1fxps/VJPi/Qbp+u30
HHWi6bY3oB4tg+AuZ6AGRPN/4/1SGjq8wFhq0jpEsHveF7YnTbDn3Ml7RYUTYtDGwh2msZmZx4u0
aK8vO5gL2hfelo5pD+cS/Czj7f5HUpEhthHBlcPlmEi2k9kQyqIdF1ERBoU957XG4uPtKuvn223h
I7vCL5e0ZX6eTnccOwCYl4/9v+NOmnnHHacRIwlosIVmbo3trxpMywzk8aVXs+zqSeynak3gCWov
P1cC46Jao0ZVkcu5aoe4IW+OVMSOfjkOKvhhtY1bWbJB3D12QLFs0By5hZ69EmyK03ICqh6MZ/s2
UwbnlaVdXMOeIhKkEXK6GjsUYsZsFYMLNxJLpPycDaQk+wQ3Ht6WJmhz7Pi68uVw2E7bcQL0v0FU
EnmgKzH7VY4sL4+yMrV+/0w4Q2cUr3O570cACSdjOb3reqpezs6xvQ/0DSS8d8bnb20/m6xI7IJe
xL8XhhClpL6ZuPhLeevSpRPY40mtgYBu9REdxmYW1qnpqyZNVS0lkt/+CI+i7k+qY0Gwu3U7X0iu
yxIrTtNUlJvHE8pMt4HtcxYXufLVn5Aqj8nQ8MjXwTbgPwXfhwundR/6mNQerqZ0y34pRg9EyIeL
vXYd8vfleqSQwLSxmq7HKyoLondbUiwVKgdNNjc1lulRIw58+gRPRMU97ODIq0WFtXBFZRdySsVV
6uycUXu4/qcW8gkvyuDoKhjPV4RKH/gab6UPRgcv5oNsKUcuVZJkVRIY2okXtt751uGMoOQ2c9tt
5jCIgdeheB5L5JIgL8H7sgYXT+b4Ew5ez1pMkxWDZhRQ+NX3zayJ50yocQnbEBsNpXwZr3aNJm3r
7Umo8nwI9JHX6tfb9dJQDY+9vQ5f7lzu7Vvyh2A16wIUpo8AOzXZrmkUeVnunGL1N4o+1idStYLo
9avM0tpCgxuSHn4+hGqXH9OugQx92pr/ai2EO+KR6k7PjMU/ajRaG9xe5epjPG40oYBsu922OnnS
g8ThZP8BZ9E0y2sqem7KI6uPUCzpri7Pnc5c9yB+wTW7bKkMH5mPm6lZlJv4Mo2P118VLToZt1Ku
1n0ufYPuGmntJvUVSwM3nrZCb2ua5oR6LPQBV7L57ajyPqBc+OymJLla1gEuNnQ+Oh46MGszQZcP
AzseFjv0D/RVz8BcT5fWPXi3oSuTG8TAwajRHJyilBRNYKBnrkv4Z9YbXQOiy3JK5bB6yafbC6LV
PfnHIr0jC+eELYn+0NHO1plgYt50SDewwaBoHfSDNsIwWTx7ummspLiPUvrtIaz21yu/NrKBawzj
AUGzhQlK4jY7Rv70eFgG+dfp5tVDCf3JOlXdAx9yqC7xPO1s/53nbliWt6+9S6Mlyy0JYWY98q/T
49ajxqX0kde19G1+jgQnwG9kwFG+/Y+J28UabvMRiKgR34p1/IfNoOMmjjWXhxeAWt6Kx9ZJpD6k
fBehVUJ+2S8ifNT8ESmyPD2CQqyqfj3k2tD7euU+ZAcbLoOhpXAJVtrH9i2Q8S2cdGKLJuFEHLC1
USHIj5BjLKVcY/rCpsPq4NDVHcUbLr9E7IdbOiEFpKYjFWNLeG+wSgK/VGBPsEZUTbrtRnSo6R9c
wzAEI3pLE9CLbj6do4zM1f8JrmDvn2xKjmggQnXvXZ10s+NehzWqEllB/drUlGQNQxyl5XxQwyGQ
w+EKGv/s02tjt0FJPsjafxcl25NPDS1ZOGOcxYkKM7ADsBXvMceig7JjUF4WMo0vKWSYteHUqSqp
eo1HE3NbHIzJc35A2vVa211983tUIcFZgbBveNqK/6Y3Y1O8EOrk6qZIg7dzxIjIZXfGEAjQ7x0f
1wc2m/lb7OVwA3/DumbuMJcC4OPsDVuSVo7WS1KP+YaRsaFRCIKFqqvElo/qCSbJdceV+ysS49lP
qVdv5JYVg615iWJa7TiW35TAnke6p/+W5Tc+iRU4vs1u6ap/zRrfzmkKm+6Kf2jqrt+J21QEHkqr
O4sRkxz7FwapPBt39qCAsqCVmsKvjZ1gDFmKo/lGgR/A4RDk1zzvGbRdItORK704l2dMnFYpkE7o
2n0ElC3ADLgbeySxD058WBkpfxwnxEd8lEiO+jUeHHxSwsAVIDmzuE8lM8YlhcJ7ZMjDSQD8djt3
ib16HibkEOVo85kjF78/oNV3hhZ2WNbZkSH1Am8jflWpTjAoO/xj7+9vlRtj51/WhkNLlNicR/ac
avqNkT/X5hHN7h2w9CvCUopQPzq9XR/LquhdP2yu3+vRV6F3Pu9keDfU8h22Qn1rPBovWpE1jjXD
RlHkGQTa+VJYv+hPa/q6phwZwsHtwIm6/lqMbd+CExtkYIPdEl4uOCWydVq8DjYpU8at4xLHxtJ5
gl61VGo2f8H23YbqHNf+qv+WZq8dlq5xcpZhyk1sPwI2uj06QfeZcJ4ndeFICNnTfkuDgbIx+xut
WRI6NYPMOGWCxJSIIIC13Wz7Y9Djy7EkDcsTAUfMFiD53uDRWZNNqaiK92ghVq6bfJDbsWfyxvCj
Y/S4InC9dahYg08RHQFRSt62dW+V0G4WvukOS3LpRAAPdsZIvcr0+caCwXdHw/5D/B0jdnWRg9Au
kbT19DNsO72Z/c2u7cYLNjOxPL2PuQZhepKnlEujlLGaoBddXZ4rXTrSO4fpJZLvehFVaYmLzt1p
UiTxCe7dzhxXnTnR9bRaSpqQqOqiX6UL5sJu+ydoSsTIDouQdil8cWk3yyRCybgTDtosxtk/3PBG
JdBk4Nmsphgknqs65/lm1E6wX4Pnokxm9IJ2cPHd9SPavL4ZofgsmNvFtYz0SpppPnjsgjGYcADe
x9qadKlyXHxkP9xXdVHIYwY64jqANznupx271E5uMLZ0a9ncOW6M9DR6iX7GD8spXNQAZnNPUwZ/
LWT5biU0RvlALWPYmmfj3r0TnNFlkEOh4rNv22C+C2fWcu+yeWtsxMltkL2Bcu3z61c8lzvdbfm1
0GpJkyjLVJp7OxndcgPfpm6bQ4Lh3NobCywKMcIqqjmYqXutwuJ0py76QkxZaRPAZIkbHfZhQqbF
uXCeQx1v09HkdcHG3TagWw4ebOVoIuExUnVkmcLat6l/smG2Xsw+vWnrIyjoa8VPU2eKA3SJLUZa
sMt4sno7/2vaox8iNLFV+Rz9L/9QpelzEJ/mpGq6Yeq8Aa5YABkdHYiSt3dB55dJphXuZ0ETnuQn
qCDoRUYAjfqhGwzn7DUKapy50DoWG0snag/6xN8YslJKSmAZgf3MZKkeQwjL/H7u0fEWN/i7IzW1
Sgv/J7wK+yLk9h4aED0GUCQjb0tF3XQD9W/zUy9Lz+1TE0jnzBZN4y2JgrlbD65ewSoMoxgnQ4F7
NNmKstAIP3yihwuom1O/dJJPdjTeQ1mMcmgyBCE8u6TUp4uswYqSZzMw9c0yzJqLkz4XRh8eA7kN
+wStMzCg6M7KehoduoPBB/g+PVA+X3XqmnZJZ11azCVcZSUfFsWzPI1YYlyrpHt99+XAzabY8Adr
3B6J6TKHlD5W0bW93l+pEKetvFwUDg/LFK3q8CSaG7x59qduGGu5XuAuy2Qn9/irXd0K/YSxkMs7
VVgtrvNJ3H28OmeTLRH8O1ea8nnUIU6JqNNEV1W+KO4Ipm8D1bxmwnWd3+qlO6pkSYQkvE4PgUmt
WEjnqJqu/VLolXXWx34AbVgKmU8ffsD0d6IMDTJBlPjtUSfbxeBSOoGUoShwepL/K/vpAp0urwby
d6gw6jUa2MBFoDYeTEo/8ihUZVxq5dI+UKGsv8mwpn/KyqXo5zglJVVFnmjxx6LurQQoqEhs1Hjw
wW0b5gvtUwBXZcWo5jSCejb6GjtE+/8iVCbFLCLKvHqMQs3wTrV3HxKGNIsnwP6cgYcytNcHmYfo
H0NxQQiprSffKU3496IS0o8yrvy2sGC7lRBVPZqUDBIXw3+E+zJJZ1PjaoKZklpA3EU1TrAi9hTZ
2Ai9K/tMoOY9gpnMVveJ9rHPU1KCiffBmhQIS3DUxvxcPc2FaDV62Ak8XxWm2rThNFdqMRCE/p1C
0ib7CVx2lEX1eDzdssvtbiac16LLMacFIk14YdUhb1rwkHGdNEjlmJWJvdv5TOmfjt3uDfCXkpek
aiWxihXLns23DNmNH+IAjjRnWXKiJ6sqMf0MbE0zjVSzV6+r1aNeGqNAlhs0WldWDuXgT7Ncaeru
GbpADYwROSoOFkY35WGQWY5IBGEJ91ibb8N7z2FX2vV+CeQAL3lrMaoeSKXu83aqeDCYv5OeS91D
LiPdx24MWNAmNHxCf8Ot8VGNXw84bjyEA1sWi7fN92PCGKhe3lMge7Lm4W725KaJkSN6FtRpoibq
QMLoiiGyigqeIjs7cBr33lamVfiPPJ5NTxJ5KHq/XJXSqj+s7UDTZ4AQcgDG1G80nawe0GiCGwsR
o+w0gcpS3WDD7HVHAQfKHT59yTBZAU4dSGrdMzyvR8zI5PHpdxAc7NAkRh/ol8kaV9uDyAFO2elc
XXA7KJ+V5G3+gE2Gsw6xYCoUvFukIqkOfU4ejy0jqEMLRAGDzjlECZ4x90KO1nGaU8RvIQzluT9S
IVTkqC2rVukbw8co59HXF62GiEfgAjqlmutl9lUQNpIlk59UOkkgwsEaE6o2aituv6GtHJO2MXtH
GDSVgt9kX3HuzZ7vvAa5FYX3oBKwOUzxOAkaDUzoiYJslmoPLufrflyoC1pwhXkd027QR/92PxKC
XUJJBVc2JouKYAumQ7vdcZOdnc3MILjD0yILAKl/84iPapsh9Y7fm1UgOWogfPhPcZVDn21HpKjs
UUp1WMM3wTagnU6/CoiDLLAasbOYJe6f9Yccg/E7PbFwK694hkfmwm+TlYmPuJIS3KlUGrAxYnH1
MnOG4stGIUhjitgOD1pu/kJi/T8zHW4f8Lzg8O8hm4/VBMA2FdYB/PDQRzN6paHA+5uBDl6B1G2n
KFVmEofjdqXDJwvjDRMtEeNrslbzRPv+/tkX5k0qoWKxny3/mPqOjSxv4BJl6NEkQflAhP0n86mK
uGqowJ/pvB8od0oqBu1DtZucBwycTGweaZOMX4ykJ0cy+QX9BzR1rypn77e5rm/qvnLx2oLm/6hO
frGKEzGYVt8gTfa4KDNnA8xj1fjHDnh1MlREBhIe1WZIrl2v+kM6HbRK9mdsMv6bE0J9rJkFTWH6
GpuNGTtrvcjg2mH9LsklExd6vwCiuQ3ptGIctW5jycChrGw362YubOnJbtPURQTk08y629qeeQI0
fEVMpMtxahuNuhgOUoy3cPn22h55EMmKbfO/ppooYm9S9l4ltxwqWj3B08st/I2zbh7a+juHGcCb
/Uem0qkP37j0s4POcJl9VNHHuV9Oe8mADTRZSDEVeSKqZVPIObxr0IAMOOy/BDpvB6l86vb0omkj
jkPruK3wkbZ9vwq0W1Fvu+QWiwLf+GPHehIVpocqSJyzMLbNqePZ4PACxJcI4tWzY5ELfPDIzKEz
QElD22U5jFSrkU3JJzlSFih7nruhJjJhrM+xxM9ndj6n6x7OwtjGsdpryscJZ6ZnV6iMa3hc/coV
slJ3aQ4Bij6W3Ijry0bQ9de1Z5oiqQHmnpXWDQw7tvmGarj4yrOx5QKIYaOnBkHCUWH6GiTZtxQ7
WC8HVnopXGihci98hN9LCYTGQz2/5jyN/mjWdd67cN7OAEgl8dioa1ST3OeXLXucYvEF4Bj8Ps1U
P1D5l731ZUBuSpMRKx9m/7KKpityws/mDv56oZAp5AzOiYx2GmLnjg326SF/w+KlRTldped+2bfP
ziS+8cRDYSIClaqaMnqXWpJMFhF8ndagYsqJWl73lhMDhvWwMtw4CHeanDUOaw+81G7tN3v7EkOy
Y5POYvXqdMiwEy/Y/18nH9izEd/TRoi5DRcXSf6sn5Up6qVihbSP2aMC0hop+on87i1Y48JzTSa7
ge0dqfneQsXq8MmRP6YuEp2HDS0TmjAYyuxsJM+M2pw/fxX2uFkb4o+CWIb35erecrhfW53YZUGk
grt+jrIMr8buWDq401A2l9mvqGO5UWVoJOY9RDiXYEvC9SdQhNg0OLvT9LAAaXXhGttHK5lEoiSC
BPulFHiuv5c8M7q5a/NbSsF/f83micn6tqr07rDaVG3qZlj+4vyKz1xRajPUKAJnq08cwJkiKvu6
Iu6zZLNZ9WvXLFNAjT23YTEOelqGerQhUKukipeQsJOQKTXLjcaXZZpR1WwK/Z08bOuIp41LmxXt
MN4+D6WYGKyZORo8rndBehXC25EDxbMOiLMIG1BXZO9Gcq8RIIh/nTr95/lnvm+QLiq4daAL4xWz
Kc69UQB79L8sM/0urfv0Q/0YbCcnh8ZausU7SfJhTjyrQ5tYLBrBG9bNA6SxQYAHlkG/JvKvBBLq
w9LnYB/vjSAS+2pQwc2NTpV6LS5fRmb8tYbW583BlC9a3zUDhM4drJd9raIrAk671czb4zTuu5vP
IWMm6+iY1D8hqeneom79hcIyaasBsvxPOP61WuRdQxZb+JjUL2afWvr0BYjvFVRjkS6La9sqcmj2
y2y7JDvc7i74xTuJ5hqKBeMFMBbHcJaCVpxbjCNdN+uW3jgZhSZztZxVf5G37hwYpG9/KwNJccT0
RVVokgOKGOjwlTkJhu7aHWSknK81dpnZUuNQx2kOXy4LlhJ9QR1rrl8PCR91UpMROSwcXNcKTySd
oyRYHcwUksOgKyHGHGkfp3UC1nJVf4cSeUZvYonJaHPIcWphPNOeTpfYm1CLpknnJ44Nws0K+Syc
Sefc05p+lVMbZ4zbyU9T+3lLbK3dNEVKQ7K6o9n0pG0cwXjy8sh+1sbFi4x3zv0kWJhR/LwkbQgd
lw+b1LkCDKlhnfSc36qNkg08abDnd3rEVQtcsf3ADX2ERSJb9IV0YrxnkMO5z3zTYHefWYtaX7ci
Ei4/TiKB7Nfq+TEJtYWKWX0yuAAQq/Lj1mQDWgASBM6bN3T+O+DOhsLG33zTSL2mmBU2WBSZCpvs
8sBVQ7F01AVolO3QjhIfoBWpOQn3avdTlq8N3fvTamFbigyaD9uti3bwe5b5XfUk2ddFgXUedyZg
/89TQkC4AgpkvJ06vTGiBeiatgFVLOjrfLWeQIbEKR3sl/4MOuMtWQsG9CgeFgk6LcqM0tiq5Kob
4KDRer13hMdZY1c5baEevaLn3mlFwaF4EE9BzcSU9eAa5BoCJJJCGRmoFjwoT8JhjvusQ8U7q3VO
cTyyhMh9DNrAbhyiskZiMflCcyOACOsFXQoMfDr+STr5Fd1wbVdYDa10Vlxk/0KUzNIycCEoTclM
bIo/te9cSuyasF9XLxIwa7lxqUqDIgDdxl2WgMUHtmVlKDnodY+ucn+CBSTGJuT+jUhSDCyXyC2m
yP7fR+lFpmYGeKjWaY6IZPCg79LjZx3ADJ/uIO0xwwQ3CmHMSctdULdmiCD/IDzS3AL3+WMqVES2
K76FpA1BaeqCN/LdbvEmF9RrfienzPgo3G+uTb0JZo7au3SP6EAgsrBqeQukU7+Mskzj4i15Wvh8
4TyDQOVweWVMWtNujVIrPST3C4r+3uz09xiDqkUJzpAk32EUKglgsrjl5c07Y4MRCppHrmYW/pZX
59N6Peygk4dAO/z6uWzXZemiMGOov9Rn56yP9oI6nlGLsE/D9HCU0yFvBD3LjVsfCYdgwACE4H/x
V60EYYlnQ5MYk/nG20bPmP/SodQ35QlCncUvKnq+AyOMk5OEIqEh2SZCpXgtjthT433KWk49EI7L
QGLljOKxoHGb9Ae5lScAFlZXhpt8HPPJxJHd2JYdmcMkJ7DfQ86S+6uoAZ/ygGweB1WLTzq5X/7U
pKkoMaOahe3qsqQmvZ98MkiHrWHSWSKAvmlVKib8rL8Asq86GQPJJI2zmDv7Yr/WMNgBin12NFxU
uZbw7i5y/SCnZBW1dawHb2/sBYFysTZ44sK7kMxml+c1JVahv/A9jkIEocZaRu8ZNQY0VxLurUc0
JgBFkpcJ2FMgkPKnXNPhPElYO50xzPHTKWCelgi/dV6+irdzoZ7boN8/jy636r+mTyjwIrlkma7l
aSyQ1EPPV7eNh7ZTHNMLpymQWPpA/+FMKTZyXtBVU8J9p3xjTRqTPSOWjPoa5SBlPYS0BQJc8A4m
y/vFEzSh40j4zMtTXRYIEVoz1xxYVTeiCIySc+jb5KVJEIR+nW1ce93mtu/QZKVAQdwXvID1bEXH
S6mR30FRm8AKoH4CZHml7JMgQ9nPb2MVkaRxT7JwJ4KY5YYCIS0WAZda0NtwAidmDAl4iTdh8CSj
rbEQNUD7igpfvXzlvMduF9KkY6CLeWUpzHA499gNVJITrPfC38U+oCZgB9jb3WhmZS/NvIkwrQd3
qna7HsqQVTO4sbeyuE+oVNN/JJXQD2UXghTVB7otZ/5vqYkzRlPQBbme4VbG6A8yiC4byxfzqHzL
i1uUEl2ZGm8f5dsZEHO/K5nUWO9xI7k55AAgLH9MyFZTDSKhvFACx8eNGyzWrkBvP/rw8C7SUk83
6bYcjmiYg5hEj3jr1CZsFPl8wDukbSEWwhoxa0V9L4vvdJ/5QceKom5lxsaQbN20vZsBuuN0eTyl
ZFj7ns2qOcnJKLj+R6xLPKCDQDnR6UpJ31P+Vg37y6UXLJSrLfzjaL9lo0CrBII4DaGqr1oqrucz
XEOAitoMtXqy77GqwvtzXSLtHLYTdzKIaUHmGW/nwqmkXUWe1qhAX5MamA6hU7kPii8WCFatMcjh
zP5mH6s+uvK13pS9aQdqPL8o9hm13ZFr25T9u2G0M48igE/bgxAlrmbdgDbofCjAVbuYYT1vlhXw
skN9/vUA4JpdceIeL6kNILQXkqexqq1CxWTs7t8QuSvY9fwf/MUsbjOiSmGneZRDW4VRMm6puvEu
bc0MKFneosV4eOqoivong4RRMH7lZWBYZn/DMyWRovEAURSyL6YXDzYWggfayVek/LHL4hrU9tWd
HhJK+RdIqMNNRWge5T3ZnJN7XLK1LUlFUYDcghqgsI/8Tzqp3cx3lmmmPaQ1/ZQIcKq2hQhJtYfp
GxrOBxRLA80E5kkUNSRFWPAt+4Aj7BHBmH4fJfACkJR0b9LWQgvKA4Qd27u00CTyrKWOq6sNOzTQ
+ax7B/j16HfyhyH6mj8oceWBG1U3Cree1LjIa8Q/hzkr8/sejcjpzTTogAefeidMq3tkfSOFHK5u
geRwNDt/r0tIsAhuivvZLRoZdHiHIGFvnRLRHb37asI99uwUhuuZ5dSI253oHayOuwrXpO2+cqm5
U4tS7E3sYJXR2DNcBbIYI3uQRELWzgTvh+Sn9E9U35dDhfMjaZ7OAsuqpByaMhjt4gZFpNhGl64G
ZulJlx1ed4MaobNHNuhbr6qCuEQ9loW3MonFoeqIJ725vAO5HASJx12pqxL+69pfoj3lW0OH5PDH
75c5OknWPrJqEk2IXf5KOaC5khpr4cAmt9YsQ6pvRGgRGBV22LnyIoYUSWgx1m4MnFjcZu2J+CNr
mL23uQkRwOtvRAv2ovuefAgr9q1AtPlSUkE045W7VCSPifQRVQWsMgaDDWYqtNqNkVKcLqcCOWjT
7AOsHXAhSZlvim7EKiRx37AXH9fIJJbF7GJJAOXUkGKy5fhIuNKdHZxVKQQJaxCoPCn5/hNL8mrQ
CmFmzhfj8PdFdbOLq3gR/xvfV4L6iW9SKdhmFxOERrp7r5msMsDUBbqH/jct/eEtFIp8luS9NU9m
TSqdKlg7xPADcmUgRX0ITlaRi3u1KuBRN74fWonY0vbxZqmK0RUCaqIJreWd80seEHByFzzanF3S
sXTJ5iXzaBp+mReNOts/ItnEWgoi9LlcUO+S2WbryAvnhJs/j4mKvtNB8n1Cib1/HZ79FhXIwMz4
NIKau4bA4yNlmAXBcOvvl8Z4jf1D5cMg3C8OitozMxYygknRNhi0iqJnWkDjVpq5Y58HE7ZGgMDG
szY16dz1v8/Bhq1IPuH5R0L/bxANW/xJyi5ExFSDfPJGIsHCyEhikQKzBbxVeSNDSSUeDxOUzO6d
PDJr8BwFiL8GSzx/ZRGxKlXpwlcb29jNxfxBG1Fj8iyNASDpAVUpu1V1i0MOzkTr7AbbpdOhNmMD
bSMh7EVLtwujMfI/dKXEa+++WWy+NJQQCAUbxgFqwd/w/gFt593lAdATzoVagrx+Pc3js6DwKACd
YrUetmBRw6OWgLxmo4YLWh7Z94+nqXEKt0kw3rgBbcbYFF1c6lxieRSH6JUDzkZZUNSWlRHx37Bl
hHvxGHHL3FkghMw5gQwlTlspzjG50VngX6mFXem5yyr3c5c39zCEX9A5l0nGxZQK14ZNmmUeKC4n
lA6MZz00jdfpVYrjzzMichAicyN8gpvXSSXUuyg3F+tw+nmhBnM5O4mapBlQCIkbDU7IkO4OPd7t
L//Xq0QfDXEees8jaFDemOVGdgaFdQFyn4NK5Yq3BMgIMdRKim0JE0uda2zj1U/y1Xhm48Sivp3D
3yOmXVB65sarbxVVwYnuYZxfnXbrXC2mymdoYxf8oqwSmKI+2eesyTAykW5TuA5Q60uK9CO7C8dE
MO9fwJgBpkEEqEbIMULdcpaX6qbpceZbjIx9SYDZavVYfi5qd368X5uxaNlrJE5oL4gAiiJBdVjo
59WzrvEwMnYhQvu4geLmqNIXezQwha757zTHJB6G9PBZkMPoG7PlZ3e/P5c39VbKQWZMYgrHnnZc
KPdJWmpMGlsC6g2xDxWXXJaXgts2qHf1/mBUp/hLUGITUTU8EZuXg2agbvtQKNkiJD9k0UgQbTWG
GLC+IRL6Y2LpnJiVM5ss3DLlJoRedK1Wjcvu7i87L4FLcSQuVgDjsDPJS9fOMshvXi4IAJc+wzGx
vT68DzwP3aF04+d3lvqfonK9uIbHjw9sbnt3Es5rdK9j9YSO+wpAoYNlsJJ+87NhrEXWDJnuKdkH
VukVK7GleLezSadEEhwQGc+pxjstYaGyQacJ9o/1uZoF/4902lyYrYIUTw+yEbNj49pYKKRilzbo
kkWOjF4PXImOwzq9gj7RDlcDp06CO8C3hdhSl4KETTluIe5fAjHcXE0M3Yp0GxzvKL+m9CGrXiES
rA2ksBqUar+W1m9InsM8yB68fWr8OR1daKbf108IIOgMLIeXimwl64uLYBIaErQSWQxtrZgSzapn
pO/AFqrf2BjoP8QfUSHfoBGBLNeMDSVLH6qBSRz8iIyBfFDS0LUZqvZisx8+A4NmAZUHb8/ZeWPr
LQbvIJcn9/7TI3Aiw3pVTCqaSfdHkZzGaI+dX14ioYojDkvPqd+vdJjMCdoFeBWb/j1PHkOyk+EW
x7h2xYrOiq5v+VdICxwV6LOP/BEN+qj7OvbzWYF70nmDo5TtLuqxL0B3PI0qNfjKJglytmV82ccy
IrbjEc9wcZYROt9igCVcQ61WzzxK1YMeb74l6Uh91G5BVpEd0c+dF3h5iy6RqyKnIzlgZKat+itC
OE1KtQu4jf0YrhINpuukq3VZAwlcDK6xxDOYNzRBNRdGhDIY55XJgQi9biAT7O8+EHmeNtl5QWtM
LP8ViI/Ezcs6JRlp9Yz2HTgB9gvkP5YtCasfBsSqpM9lWXffAMTC9XjxqheksXdyOtiesY47n+7d
nTxJr4U8OkpNtVyhYxhVGv56nqyFQXuI6T7nkbW/0SQx+8wbfZ09fv8zcBOGDd0Sf1VHNnB1havz
xzVBZ2uDjaD/HAVnFJsgIdme2NVglLey2Fp5dNNXsaOSP2P+3dw8thwwp0RFCZWECvR4hTq8rdUH
tobP0OlV3pY7SjCxI6A01MHvbYuWkq3GTxdrR3J4lu2bQp1Qo7YxHmPN1ZMT9ST8veL09k6GB7Sw
mTuZp1Suhr9w6EYcQnLP9t8JiVeqr3eXO29EMtWzYPgBjwe01R8D8Q8C0dxs291zHIPyF1+r0FjN
Pp4gQtyS746szvc+k010i3V8lQLBCtHRadNjpeA/b6hQ4GJP+3zMTS6HyXscAVEE4MJUndYQVd1J
O3UrQkng0JIhx4pb6jvmO3te0htQfW1bgaKbToR+IjXNt0TOyepWP4a7htJ24GQnVSVeL2tKJj8F
g5VlEjdwQIE44rYze1OAxd+6U+R+XJm0aRlO0t93qzKEeUrH3gGcFMJRAv54IdqwcZFE/7AmgFX8
DH0hAT/wp+HD5KPKLflqfB7jePFSCxr3k74DxZKRvZZq2xM8+FokmZMCX+YTtyIQjMjrQWfUSlij
eGFJ6uL6krzuMovXjQ0Z0bKZ69w19uNoitekFzTxabhNjD0P8rBxV6fZ0ZCYAPFK8BPT9+paKFU8
E3ECXt1RJclTnx8T9vAFZ5jNGb7xLlmjmpShPHeAsTNW2kVWpi6DYeme9vKAiVET81qVrRzyjiDl
TLcj0iVhx+n+mTbAtxVmtwH3KsCgSQznRaKzs8YzJRkeMJSGhP20F4oEoByEK5o5WZgmXwqOivKw
rN+s67y120joVo+fDCyFP4lDxmtE37Or4U281JfjZSi9+Bx914sI5LUVvNcPhqmdorZv0SGnDniS
BmMpHOzXtjloXeCVPEFDoaRx92huGxWsiNt6QTkja9pSQve4e4fT7xEbmBswGIUc//hgIxj9nIcu
cSvEPUyUZKmGO1enh57GdOeSfwg9i5WeKCzG1HH8CezceibCKZvUHLz+/IkX0w85hH3yPw4uZHlO
k+5o4DzQKY/qreRcreZUR2C887XxZsKa5lCpd1PHLmMbrNbTHDlMQWje+EFy0Q33nJrs446mxw9i
nhh3CyRlS6OhIDBLxSvC55RqGNU6ACofggZS3oMScQL1184NCcpUBXC0i2jnikK6rXRorWHINPxf
uPsZCLbjbGiS2wnZz8F/eOs7paY3y/gt61bIgJEfW/4//6AqJqJPdSQZSapbcltSCfd3ooitueIG
P1bc7EtIU5cJCq/JofP0xAXy4lFjsvxq3pDXiLx7EiVF0MSfDEeFT0RoMNrg+LFyMVgKIybIaO5i
c8bRAtonbEHygYBQGqyTCR8QsCdIeV9yx+BKclnZ20ndCV3tbsE8tt/VVnsfbtQeAbKYZNU8aCHS
7DAlTgY8m1hHDTyfocpG7ecWMFi9u2eNvzaHeU55tB+5fu9oYgcSitqFoV4i7XB+0/k87Q1HoyjK
jHfZQKCzBSSQUVcomYcZav2xo/NwDV0+YWJ4ua00likT/ZCFM0Nw26JCoKv+LwZT2IaoDCguVBQF
eaqBQfiQXjFyqy74MnGpDVH5qUp4xBaNwxbHu5P9ZzXSE60nfTjtzJAzd8k5VqZ7tuQDyyrHNTzX
3ykxZhqFURKuW07Ipg+wJlpJyU1m+8mc0klChgAal+1AwVZh3pF9xCGUCuAQLK+3Ok93uhSAdEVo
NmVCdAND7MmHlP3+YH/UBMPxHf1PVzM6lYAXWQlMiOumcl0cx9T1Ro4oqsZk3Dew2QZSpzRi15cq
SpjxzRFeiFFuD/R5KZD6nh4XhfFXWOdiR7cdPLiEJ3PNSdb4pyCTpWLOFNrxToa6XtvRHyQD+4d2
NGoWNaV0/MVyzoaHtW0NF1jUcr6Bi515QnEbOVm3YMtxOIOBjNpS6PznoKlZvpxRuvLv8reUbovK
SxcrABf41BMB31SGHZ7Q4o/jDuivrZwqebLnC+SdOjkIexD2BRPnGRA8fu/7PbFnWdehUsxRTVMe
gSyv7TNnLeHvOu6W3wCAEx/twpkb/3tP4AlegyqarQVuqctySgUg6R5GNOf8yOOsGunzaYVtQMIu
TKJZTfWMtcteeqU5m/IlNmYTzeBViO/fIUoPHW79KoI34NhlcVPP1eK2YhkPf1KF18Sjb1m8BDj/
1POAcPTRHXqUomx6L5IrB1u3I61+DLHErYlw5YF1xFzw1DoxuFeUr4eBtEp1NBx4FBwxOInMu4lA
7ulRlB51Q5MRHHOG8JAIN/Cr7iKp9TDu0hYvkg211D12xjRMzE2/4kpIYrIEo7V4O5p6yj0LrDp0
zKO3jNkcds6R8YkoLUare3VNZmvDWWO9tMfz6TN/6mVvxCIYg6P4N5h8ryhTOKRGnYWm4gYlNnyw
z9c+veW1c/J+YBDkOqs4eisIFE5TZnPJ1aRLc6p0h/uwFO+WS/q1TBDXH/RsWpW+pvJKDaQ8pbIi
1HN7A/ZbOxpJxNxkov0rVKVGtXjak6LDg/tinL3E7sU3+yX8T/WTd9c36sXRC3eP9oZquIJBm3zF
TLO4HiTic4N3dEpzgAmTNylzTbWwo0cPrJeYoVM7ijgk9gwDGH7U2xhae0uHMlgKliN48s+1FBcO
XjKHgNZWOkw+5Zzdj3w2jZvpVcO6ZSZgU0sYPyj2HCz2g82HIZVez1IsaUyjpsAyIR8HodQU+ZuF
3MFELH1usGmM90WVHjGPokOslKM3vw2Bjnuu/WvwF8DEewQ7PBnO6l45DLeesS4ssPqo3SX+uYvQ
gEcj9ED3rsMcH931f5gZeAjn00TUnNHqf71Z+jie0aM3U0+R9ushOKdSviDI5ebLsx5eH9xtj16L
rJX6uRfAqUfdqZiw79XqnuiyK+A3lOWodpiFWcPdXPhogfwlwQjT2QvX30dbUyHlW6WrJLIxWPRd
v8cTJQ2keri/zhqnjZ5OVdtZ0+ZPw5ngaUVI6MqsCmzcgjH4Id7/Y7aIoiMRDMUesJTbUWxiVzcJ
uvCHPoUjvwQ3QEpF4uyrffHORVbErd0SJdsOytq2OZDlpv0/J0YR9AIRXiysZ8dWZ9wte1KwfO5V
sJOzAhZsaYscpYOhtBQVlw0k3WkUhREGM0nKoZZOgw/HKocEOgfSbckMHkImUbaf26kw+mhJwqSy
JXZpMrcDZVzGU3mxM8WHo78eruAB8RtZra+vwxK8w7sAf7P3pQpU0pbACqm5Wo+gJ2PAmDA95aAR
uIARgx8gLB79ANmF5TLjbjN+YcfP78ukXd8lVpx8aEHsBWP4ne/yRqd4J8aqcnK+jjsBCSolUq8D
l+8MOtCWId1UL7FBbco8OhTn6aQr6QiGUXTtP/XaEVevq6tgVWZb8vwNP/KudW3WF/8sX6vjwYQS
rVDmG7KOGGhljYjXCUV+nPgHGGPSMESydBm3leIFIxOJFiS2h8w/0QDx7Qa9VbZaes4Ud76uCrf7
DZc4dGA5NkDxJ4RERjJWxluOVyJglrldwUmbat/CPS8mqGWkidhD5HZSsUn4K4Q370aXeW0hzRYq
uDLvGZ/df0gV9N7wZdlz7HPMHI2Vw4yhea9xIUChUjk2KKEd219dIlUAkUfP7TJW47sV30iSBvMb
mFfzsY/zeVKf0fKm5uTpe+XC6Rk0ELZDgpzxGJUxcydO/DEEo+CCKv9lNKLqgPyjRZULI057Jcim
qMREJwL8LSpMn+OjuM37sQSiXIY6KP7KmoF84E+iiMuxr1x6RIxzQw6mz5spjGYaGJ07pMRQ4U5/
ksIB4bJRZyBdnKGED/GioO3cMZjjx4ESWOU33T6YnhILGYF/j3VYwSPoRgvQ/QuASi8NiflCPJhc
FeFWh9OgSujgFM0gSYpfdOAghK9NMg0gt8m3QVyhH7IMgN1cdLDlhytvShrkOD7D4J75WWj7wq37
KsxdxSGGRTsK/Tjxu/1pllwNoX9RuC1BiRlGPxL+Cv6X4BcOzPxdrYouh7IPYC8uJBDukILCeklR
TD3B8+WvkR4YPowiDHFDtTlQggssugGnr4LMvG3Fzee4kol8L6qxmc7OKLg/mS2HuzTq6uW3Z2+O
ohaWxljW0urGT4uEk7q/eq5P3Fuop58y83LXT+jl9hY+T5wd938sUCM40Q+Y1EQMO7akJIDu8war
DQ6KJ3alaP7M0xn1Oes+H+BVGxlWbPO/BL02HS9odrBALbe29x6+Pt2lGnxwQrCa9r+OJ8sI5uCN
DyGb85hkLzM7SHkz4JF628ZJIda0dImyBHZXae9s2r8WGEfgTCbVr51YbFKjsDkAIkXXNxCPZHes
R/tzqLXoIi6QbACu/LfQOTh7KYT8E2ci5cCyP6+v2l0hfM8fc0mAU6vA4/ORKQtSpU7ruLKBgNP8
PvtDKF+UMKEprlAIxkv9Hj2Zrs+JNR/yV1GELsc3i2VdNzya/OEi8aYgfMVWn3TJDa/WkPx5FzRq
kogfbWxSlyeNBiOaiv0dFBDVGomUhoR8b9BlHtTaz/m+vgoXmjByB6/0h3qT/5qgYODa2lY07cfu
RJVydRB6OriRUZ5oOfoTGXolBQ9JVh31+TAWrVDcms62LbpFvk6Yu575xVioB4Z978KGt1KB8u5P
8ox7R7Zz+jd+4snaIHhdEV4VUBketxJrcj/AD3MO9m/wmcA+3MjbKL940aq8Q10X2fNwSK6FX/o5
MKOoQGqcSNa0UlGuvNk6ud+cgUn6DQ5ZLaigi3cvlYXDPkzePWzjHPbk9AZkX0NPb+NicaaWCkxt
CiWqdrLFn2+p2tzgafC4Ct+110VSV+V7OxdaXX8B9bHb5CmK0hQbc2oQyaK3zne+sHPD6xSmR31t
JKLtMz/0viGD8CnU/EW57IxXlrDmZe5GnlLdkEx3bwnJhK+TRGdarJU6j4pkMwMs45Fjs4950fTm
1lWETvtfZCmVQUxHE2pnc0nRmhRWzutWu8NYfqqU9h9SM9udCjbGct/Vm+4AoGhvlHk8GlWtie1M
fgnDSr0UOJrO9W962VGD/sbufIcvI3iYJgxUeMwbDvKYcJ2TqFOYce6NZbMnCpqwzSi3okr52P/a
CIOKQCjYc0/gT1pH3nH4quwyM8g8XOgSPTkN3e7di3TaNiMcqRrEIIGWElj6CJXUGA2cNmf//nJL
ze6JbcPSEptwyiF2MxwgHon1h4zNR0Jo+SWtmuM96CxsXxjfpwogbjSeH9oQTeQ8tJBlm34/Etoh
Xoae1l99p4cc1nRnhE8pgUhYgm/A6mPe+KsGiXiLfRdjzgACUmSS+ca1RSwF+og0AugsB9GDz5su
ASFWMBBlDhtFFKNZERDWp3nh82e6aO+scs9UH/S8BDqXMSXRyW3UyBQqTgT1a4PJKegSw665/rVU
QdUz7IbCi9MT7Cv3JvrDl2/+f7T+DwFTbr2oOgM7sIyh5RoH24wniaFHlzntUYh5Pa6LlbOfTdrd
D0rLIqdDRQmz/Z6O1MDZ2F31KfnC6AWC11c66+ACSxqDj6wGWbcPGFFjTmcIQanvDN8NOwR/9UVj
Z8+rSmT+pVjIJPlTw6K38Pm68AC9Lcnzm/szeDPWhW+HPvmK2PSR9XXp2YX/sYwnAJikfvqiSj05
3jxWXCeMKBIr6UiCrkWhyj5PiSTBDblc8816bc3GXXgZGD/uQLFlLxQmyH5LVjCf4zT+H6nUu4np
BfUOCGqGSh0qRQq8mGusdosrKayBNxmdYczZisXlHigvNw2K454jbUsHG3IRX32EOsEs0H7zmz0W
c89xTDhYVvfWwg/kSKiwWj/yki13PNCgJjp1pFXcdGdxZ7T/PdO7mp7H+d48jM7t5L0k3VT17Fo1
zwUy/OT1VKQUFknKLsOF8wHKZwxskDr593CzURUyrg2/6wO/rloYhdnqNHVWbQriqKl5ecqFqmrl
OzvimvJArvMZM70PXT6L9LOXEmAp9ZzkegobtWdTXU4XKgFvA2hMyicUUvZidbg4imw9lGL6fWgb
mh821y6WgcRIn6MG5WvZGBnbMdeaRRs+TTjWXDTMmd8KwBeIrP5BfcqwKGtMrmo0UNOjtLxG+DNk
mQVasK0lKuF2K8GS0D6k6/I/5BpLBhgP7UiZ3f7QtbGRcgj4uLdsi0n/9hwfR93XKOkr9QHi+TBq
LW2KBIlUYOcaHEGl/LAFlpuVgTh6G1nXHGw7MDdYxFNO3Ic1PnjoYKdFEZ6WIg7H97iDM2dqomKz
BWcx+V4MEX7qL5Vv5BP4N+M6ktFw4r4/5LakHUmhP+JNAfjaEo4tiid+ZYw2A9mBjHagarzadXDp
9AuvNos6oEWMVw0QLOdC0+bQbVwQhJkc/QgkB/kdG/Wr0zijGKloLGNi3fLs16iGR9WRrbOe0mYE
iMxpJBhop+c8RtvUyCTjFNnKmTORhhn8Dj3i5m4xovpNjiTGsYWtdsSZ3QhSvjerBS6vMSJ6nLbz
6UIwxhRe1hO8mA6xvgpPEda4QXVl9KXnACdodIxDCapR34Bm0MtMgyY2nIShbXvdvqGpyUCckZw/
+hgiYdv46nXkcz81i4xLkZuagZSycoT+ByBYf8KiGCNEQg7cr4lxPs/G3TtnMAH55aAUYSVwSPel
aV3rpl0jBMBw4u4MxRW6/W0xU+PEkeJ7htrfalKM7xS3cKWfWX0drfNykcutx2swflIBJwyhpqYn
UktP44GKH9ldHxhvneZnjEY3F0W4DG83D8BdqtR1TaCvA9hNNo9/0LNfuFC81KNL8SpQUHw+9ZiS
uDdJT2FBxpTWN+uPQlASgCtaGC4Canw/46QV5TD2IAvJiKqoY1nsUPKJPhrO+JVVI+8/8c6ksOl/
vabyrvTHw3pq2eQ4eseseo3IurQDp4+EeS7WW2dAkdspufdxE4WoobURw87VZAvOjpRZ7bGvatMX
GWfLcZJ9v5ie1EEZrayo0VrFDfpoSKs+dxOH2jKF29Xf/zSsqOFBMXOEA05huIoHTfnL4n3MQPUK
ynEgTtHN4c4Bxh98dbtM2kV+sbzNeVosdQSa3LiDoxfvLAm5/MfCZIOxT1bp+4LVrRDd/GJwQcR7
k8i/Tbf/9nCDvcTQw33SkFWh5gpjyliC1+spktxqCVTZ7el0UZQn/aNW+AGy9ebTy067tszI4xz/
CsnNesZCk7jsFlCjm6RHT/mjUPzjf5yoTNmk54tXDthDxUTa+RFg4JZDIIgNbz6D0vzkA+Sl/Bm8
ovcyBTiTe2bWXGZOtVZTCLXH4KpDlHgwGnZ5LokBKWzl5uW8g8+6x1RcLBIaeZwjXJN3xO8YNLdH
ulalc1pPs/ht9cllPCefX2+f0GSheI8MID3+pzvHH7CaTcsUTQVJBV7D1GAEiCvmHm04PRZwjydq
B+G2LWMdfucfIBjzaCOmB/sKYlka3OWxdKc63gree3esH1uN41Ylt7XK4kWOspqJTwAPiKQzmq/B
uJwekmTagvGiTDRXeKW9igjZfvQtgQfsiDEHEE8NZz5X9xU8xIVDj8DK1OhYx4u7PlTEjtIJbfj/
atqyQKhl0cT2NLPRJSztjBd7Co6JsHmQKNoKVC+XQXDObBf3DSHjiATPQBNtxyRANyGndxpHpI6U
4L6ryXQyHLf/4bHnyccQw+r7K0keUF9iHapQ3mkDlgV39m2iXZ/OC1rGdBHyGuwzT/ivzqEHbj2n
8zIeYn5nM1U8k0sPYTfpzLovmt0UAXp2cXmv5TT77d1pZ3GYB4cQNWqZGFyioPKGY3G7M8y8J+9Y
6XELXC1jaj20pr9sWpRVLzD0S3PRffYlTlxdJcgW5G3iYCW5aOzu2j9fWczKiQQdDG+3TM6XDRdx
6SCO25luqEoWWIboaHSBqoYWDhG67cY191MywEtDn54Lqo+2R0WQzjhLvAefjfDfWhKU636nT0Za
1ec4f+43Ovln+mHvRzRZUHydCK2urWe62aI09Zz8+6eKyJzQgkvGYQ0liMF7cwI4Kpws1JiNO/Hm
/LCnviP74T5K9wQP4mfot5wafLVzEZDgXYFboKDWZx8GjZHBpSqs8cCLQPGFfCo+NPHsds+nNRuL
3F6OThBDbT029RBz+d1Mvds57B7khiEMRw5updxef3mpOZ7vweVDv/5DYXzS7bQJpgYu/4LD1JI4
c/PlhjaexqiQ3ScR31xv3/7w2q31t4jkng3ca0cK8LaWpkHgMxBvHQ98dB0CcssXCzKwZWDe6xxF
SJSM+Mw2wTBNRKUoRevb/L7K6AWZXNKA09Gsi6YjHDrSzVCUhS2VJ9pUoUh1YWF9iaRHTOcYg8sk
k4NTs17r5gXrZPCDbmlL1lDC280DS1ElW5y3vfGaFc8GqN1bT65mEfF2u/XfR+AjxHABxfk6KZ0d
BlZ2BgE06FSJR1ApA6yhtOS5DbfkkgIAAQO0xPqgOXr1dIBp2uzn3o4uqk3ipmz1N1KTB5fc+bUo
1yUW/dzTzjaZkJS9beasnN432wa6DQAsVRSAyfSR4tTeSIzysoNduYyDiRU54lgyW7+Q6eu3SSCR
SKBT07/KOgNl3VI3cESCfn4TfH+pD6CS03nReBtMX6V9mxP9oNuM3gheMeTtWbDR8pXnYLL6ImkC
xWk/qElUVbtMMOQzDFrMSRJzzdSPJTbKxrJcC4Z15NFzP7SQcXiukELDPATQNRS65voNobW4TjB4
teL6lnq7Jpxbeiya5EVPplhVXSwTY0ogdkb2LmEXSeMh0D2k3rU8VzGluwxuwnQBVJtAIyzBsC3B
sJSsiGWuq2UKhOJrXpZnujAnxEc6jm3CBv7cu2HyYHhQilduFzUK6emNmsr46Smt9tjhQyuJFjch
2dWklsG9/cRs2eSmSDmygy+irtrxdv6Q6PAxoIWBNfr4REPEgM8a8JP6raqXHMvmgH9FBbZSEmik
QQQs2WFpT8kznbGe7+o77EAgjd9v4edLy03xko/0x+7saB4MGDtUyjEiic0t7D6HvbApmEtUv7J3
M6xfbbCqgTJSQNybyPpusKKxpLn2IkmQKdzFdDextQm4uqS6Ogn1yvPxyoBAafEpTyY1+a+2/WxE
9xaVmLpEuOyWst0BEaa8eEcT6WcD6rIra9iYG1KfG5856c4a5LxbiYAqyRR+FSd+gQcCBebVjeso
Hzvy6HdqLtY2MjASlfEGlh8nWooZFfA7DpLxdJgYJb+x0pP35sYYSnLlj+2BQ0tL+hXjBLwyVO9e
A8Z0xfDC1GduCDlnIL8ArA2r80DY5KO2dOGPKGt4X4RR8vcROdvS5eZzhtD+RoBXWfRRlWYpjzPF
xLULTwFpQzvofDooQA64I+h7nCDETZt3rYHCC/vAzEMXTuVEICixMONmCJZVKtgP9wiXeDOLkS7A
V7JUBnJjWn/B1tPmmM/yUwiUq0Q6kv6BxjgeBILExfQBwy8QE5+esith/7pmngNOG7R0brKNXSll
yB84Ed5jJh8wiW/Xmqn4oNnSem/S9KqO1h00jAiJ2ousQnj6fRt2ewB418MKniv/NRNR0kziNlLS
xvbz02SXqMpc7p0NPtvWzYIuhKXdGSEPsfb9I6DynOZgN0+Wgm+gS/WCQbDL5t+8hVQU8DEN7Q0X
b7v7grhvkt35M/o8NjyIdcrm6utIphJCa9xgUyE8aoICdnsxN6/yx/mpmNorVtTzz4gOk40mEpRt
/V87CfC4BE6ztMdHmbyqNmeoCxjdB+k5bdce/xqc609Iw1UwRP63TD0h8pWvc6WNcCKCLDSN816y
LAMjiNxoEn2m8redVHsW8ajDdzD0e/xNl94R0xsQfnyUSqAyWL92YHgXaVVfr9pfeUC9Ha/JqWFb
RFbhUHb2JK+Wm28j/Mnth21x/1/6AkpaY9h05CXt4IWPpLm+hLvsZy5iBocUHM8wejqQ95FxSnJ/
QRhi00IVUV45CYtW5lzpZzO1zdEjDeTS2IkG0QCCZM689rnUCJzcA8WvgVQnQaeqrXTXdM67lETZ
wTs9se08oPLKAmeYi+OvpZURuqkNH4HNIglvY5eJ2QoCRIW8lapF1OkblQEzSOYwASmzyoYrjPWM
tankVR7GGns2e8lngfevFfVL9oDb5liVghv8KcPrqM2K0JmMn3PeGmanO++ErEpxP48fP4Or9CSQ
z0aYOJPOX3uctzfhhUegbD5ngtq2szSuQgFmM+vtJRMylFwu8jwZvzXFst8lFK69Ywln3HsGfb6I
fKwrVux298AaGHnTqL2pwo6EDsHfHx5HH04PteBsisZFIEQT8g4uEMZRqfChhgnlulKYG/2tEVt9
2qoHrC7m+iYN3m6hNTgHon38BGq78MK+v5QL15Ny3wZ9Q3eI9CL5snhe9byf8hvd8svEfHFcgdWK
Fb8SVgTQ9HiSnPPc8/bFi6HLszcN8FGvXg0XHp/emNq50TCt3jn1hRi1ZWrVYJcahS023IPmYEfA
glomxZdK/ZYAE/ilNcVjs+JtKxOqn5S//kRXY0eGf0efyQQDpQ/uywdBgvj/p7fRx2sHAAit/w84
IV9ZeFPioaSdNsWzF8WBclUz5yZ0EOKFNRFdNKe98Vp+4ae8jwiwWQ1yu9//1JCFNDIqtChYkcGx
x/4k/V/rElLq5TWau2iAGgCxwFvlTB5CnqdDS3xW5EywPlXKfcQTrTpGnYXMCOf5kbrMGgtJR6jF
HYAtjaSOYoiyc39B0+CbICvEWy225jhW/L7KCAJ4WdIar4sKxepE03slEuVG6AN3N5fggBnBEm40
XvCwpUEBAoP8Yjmz4RbX3O2EmlYpgZIAPx/Ce9yRSdgLB20wP8pJZy06Nib0WIi9fEc/gQk6yBMu
Q/o1jJvGFWH7xhqINHybTgl30Rt8Tcki8o9Ozv+h6GFPxpHTxiYy0jQJooL/hNQUYLN2GPaypp9o
kHY8bJpEOeiWOp8nhd948EoRpwenebkhmdQ5l2+pyibWSGuijE7CoOKXwDHVDee0iY5pxA7wfmwQ
qBWiOGLpIy7J3/qBQIQYvCjhK8srAb4pxIhxNB5bjANDbJiVa5pZhOlcvD8k+n4vwtJkcyDVoxLs
EhfShYSHDBk2Gz44pq7QhAXC9pd0R81vu2YqC7GEF8SGa36CKQXmxCjlkKEfsPlbVAJczqG8st3N
6vV/7VQCa9ghZKdx6QMyIBxah4Zxf6NqR9el+CBi+kRI2OV4eEVRts78wv+1wxO0diD/snBIRCO1
zra+x34F0DdGbYYp59E+U13YK7Bsp5xEbHAqcmZ7vOzY3vvl2iSOCB5Hfe2aFkjCsIJ2HGe//cXW
KHdNPYpTEj9XF4ifVATfv/b7FN4ibACXli+fzGwBCLRrpc+Ie74L2BhI9ghGWzJxad0GE2ZFKoBB
7mT5+veVEFv91V7vWKR4nPiLoXhliOeGzwBwTl7BxJnQrnE9c7G7+t9mgYDMLRvIicBgpQxJaN0i
/iewwRVkvqbmck3kD9qqBDtrA1jyvT60pq3AJVxUCkePQZ0Ak8wr53qLeGChrEeSDzRpEbhB0cnG
rJvdjdNDKoAdwB6b8snBrtb5gk5/kDHIXBiE1WKTTA71IUGs0u8srD9JaJjBadEku3d2zYQR1ddJ
gUARppFRxVAUZzng+GY70t8gMXGUVrZm3X8eHnlmQ24GH+e6ZdSfmrNhQYbLiuyLccDw6gWHFaM3
IzzQJE4JnsPncvhjeKn7M45WCCBE0cDTcRDx7m4CJf+EqnlOjmWj4ftxXTf3Jr0R69rrk6lDOrTm
+XdgYoff97J+Ulgp1FxR3BNKYwtqU8sjRNkevey3tzfjyhavFUTR73c5Aqln72LQNzkGHcDHdCcY
b5n9iu0k04S8OgIuZAVn58sNeLGrC+XsR6xpf9KknpvDicevZ6WwlXAZnr5PleMiPCviRev7Pcdm
uEYQjsrHGb/3NyE8AK/meSUig/4i4qSYS+1XI7JsjmaxIVMEouNBazXaVZ+FzmYxhOJLKaOMpfbK
xFP6Pyp7Ktg2PndwMGymuVpmPM3lFC6qidDoDXGnwDDU3SgzPUlr3eMsnx6MdxEGZcaw5GyEGaH0
/1ZpJkCsKJnK04FiWs5s7UNoJ8M2pxpQO7neR5T+2Nr+kIEttmUMwaxpIH8I0ePANcyEAtz8l0T2
fHC1NhPkjMxf2SrKk/JvczI9p5NcIRWR3IdsM8etwkp1II/+owZbGnxhOC57DCVYNCDYnir8xGEC
keZoliUjBBhp8bRuDrbbKIyxTnInRpHJDjrgh0Q3H7VTlSdJ6FEqGaif9np6tTgnM7qjhSTQJmSt
yh+aK39ccdYVQWEc5mESde8ccXIjhKUdWZBCEt6n+cBGchLEIvgtU7B5LPZW+3VvcoHH5ZCt/h/N
B1N4RH6JfH5UqVXkd9cCpcQmHeeGWZ97uV8eXHJV+tRGaLd4eESx7wl7WZkIkyTutHGmG9o0dhn/
U6lC4oIkO3AzswQpF+WAtoisyEQdiivRfPx5Ja7h0zguT3fF3X3VD3uIJKx82tcfZsPuUU65Gt/z
zWyzUuN3dFcmR3shvHdRlczI3vJ/14QNPfHn2gy52XfEZzs5RC4GYnROkPoWhHzYGFdIsXP5Es6L
8oFCaZMs0no0TQPmlmpOJt2iwwrHjqjoB1M30J5Rzlcb7ly8d7JpVO3H8l0Mn03Eo1MZUEgL5hVc
IRUZSDiT7JjU2HmxxTRoLcQ/IwQ3gz2n6kV3IgX3ahUZwE1P6d053o88PCtI3rKVR97dZGxYEFsM
plp+pimAaVInjVJXaO1IfmYHd95wccKUkSDoLENSlHZvyJsk3+PsYZiS2nsLE2YFsGff+P7NOOq2
loQqAwnGaHpJkClXiunUA4jOpgMqG6N9pvwQ+kNxW3h/8txr75e+wW5H6i/ROvne3cPIqOfLQK0y
7mUXsF/M15Mo4G158DZlKXF0O4PUP4/iXzK5/R2jCtvDQRiYKSZ2rF/WP/FV+2uWIijx+7cKQZKp
eC+jyJJneJguptQpqvolwCVszuNV6T7oOVny+xBsACKTS47u2mScTHJNdUUaOoAzQz4cein9nZTy
T7QNaaOfI7V38YO6jgXjkWJRWJRO4Rpm3pnVkdiQD68d90qBfzYrhL8Fd/fdbmXw10r6iyOPUVOR
iCkq8fzE1zT6Ge76Wlm/Iw+rKPM4e/Dpq26XTHx7Kak4iBfQ3paljPSY7YLgcIanPMbPKeHzHnz4
pR7uI2kpionlDNZZ/AIQZMmlc2Eh8/fTgrLllyYZgF5xk0VuRHsCg5x/pB29HaOUEmReskIfHktF
NM1bh9huAyNCNYKk//TI8+LF/130VVBeMo9COZumsTTmrt/tZ+9kmJvXtEiBpP1ziv5gw38xgbFf
ozZ4JMpU9biwA17/vkTKBgshWs8Lhe8DQ6QvqCrnstXEGXND0rihNNLFkVgMWVg9xRsQmq0FY6Q2
x8w/ttGcIhHj63Xr/2LkJeK1e0XBPKOCMMN3t/5XyVIZj9ZiMYiJKgOYNSGtQ55e/eSSv7+QKTIq
dBN0ObJSi/24MdMESToz/HYQwtNDxgcR5DYjd6wyxbqfryf7T/Lb0LSz/WQgogcBZ2XUoln8caP+
ecFZ5YsfaqlyYGCzif3Mm6xfkFlPN+8Plhz9NMGd2aDUqiibfFrJeA6g1rMQqV3sKVm/NhaLF5fq
u0yaHWWwjhPseIalVfPTbewgMzUowlt87Du3Qeti7vjtFTx3TSIvDxcPqCcbdzQU7i4RoYvOuZIK
Wj8UgaoB1GRSc8UCxYdoctxiKB4lVrtD09Tj6PeIq4DskPpa7rVptcNBWHzKFG2CWC4I7VZgmqCU
aq0pJQwgJIMH0Dg9JSJlooTvpaYaKz+QrKQ+bOMLePZbF8PKg8tw290elXuCH1GYEhoExsxNQ+Oy
H6Qw6bcEp5ATgmqpOrwCMOpb3RDJvBn7LW7mAlePHEcYdCBlPLzrL9X50kSjLq/VinFlUTpUpu+g
tCvrHYpruiIrdtxSO2M4UTxJCAynb7Jlzntjt8ICVmL67vtWqjyYxzgncdH53Q5fXxSzi+c5vChe
Uk0IqH5R7FbB+9pg1nR8rOerM2LtfVY3ZAOHNhvbyqwBfSqy/gw+4iLZKqaCrojKb2C0BdGnqrRj
JIt2js1LHsurMvEvDg/cApSITBZguE9gvzNcEJK0QHKju8Sh30J5swZhEmwonVJ+dxRH2/vKt2l+
K4GFxvVrw3HmXdnpseTaT9fzETKDA38M0gz4Kw5/ftOwnl50bXXD/REcAKdCQz0f9lbXefEIyv4G
63LIlNBlP6z6R4Bb8LirHGTwVdqgfKz5j3GrrhzYrd/FssfpCvRg6gmF2wlAgPDtg0ogFXQxoe0G
SH+FhJJGy3wh+qYq3cuKhkkzs+Nv0LHx7BK/U3tFLTu8AUVtVc8XFVjsvJtLJ8VArXDJRqmMBrD3
SHLRe3yKrLLaL49IcpOCd6yOAv2T4hvaz77kemEyZBWv//wmjni4H6/wln7imnOTmicySVQ8uVEu
jGgBhcm3MzihP6lTagBxPBCRKwG8mCeLMpu5aStRjuK32CjFkPXNL6qvCtsZRj63tYU5KjIu/WCz
CQfy/n44r8ua3N5Qv5IFKf3aJM29ZCxc6if8OygS41vHELHVU8vX9xchZltic5DY6iam6EofJQO8
yeQTD1dkBlUDZanj0o2EIRC8DdSz6Kb/STTyLmO1JHLig1BpMaZ2P+w5pujZC9YeMEnHnxc8iBn1
0wczcluSk5ql+XMtU/v6GxU07vjQub3ZgBNs6DU2Ch29hCG74qlepIDLuhLPLAOzoa+OY2ZJ20T0
B7FLK5Zr3z54kY4BV2M5Onf1/3IMOnIFmRI2pUZMmDFATVKtL9f80Mv47mhoI8tYXawOVE7oG7E7
4r9xkZyTNtySSoNXZmL4CANQnoNMXlVlC3NjdhEja/4TND0TGd7YDKJkgHFQRAOIbVoKqcQULgBt
xIOM5KFHKdQy7qr4pAXx+M5yUubAwn0d5vqA7CgDybO1IfAIOeh7gLnvPi7OxcLpYuoYk53UdHt5
jTfR62yV/LPuvd/peXh35d6lhFDH/pyYhrxHF0fq//Igeiit6XGCgzm2B1RPXHksFE/CvmEVA3gj
QxlYbqrJfirhmOCr32pWXngB+4xCVYnLx4rn6h/mMKUmrHAqUSuAmQgqSIYHfisdE4meXQ5W+cN8
n6Ljg88zTilphcLM0IOOawJZicPOD6KQUVpLWR2FDPbEwBzlo4ZCv2VMkIC1mPFh+GiBcOzB5yXy
bLXoioFr2KoRh2k+v3k7N7oReUq5io6zoCAq/+weYNQ7lAeL4R6J2N4f3S4PEK173x5QhID0PSmp
Ih1huVOgicySma/S6TifCJXThI3d/p2skxSHPIliCQhEHm5tHiNciUWB2YuThH11QuRxR4EHgwVM
gG+BddOEcA/BhJEYQPEPVEeBTPOoLRRxCSge7iz+S396r27nynes608/U/HRQvTWqc6O6vxI1f6f
W0q9Q6QSHsp6i/c1JdoD3aCbYTCtECHjUxZbd03SvvYNzMJec3Xez0MPd219n/7eLJhYdjNcUX7Y
4jtZe+5aXk/DBgs6vYLV8QhNs3cfWec2ffmJnWXnGaZREi6p1xv8Xn2SdQC7Nw/t9oEnSxbwN0Jg
05Kwctah4zEpfqhCOME4xMgUZ/RGy4YnRKdf20M/rzTO5rXj0iPhAWAAL5zO4cIIPFd2WfnW0SdY
QunTASEYYNJjpZDTXM+FVfrxnucNfuoioDapBR7wmHWBc8NvnudJNxCREuN08gSKEQ8eeMj9ZmtS
dy+k+r5+P3zl3IbYCuwAzxs3LvAtdbBo34GTp9j0YEcF8h6q2VID9sc4KyW5u1XmAJnuidpTptbo
nEtaH7o7JGiwApwsJi3k1HN3idV+4bnsGlW6NvUHq7thdt5vFDU4LPuTDbcGGKKw4RCmf68whJN7
r0usfgFzVIM5La3pQJbru3F21zm6FMmsEiHBfPZbG8zr3zfNBd+RJtwjmnzxwcGcYlKL90REoMJX
N7PKPNciXAOskA0dh53+BZk0djmJbdICpGHKhRmD4E+TD1K46o0MrM8evNfA6Zs+4TMdK00vBmQi
2PUTXfsR2gngGNJ2wRkIXxRmBgHHXrvjA9aZK9R4OIYbCOM8k/K3J7rVmwgDi5WLBfQpJpEP/7To
DXYWLTxH1MpSIlvalUDc9MhR6X0asHMfnlHI7R4vF4SW5riUuE1Ia4xB9/56VFoMn2M+4QBjPPt8
Brrg8IdPCQCKB28JBkmuhPqhRKkYTlmF7XrmVq0i2kkS8F9w3+QG2sGj726nZ3nFbbc5kZ68ibNr
D7t6j8OAxlIYWcH1m9N/2jEBfuzaaJX60k4xqtwoMBArISx/rPdg4eHGl58rDiSbzR0rnsw4DkW4
r01CjNCo+3hEVQ6CzlAdPCNQi7RZOAzAXlFjkryuLK3xMAa+1FJ6JkVMxq0HHNRL9oGLXoQa8n9X
dIVwTGBl6PWLl5rScxbZtv8aNqOYz/Evt6nK4ALfmKaQEBFfflUpLYce7GJ+LyrG0D5rPy3V3iQB
+31AUIaV7/vtA8H4eekTNA+tE1zuDDV4SIPqroGnr1WSSZPy4hPlzr3inoMAMi0zurxq022JiUpJ
UVqUMf9Yv9aXt/btm8LDadOni7xELI4pMkxClNjDgfu+wNyBpdGTDJ6l2RlPGBd/fO36r5W7p/ZX
LZVeOI4S5tn20mPtjWbOkGUnMwBr6AMQ0gYChRW9LVHV53pN4brxtZ8Wtrk2gyfMUxdvPyVsuZ7e
c2Hja/IqQ4jfOVffpC5+r4ll7Nwiuw0v3F1Y+bjYaMKdMYhPKxyjq3GfzWD7cAk+xfXTYEnJedCU
Y1usM9qeE6RlET3pc+q1/Ft3Bg+0YjS4nnc6EqNdn5IGWdb8ce4QYx5DE6BfY1td6Ojsy7V80rgN
+u6gG2rf51Ky77K0nsaMr6TwzpXQbf86lT46mBMhE72vp+/mpjJYSfOwz6Oiaio/DVbjL+Zj1VaT
yRRTw/iNh5qw6szl3pgNKomLX8lTpZBb0A+rIB7strj1AzzpIqHanMHM9S9ZstzMXEI5izKpHZ7Q
MTxXUDwWfuwS7sRhBW3OHpNDXRPElkiBN8KRx1DiTCtnW8ztWESaG3Ef9DjyeYzZHg8OLHUwYHhe
U2+18ieAyK/8dV85r2bmy4vLI9r+WMTl+1dGwGvxrVzmYp+YUs0ox8FkZktvcJ6D/6i7eDuCLZnA
DQbXQ9NC1KNYEoiRHs+Hmo4jxb/OAO4FLBlZGTl2rja7rafZwz25OVCHhYKPgNeL+LF2eqWgJc4i
4r2jEOdvrdCLHrCV8WPEDR/6DBlXrmBJpvJ+4WO9H2DlY73uOX6uwUMWdy5tGkLxxiWahiaPco2S
O3NZh6dfDsC40WG6jf//1Cv5SxBSJDLa3RxfKK79mSJCFmySA/6dY1t5YGc8YLyzdmwMPUeecBnj
EvTmANofQZqMgUYEjPCw5flgrIiEZOCVUw08wzQ3KgkWdi4MDBnR84+HrGRW4clyyX+yiDZThUpI
j7U7VQDdkUIBkrgeIxh4gVio0v86/ZV85tYdOjU32MXApw1EM90xTtS2JLt33jTcRd6WRLMe2M28
FSnLh8ebGnjnD1vdw92jYG4TUdk2OgE6Ta6DiRUAompfINh2IpRck8hcUawudZ1GCn3LU3oGnBFq
bNC/3LEs52s3lT+JjRzXIZGXgO0A0dwwrVVtwLZ1xeRsUojx2dZGJPiPtxZ0n5oadU2ArXrlKd7y
+Zf0PDxL6Ss+HnXYjBgliHvo4oZ7VOeYVY7HqEIu6QbknQOoiu9aQMdmRuZcUxc2aOh+1fomT5Rs
ae1nRQr6220/aPc1LmWuD1RkZ+NPt8V1Er40AGDS4dUnaVgb5oOt1BgQHCnESjdzwJpspUCi953F
ObArUyrtc38hYp2yJKBwytgrIItBF1UkIdGeIDqen3SoaIUrMNdGM65NBAZ/874T9ES4yLJlhhuw
KCE/lBRPXlzYzxOPiDmpG4iAo5xQ0EPcCACz3t5kOKVUHRd2DKOLvm4H8AVqIVg4Jbo95Yqm905e
VkVSDRdLDS57Y2t3S9CufduS/Uzj95f7PDR2v5gA9LLgPy2+9pwpWMltcfNQQbmhe06rLqkrO2t8
WGo/ltVzwRIBoF5Vs3ZfrdympcVDXsN+crS1ksqX3ooCscjkaHugZZ5heJCvDgUAug6nhoe5yHJm
bv08BW5iuEKVQeT+BijdSIWMstS4uW7WiQs4ZCSUK35oWWMV45vUekKw5adR/wlq/ml4J3xiwcrK
MtgpOxlF2KwMMNKaZbz8fYUJWi6ioI8jRSIKVNsYGmHBVvt3ab1zrfINbtlgNlStRa2hrHNfclx7
tlPZIV7nS+tbCsWGBELCgUL3OCySotcJjkvy+oaMaWuhFrMXemQRmp0jsYdNSGOF+MMA3tzv2l5R
kX5OAoArx9q1JZBxUBwBraXPLNVc/nLqq7izWuJd9FoJeKB5wws4xVcucHRswuWtLIF7P9QqG4r3
8F86ydc7/lvTiqy+pXtghNhtSUR8AxHvjrHMqVkw+iS0payP8z1GlCpCULOqWesJVGmGvknRMID9
ugIKdT0dcTO6z2BLhF3C7ojcbwW+hh+zraH6n/JBE8F2+MwHxgAF3xe6ngkY1NpV/I5G120yuP7H
FtU7vnJwB9txDVW3xSYwmtpLP04STVkg5BPQni6RdB7mgtqiOce+UMlVjDodvcgKRXyHnMIqfgiM
4q9EmAm6yxNB7pQ4mLP9ARryCodPQJOQNQeH19wlOIikw7/QqMsmIjpY23WskeYd6dl7xaVM6wET
/EIoJX4nrr9ujhuGVXmmTSQby1CXv8s+Kp1g3bCbqJaNjxLrye1WK+63tU/OMz7wsj73nd1HEamq
dFD6q2owthkUHlsziodo3YS3pGi1D9s434I5piSOGWoLgccPVj/F0qiSABaz+eTR6gpVX5F7+2xn
efNvHcVXmYJ/SnMt4lVtMuxGtV0RL0tWlDpIfO/JzMPihA9zMbP6pczXFp3E/Qs1ypbs9kjPvKGq
hxGUe95B/+b3jmF+jg6U0ozg54DF14dMaEkK01dmRjnprRiQJbSgYCB+zsxkbZAD7ad+40eAHW1F
08khf0akvCJ8T2RK1/uyXBVgdDTVxNlMLIJOlOfKr+c50GblH7w2XxI6wsT8WBxYlc5YJws0mTIH
f6BsLQaeipr2C1bl/mfKskzrzq6iLgobTupOIgAvcMlYucE+f5UGsROvr+FBTzUACvK9JfVLVRXx
E+0LjXQoTOzb1h1TqfTYkH2lp4A4Gx9ldUbw/CyFdu1vrpCF6GXqo4wAPKY/L8EmlmskytMj5dAf
tdYhM4sRL9rMq38ywXHP+fZfr3wt1R4cEbbklNdRFDwF4+FXoPu+MfSZYXeThGDs9Oq1HcVbGYSM
xUwIYQAhImjCYftVPCXzsOtaNYovWYXShDY2s/+jR3qpfVAKrFsjJeY17r1BeTs+mWUlHEZH57x1
csIVJ5SXN5sgReQu7TfBRbpqCiQS0PIKKHL5+3t+oVQApCjtzegBI6Px+EuK8wYEnXpr1+qtwY2C
x9+o0leysmuw9DZOoGqk8CEFhmSLlOVOrVvvb7+3dClvYcCMKWYWbaLg8fnDsmRHrynTgDqOgzU8
g8fuWc3oxQ2j/b/cuFuW7xvKXQZRpX6ZhLXEeWjXmqyHkocBaeKAoOpgMqEIdE27Fkl+DFw4lAsM
LELET97EfXEYbKE/kkxfrqRiX5azplqVgQLmwzZZE8Y0HxlHOi1t3QaVf3ZrZ1T9a7BLKJ+pJSgo
yfJ1IWIKs0ZQqM+aYUBtezUUBgIDEtaS4h5QE0aSYADv5lcFVsu28ofbI2Bxfuq0o8QeC7l33451
tw0nTub4vHQ78NGtk6hFPSbr3FMpsrq6QCmMZfrgBSEEIvH3+HnsY9MdqafYPMnd3w9yx895ePkK
1aSskfdqywSDpMwUY/16k4Wp0KCZvzqigoQ3EEZfUVveVAzQWVy/YmSJ9WiOS9QYCBFXnhLK0pMz
eBnhTLcI+M7DG7AORcih+hg0gfxGahqFSIKi61sElp1KQQiUNtiaF1uzuO3EPQTavDXg7qPrVthU
vp7iTPb8qP8IAuuZB3KopqJXKer5beTJvIvu8GHNwYwIivTVasz4t/wt8WajVRcX6UsvAbOZZe8k
U3lBKvA7PbsFSDvr5LRCh6ptdsJHzJ8hMMHixPbLNcrQbOYU/8pJS4yp1WvPKGeP7ZBB88fSJ5Kq
OaMbp5W08ly5oGwGuYaBWSnLe2HS7rAkZIa/t80RwkA5V4vms9vUFOovv2+VhGb3dN584cMla0TI
3UdF1YjgN0wO+xH0QcGHv/a8VIAEaqFru1sqc+Pp7E5S6me+fbycu7DrEeImtpRXRIMNEoEZgY+A
Agv9U80UF3MV81jjhEAAqRUKJ8FCvP6xTLsOknWuOKSijnpunA023Ka9cWhgAV28LghPOx7X0pWh
L6q/D2BGhRZuq+XvrJ2wsb9ZmdUsk0h/DbxrBImIIQzdRh6mfxK/VXyIz1L2jbEjIqZ7odCLpHif
m/U5d/8/0QXR8+m0CFCuHTV8y55bLgupFKx4wwL5aYq0yYv4/xpwLZEdTfJmQkbxMrm3JzuZLJrd
o+RxDxX5+b6mgb98S71VKbepwzPxEuMsWd7T146SCQ7z2Mhv8WMAKDDIHZrlCr6KViuwD1eyCKtR
atd1E+ZPPRdmyxQXrwPCctxpxnCP5OLWt/teutoTk6+ZYREgkVVUlIuqyiRe5PQccm14VzHx69XG
I40NxKm4sx6LUXyyAX626gTynq5D7PnbLBvXLqs7eXURYLaiZySSTq+JUp9RsA3QqitBelh0uDXE
cQrFP2ZKtg1FEmyVywFV0jNdT1n656ztBMJ2uQ64YoTXucDv2nfMIYRgNcCFBuMdiLQZPsA9dvo2
0jPKrVFJhloRO0mqXR9gdrN7AcVn60JkfNiBGodA3QkmeEwQV934GAt/9+hGqtn7qe2SyglPa2U6
12AoVBLFj4D9+Cecon4p7dG9fIXLnFk61bmBGE8uuecspXq89JvLeiCBd6RCptSahyIJAmu2MgFb
pyBXwX45rmd8X8JwfsXJYTKWnOfj6FmbVqFd/vPgwiEQ5upZASReTf+bmBAOSwvd1/zhmZOgLYpz
n800inw2rp2Bj1xwgOMsMl+zDvFib1DsjV6hDN80d4r5boAew1MZkSM6/p+WXZ205cAiyTM/KNiv
V0ygeQyu5uL3q91C1Rh2Ip7wpBmKZSWe41rOjmmNyv4xZJIIn5bMn70w+mpJ/1D+l1Bx8Q5Tkab7
jIZA1k0yNpUdx4x0QYp6FnerBEj6HE4nGlgAcFo2AtQ8LpAbBVNDDrf2QIM5OR0tJ6j+cQHA5Fas
nKjkiQhvtdaipQS9kETgxjQrNmmxMmnl6RK18dzv30xfcZllDe4dOQjXVYPrgP8IfXFo/OZDT3Tw
5z7x8TChB+j8TiUxl7F+advTXMPA/UrbkEEBpWhphySTUDmEpd6cMW3JGA18fLhXUPjULXdn5ed9
lmAKWm+GltRyLHc3rQpXyG51cfGcvSNGf+UhJTMja+RRyRSIBznxfDvPSgPIiFjICYsImTsHf5y+
CsLzZA808FjQTM3VDgeV4zSZwrfHpih99RCH7Km/SR4+iXatUvTa979CZWQU4MBWTyN9B+Z+gIMp
zmXWx6PLkEOBrNsc9+CoKPzw4dITtxKIVXidMdBfYHp2qKcqyd9FYq5T9oV2r6stL6anZVlL+KMt
wEn95pE+JuzjW0nWeo7ksXCRzk2TakE54QMZGp+8wcjF/VU88JScPBRtEPpjiy6qRukBVtKrqxRc
mFUx3hSibY0o1AnhcyhvIu9IW4/zBuRJgZdAcBIMOKuKt3yEvm0DgFkNRnz4kG7FjK1S0KQ5nf8N
WBiLS31vHJI2Lym0mSclWmezSs8ExGy+EtX7+RE5GMBYY19GBn6rJpgG8qrnmwQi4ru35diXzJw3
QZSJTCSyfXDJcCAeIM79goxtZEpgvsF7o6GtOGBB6oAHKrvF2KDlJVod9DmG0hbpfUcZViRLaCt3
bMJab20mQBu6Ss/gIInl/rB5hKib7tAQEC2X7kzM1PyJ8jDKIfHeSdAzV3dDNKhTDn32od1AKFSR
imWmLlYueYyVFdNiK9gezqC2Ntmqy29Aoe1gDvyAXu8l4lKboeeXZNVZix5KYV87IJ73ZnRIGe7y
Nk/KkDj0kfE90eaW3kCrTC9sNWfjr7nHHdOqFdgLqyxM2AMuuLjX5JpwxR5NZedKvM7q+jeJaW/p
Qodp22p1UxCi1OJdreIgRUY+Hy7Rl2kfr27vfQtb02C4oZF+L5L4UkmCtg1+4qnfIaNWjXHF2GqB
xwd3G72TTs1RctAPeYF5kJNU/OHtQntemWdaF2RCCg8Q/oYEgr+rY27ha1wSat/klMQL6L3H4emL
RbLTsozbCm5N+P1jrCXt4qwIq81TtsTzEhd7mffUH1GUfngH2mLdvR/7x6n08iOm7BdtvzGg5IkN
HIJhU0w51dpACLBRd/HhF9edpEAwPXvnZvrW9C0aPt6A437Mc04NYtOHBfM/yxdT+bm/6liotnm3
pyGKNC3LNxCqJXZ+GOC7leuudJohmtgBthFMayPGd6auzEtZ3hhNHp9LAx+kD7rXuWGkt/FsE99N
7eJfO7DTnChKRLNJw6cAT88q96IIiOWpZGtRjDbGniY1pWF1mRJF6XFUVt3703iGJ7KXE/Bjsrga
7MDf7ZDmge8R2AwPTO7xVohH9Me767a1ilFbf0BhsbcmseiEFfS5ohF9AY/v7TD7WXi9XRvqCT6V
pxu8DTER/M+d9ZoWgNB2/tXqeqDTEMtGUWh7VUs7pUzeZKpod0VIfCxoYxv2gpiS36LWPNw3xV8D
LkeoAFKAxynno9S9LF8xXPJujsGT84QSMwQU802EmHHnUrgSTDUJzZSJhmAtCAxF4DCdScUHTEK8
c4j1dCsCg+YCzyRp2f8rXFKKUczsYkm1NGNgeZwmTduKvMYI3w5Z0gVxuzAeOxGCSgAUxe4DHOJ9
Gyu++n9AWc32buhhqGU1nU6JUmdaDi4+yvTgTrpm0Mh75b3uJVRluUk7M+zn427MGwwTTiGOXGvz
h+sGFBoO8iBVItgvJJI4t1PrL2xVolo+LH8U21vKRHnaPIu3L/wTOGzUpdfAsc9xnIACjnP5/HCJ
2Y4CfHN4SZJcEpOgunflEan/7SoDpoNXGYNekP3ZiDC7qqnjqwbkh1PAK659cj3+v6qjYxtxgkbn
UjYqj1bBJ+RCphnh5iMWik/q92H7Q2pnn/uzfJlDkJNMi4somuGd8s+vCRE6XvjGvFg//NRf9bff
9HNhluHsAGRoLnNw48yX2nWDoaXuIhKMcUVLtIU/AZYNzeEIZLpK+TGBKfJ1z0Kk28FQPFQRTCON
VddmULgqqKgi9mdz/FrGzxxKCGuW4LXpzpDxsYN3zrWneUNAG2sxPQCyM8tuN6gUSbaEpfS6Fmm8
4aSKp1xbVJk0Jn9Rqob8TLZQKHwL3qOsWvfxLl5+5XUtt6QVo8d+ZH7VNB6hWJHBImtdRauYzerF
KRMQUPKVpAvKGzHPsM8veAXMcqlZzVzkJ26EWO8InqRQ7l8JrEBqtj72i+gloPSH7L7EE112zWCA
F1fuQpkvvD8reWdDfs2gIIhx3jNyTJf/bV8O8lmRg30oOLcMb4WrF7sMLh3/zINwSAkbXGw6RqHo
xNaLq1LE9eg1jqUPXLkNEpl9x8HC6J10BPN1vBKI8QQKPIf5psIf16hkAJr0wN4t6Fhxrce7GC2q
nXDH/vbeItPYYXworQKABB5lTW4lGglAHX8ZqDCy5LtYQtjPmstTsRb9VXf7PK6HeZwHRFKFuCZz
WFbBSF6OWQe93mhUSa/eyFA2+wieHbKYH82RESxEse0FOf8fSNaWidgN5U2LA+HEIIWiS9DJYAdR
BHBqVmfpVi3VmKhPAX8WVTBtqrDsndAkUhQ46BLyDp3ykp0OGaY4TJcIRJ5wc3VhShISzgGd/ONC
KAbVhMcnU2BTVfUbf6p06DKiMnFIlpoO85yHFDLece+2WG0ebN1ei94QChkXmyVIu4F9fwFuTn7h
QmPwuWSoN5EEtE6SZQUGpWC1mwLIhN/hhrrzQzEH4Tr//D5jC9avsgcDBsv24zGvqzk6uMOCl8Kw
U1RuXasSA9WREovgMZfJFik9MfwXVUdWoJeRZPhX1zEVgbrsJ8zPLYaFAA0/QFN1s6olarUXuSD2
9OLe4+0TsDITDHhlsRcfosAoLorUQPS9TL6VrGUjuytFbnmi9KEPDi/4HHcecP74y5tK60TEzDbP
RBd9iudQuK3jNmWfM41w4hx0/yFZrRkEgkfaUZBoCYL1lfiSH60E2+f1zkL/1zdRvdGjQ3ElmizF
7Zb+TNj04qMVSVfzm2cvtexlTtt8OzX/fBsjAMRsBHJYG+/2JG2N85az7vCDB3Ul7h7CBqAJ6BbQ
S8KDPVAEkFGAClAT21GHyoGZ4NKAlhTWH4wtzh0ZnpzpdS6SGJtRA8Mk9SspUKyTV7n1U+PtmAIs
RiMBgvJtCeKWaZHf/eMo8OEr1k/mOaFmCBqkmeFTnsLowJraDRQmUmDj3Hi0QxpTc+a4lz3JAC+p
qYd0a+PogAp52Nv0zIprlQZgc44f9He0Ispmot82lC9ely0oY4zex9P3MCDXwgCb5EimBba8i3ol
0EOOGtoQvT4kjQtP5xfcgtN0Y22RM3PVQO3rdGUTf9MppPrVALneOyO1Lch8JNK+35yU8MUPOYHm
bMks8ny8nqZBYszGMb5aplEJuwqWR4s3GX5yFNRt6fqVqVlkCVuafx1kqR5taE1ihjEYCcZlZjqp
ad/KcppU2oJnQEojXd5HfEzakXqZg7WqZlphsf4BZO4KjJTu9atcnCX7M+kWpJVco1qgQjSSELlH
5m3QagCynFtRLnY49dbins1XQ//xRdOIYMbGdKUFvyNpKqle3kttgtKRHWeXaRkYVaVgWKH2aHnr
qpDm0pQBlXEpNqke/gV3P2bWixLh5aPuGqz5fwtoFwhs9wUINRd2JUAtdgDmgLDwrT2+TkMwC1ZG
+uzeTMVuLpkEJp/+RkErVxnamSWuo1BT7rpDKO4ZktPMT32XnM71DROUJqv4yelgM4nlFDNEnGNx
aHduQ+8MMZ4Iby8NMKQYFATzItBUnr01WdndJ7DC/7QA8gecfdD591/up+4dUtfs/ZsfTfpgmGrJ
Jvrs64dkI7Otfjs8dUKjUdb5HIrYWyNiuRQXlwoCwJbdG8ifLYedN6NqH3Nmv7czYRA0LlXJb6ZO
W0yUJ2eKmsohtG5b0U34k7quPPMpmdisihYsWEEJufOH9rPeISVh8sLgrRSxdg5FV9IHq8J4+hpG
McR4Rd9FVOAyVI6q7dfhQA+UrrfsTOzG4TF9KKvTNG9euf2V+FNouIPumCTsS4zcLNYswHZUukVi
q5+ZuBkSLwaFaw8cRL9ck/tOCQk2j+d9nMzTwm9URRMkUqCLsKh2VLjAsYMAwig2PQh7tQGymQou
Iixm1xm7FERl+ueUPQKLlg39ROiTSVTkWaEfY05xqvLH0KpnQiJJfwN32XY/6bfzYfvQbX5qpQwX
6Ok2Ee6qxJRcJ/Sz81D7N6EJEfbTu9nWZMVsABag4iMF+HCNXvewxyl2EdUE/bE50TONirn914TR
QpBTHqeZztm7vXwbzP0wjjZDe/9vzWbWSsRG3hdOpFaoNpvsmDNl5qDd0q0nrWFHWxDeAOnLWuUk
faWuv3Hb2Phl3BBfS/rgE4Ye0oOv9qXEGOKsDfEnK4+nheej5ucCN2aRmotcJVh990DqnkH0NKKu
P3TX9aAWYY+t0Q2RoAK2zje+JYgbcCWsJVnkrOOg3mt7Fvs00W0vljBg4KFXJvcLttg/q4qh9aUl
S86ImJtU1atcv6fhDf7RCmw7RzIp8FCLuOa5grku2dsQNIZzkgAPJz1KcJUqeOI7IUGUZs4Hpm2l
oLtexR4yvfelIbDQtXPQqTf/pwTZO9u/GXELXzh3Uhy5zC7d0IJKpMRHEHXtiid9wceVJxtFRfbA
YNMbuh1hshROqtlWq1/TzlluWxEWC6YzBpGyscvBgA07P1gMoMVf14fVEW2TX+gRoCoUyyMxTU5i
m2v5M/vfIeM85w2P5uDpmZ1qwtMU8HQv6p5iksOIYpbMram9b2cgEKYIrVRkB1kVxSLpwbrpbKWD
YyjXQzXMXH6WcqYF7qBqN7V0vYMgJ2xPSzrwhC5rjeTc3GI3jqVSViV5kQf6lNYMuAV0jGZn8q4Z
ShbcCLqXJ8+Hk+c+f40L3qej6Q3bY6qT+s9ghYnDmVzQh4LaD71NdUFh2veD6ZVzr66moN6p8Qkr
Kz+17nVtO6PqHJMPDG/DtgwbxIM9wcLUYEltO1EFINl6hOakoKe9PUFuqsyWANqaWm4YwRFBdnP7
HHmM2ouDzaIAkUng3dPoeso8ue3on25O5LjXCSNDtprBFs4Y2GzujJ3Tumh+LbXsAwmIeGIEii7z
lsYIxVLQJ3TE+b16ElHM3DJgS2AbwYnbkUE8mErEZ7GgWjjjfteLgKO3bWynsx4376IRXDuFxITW
PEeN6Xgt6RKkm+TnFwW3A2tb1z+36v9PCXEmoUYqAqUXKvYnqMe5yPpeEAkVj9QREIAinLVNHP5v
l8J9oGqKkABIeI1MnDGzQfT/jv4V2uDZD4jbjpi8CfsQxbRrsxpnTOxt3XTdoVrPPQbIv4+Sy9TJ
JBf95aCluWKIsRLfBU4oknEbGLSaQQWBPv8Kfr7CpN/ho3M0FfNl3tX60hSay2MN0VNnLrYRQ4tV
20K4nH+IQ+mVORTzcW/Ve0VnxN/cQzpWbslwNNoMOD6rnpsCz/vE6yVY8/YjHYjsTrx8bXRNvzVA
pi6uZAMD232AXOQ6bq8A5/B1o8mGXumvgNKbpWv+28Otm1bTnDkGuqlS/Mfam6IlYlPtc+cixfwu
OtqkG3/V75mZyYc0E7rfANoX9BBHl/OJRHJdO1C5K0w5r+V/Ualt7FWr97rTNHYb0Etowhlcb9wz
ghmtTaID8owVPRGb53STHqitP9a2QvEYdliBNFBj0Vsimg6gQhIm/65bUOX4MM1r7qLkOXgAB/qG
EZjyoAPXQPS80YrUeep3SfgwPQ4hg/MfK9IExVuP/M/2Ul2shEA4uX0JLhXaXEwseG9eFmnAcmDp
wIHQp0w4ga+b+kAUFWBTMWPPn1wVqpTX8PUT9HWpk9Pna39J6EgKH7LT156kXT44WAMUlUR3fbfp
wxFUq7UiS0VKYSQrnMqQ/4CQ68ffJ6aBFUQvIcx5eHD8FwAPIX1uBgXOTgVTWhJMJDrpG6RBy3FW
3An9MvAcqazibqHWnhL1buFW+CIAcBsV6DZTOuRUN+edliSWiUaua7Vwf8VAiWWeltJgfZbki9OG
qmD1utlHh3xrBWpuPtSoXuB1Rdd3wVm8EtaPAudOt+fCnxIB+eNkNVCVLzuqatoUdgZSwYI9dt+u
VYwZno2oBbtIXsPu3gQxwQQF9/1Rv6iRCpMPTtzzlCYwMNKCQnmqm2ky7es59IOYN0L1ZwAmKdOx
SlGazH1GqV5W/kOrP3SRve2SroODIR0BBYkc5lWopArOBGQVuc1fCeO2d0ZWJAssRm/H6lOiCQD0
Rkh/OUFe8PgCOLm5eOIrzZs6R3VnT92HlR6Y8mDozAxfOJeTBfMiFc5WmlDD7vK/50dTPOdhEOjd
b3K5fI3OCJX1tS67U28rPNBWTNfCVEAuWEH6ybrA7rUoFOgSvQE4GmpQVI0vP0/iqhb+xM9LDLO5
aVOskNtJBN/+aEuueMGhiFGO6Bayn1bmivTffosnAzIjqS6HCxkxr0ZqfWL/LlMr5J4Patpp4CCt
VkpMmHBNLrKy5qIQM8DkzCqJIw4E2hhGBRdWmyJRJe7G5IUJfxftOErFn2RAqzjGbLAvIGfBwEwx
EW9R7VEPrU7CFpZgg3Ew7S478CYdw8rjwJdlCf8iPfb3G5Wy7TkBJ9Mxh9XCbocOibRZ0+L4fEk3
tNbI2oc9UmhXn7KhPYTQOtqY87i4ZYk41VRU16CyKZh6PZgueCZK+QovMzJIUFsjWtZbT5b/0SJ9
jxsYRBHvRekyunRuWyOAZ6cgHIfQ+HE1nCd5UTgJRAFPbA9RWCYpKnmDKKZMDGsq8Yg9Vx0MVhUg
lrLDrftpNQGoH2A2y4lromWMO6Jn4duYkfvp4S2dj+12z+eMVvlsAcfg3WgiS60MwJudOYRSe/lx
Z3VRs8sTrZvXE5V3r7Spd7mGe2Qr4VZIYB/xwrJRev2/7BjbH0s9QesEFT/fAKF0+LpOyaQuqo44
3RJRfvRnF5ZW0eqdCzmypoclQR3MuqyE9GCdfzumOBwVdmlOcNjAx6EnSR3T7oA3pE6GqLkYWvm8
jP2iakkZ+dmfuoPoBYp92012rJTem3ttsschhDRBZsi96Hw6fjV2xiZwU9Q2/zHYqatDwLn9pG9W
/8zt1ZnihlxeW2aRGIQpq9Dc2liliJBIqcZ2FtT5bq379JqTP2yzZ84iRgWmkHTMa55yW0leTTSN
r9UTaPjak31kA3bIDvmORhlZN+aDGsKbAneNOlT3YcCLRmu1Xu8XUd8gVGVgW/y5gcNTapbny0x9
fUo6n5mrtw7Thxl6v8LK115KSflBJMIuMc6csbEaLxG84BAPnhWva67WsQO6XmrbYD/CrMzPHNe6
AP7ziWVgiIlyoYwSXl7vHurA1gdiW3eAUFuieUAVnI3zKcsYvZSCDo6/P9uEQ8t9h4ycE0vAhTRE
HIudUJfuJXVXhBd53KhQChQK4j7uvDZJKf9UJNlOhf3wlujWFkbSgquXx+JcNYcQKylsWVwV9bu0
3MFyCyVEWt8h+nWcHI+HKPOeyZz0xaC1D8rCmlDn8nW1ORgyojla5KqhimzGj6fZdtEFbHLKRCK/
wE2dA/1m6eIrMG+FZWFdLM0znvVlmnPvek9i3cBgdfU/Wqx7mHWZxxAUlcG3NaNA8jq3dE32wecA
7AWE+zWFIqLS+s4BHYwPtGNwN9cyb5NjQjQ9jXSe0dMH231riRyDSBkQ2wrzLQ3l2/pcfHrsIlYv
5lmFnxn6Yd3R8mOtlSykTz5KqCTIXznPQbhefy5cx73MguN+Vj/gATcWGTcT1F3ZSSi5gn5MZ5iA
otFYoHiJA8rlyRAmUP6oD3oTxeOXMNTs5vuR2mKLBIRr/GpKEzDMKqiyMFd9/RBaLm/UI+k3qmb1
T56Jaq5iwS9suYV7jeWTYq8ZMUmDZrpixYxG0DsN68bR0s5/DyRmMGTXWCPmqf8kCQqBxmtJt9ex
lcu7ZWKRTlLnDci+0S9UysW4hVk8tZLtEvx2hiQHKvKznaJqm94cJIzHrakSezr2p/l/9DO9XtkF
IS1xh/DQH79XKQwkVtJzSLHO3aYS7v/IFXbl1T4+IvyV6jedvlJiyVuJVS79/Nw8g1YXPpzfHHDk
sNGc1kw2h4Cwo6+V0MwOLTcW9WKWHRRcfbDfjrdEFIMSk52l60x24h2MEwJHrI6Ru/LILs03DaCL
j3Vj6fNneT3+GdaFsKmmBzJ3G2fuIkv0o6hhfBiw2NGVUTExWw47owmmj+9uZJ/8fRIdW1IH9pc1
xg4SwbtNLkT2f9mP3KJR+6jbeqylm7AnH1g7BVdRIIOUAnhgmuBkkRGwJ/tHanq9f3KHxxPb5Hq8
qgw0B93xtjHXNRCrvRg0ig0z1lCNKYlS4J+2ZiP1LCeBRdSrGFrJYPynFzQvKnpVC5jOZZ60UYf4
RsGnVwU5+F8rRY0TEfADmN5LSBQc8sdxwVW6BaI7/Y7d18oWMKmGO+lTMc6dXDEC8RjtntQRhm08
bL6aEPR+cz2WCAjwfrw11XbEYx3xcVlMAqienLo4nfhYyNcY9/1P7wNQ6ynFOpEZ8wNL4DW0dWQh
7jjQyns0TdgFEnx9tjWqV8E34MyOi8Xg477iMrABf7ccAdduo6PxdbRZ34j6XSoxB2deqfxBW/Du
EjAkzfwAuCw6OFUS0Fw+5RTl3kdfqWeC92zkzWZqYySqQ4ZuASBbHwLZB3YH3JL+KwrAPMxe2uDu
JO9hatNw2IafA80geEp8PfT7unFMuphdVUems9YdogewcrUF/5X06sx4Fbhn2pbPClUl/ciA928V
pCwlTON/RIfuBzMVXhACk4FXXjPfRvz2nZOhVhOuOFPUaqIMpUPbqSxfzkJ69rTVgq+uQb/UJOjq
QHbaNzM5HFpJFsQNk8CoBHsdkRy3ZGbNV6wc4eubzEz3N33yml0WWrYO8mDS3Y2OsF1n95bCV0e1
N+LkHfPNOhrtK/vduqINvrRU3Yq8VT9uNqlcaiwN9j/3I4GqSjQsWibOuF3wQWiSThWTgtqpOjOX
QUFUX4Y+AlQNtfsAtcdk9mEBv8odjwX/qzfxBUvjnr5C0EEuXyJFIy9sEJfh6DDPuyu56fmVos7p
oqqynTSg9FVehyZTjVB0kPv4PlUxXEfaoSEYbW/Sh8vqdcx4LFN6FzTAucOOJDSESwhocWES9yzU
l/fi+zK+NXI7ROvT9t0fE6utTWpcp+d9jm600oesLGygNaVk/fJfrO5KP32NtF0O8hJxf6Ye532n
uSiOGgbqT9C6L0P9swbnGWKgjhy825D+6RqvP8tuLDE7k/u2pffuJ3EXATk/uWUUaidUCvYsiRvz
Gn5ap09mZgiWz5olQ9TnueVDA7rtzDkvsQhO/p96afYW6MNxz9JjSPU2MKMgP+L5oRQbyzZ0FwuD
eogFrXy57TmEr5WNz7+JXH1tkqfH0AfFx2/EnrO6u9aqc1xficRj4o4SxZwrUJPjVJwlES0T7Lo3
41Npo/NaiElJj++p/DwIw4ohkn4YS4JEJGu+s48r8Duj2YwU0E1f+5gPunWcUbwq7w1grhFq9GB1
r/PU58DLOc6iHj6teAEa2LziFMiUk0W+oRivoRxO8T2IZHZhaILiupVTi8IVSHrJasuUBYgvnBIc
fce7f9bhX2Lym0vBaMlbC58e80c00jrqXcKFMIC2ZnGGF0WLaJtNwnTE+d67y1/ehM1JZKitdvpB
pSXRLGdur4fRUCDFlB8XaVw6vNjDTadx4JTDvB78MSlrEH4MUgZaWzeG6uWV7eMP5kBvJnBdNOAD
CZ1CIOUxbgosW7l0p/8WNz26fnJhMlc2f5E/+f30DSLWpb1mBPG8q8ZlnStTXV0hxMIhO0Zb8XmY
WZuV09JqSgLyODi4Zpxkns4lJ9WZSChrJXobpxzu6/wrDV291u0lOURukJnJJWwA1VQQZ4C5gvLe
AKemNDJyewgerh4zg9W8NCj8iiDmzFAv3mW4NjBLENcRlKW6nM2PpyLvwb1ImO+0UWy0fRaGRwqq
1Pa/rQ3SXsgJ8hJZCi4KB8PyNveIvaBJUTYgNcfKMvuvh71yEIAGtpK3Qt4ka7vHPIfSVl8Ink8P
7mWubbi5MQsBKv+Ge6myY36HOto4lQWK2dR7apcgQ89O1XVyDUslbEZgP9q5nhAo/Hl2QlSy3Cso
iE/7HgeRdUYsZ8Ypc3DorONgBKkmKTNLFQk4QyWmN5zN2lnGBwHeid8R5NTb7kKJodqpnBrQd++w
YY5P8X4km/SGiPYWowD6s6fK27x5tg5MJWLeSkVLE9FmCskAmKD27he5eTTmZc0DSYdCforzmfF/
Xl041F/cjr+4l9rPF3lAhMVv3jlxnFXnhBlWrJGM0XIyb+RlUlRx8Jcn9mtULEE/w55ZoBhRawws
Wg9Rt1KrrJtmXIscmjfQzWcuCe/ZvNxbJltyYVXXmNztvH9o6egxOxlirOZBEB2bV8c3R3BJdzVE
2qI8C0nWDxHR63zqdpcqJq/VNWosmD09xUFgMreXTNXEP+wNA7JFrqHn27Ywa0+3LmhPSNAVQpWa
4DReil3ycHi4fYaxIlfxHbY1IpRSAY6hZwi6nvhsHI5h13I6dazi1cqkpTVxlWJ1I8oE6GFD2U5a
9Uz1dFUV5rE+v3GokaJg/YRfNUvLOpntfqhLGiyiFhdhlO6IpUfGPcTf0iMly0EmQ5jDjx4O/PXX
xnSZxg2biZi3/cqq+YTUN3ZDjS756XStEC7E+ax1Q60R324bEI37I1Lr527vH5lnoCaOtw0IgRLv
bb5gAwrcr14FROG1Did1WR4z2schM3uqcWmdkixbXDXd3j7wkc11g2+k2ZriNjEZirfaCqaS9iTh
9PR6VzesqX5GumQB7NUxvKxUVz55uzL8XOZDq4ofLIL8SaC+Sup5rcUhGsoqQOymg/eAhc/2puaU
Mbanktgbc0LBAkYaBWG0/mSdZknEDoYYWZamNZ4eLznlJWN6QOikdA+Q774pQjInn2doecB2qPk2
KE5BdGLfU4oEdw7DkdbMXiBfJVg1AIAc1iEMjklbBwZE6RmDSUiK/TgHM306AyuUQK4o8rZiYl3M
Agi8q7K+9YOR4n2+jrShYmirSZ/AeA9q29+5+Ar7ABk2sFSG20U06hEESK9OObT0S5UuYHNl+1Ba
SZJBz/pKwcdpyrU2Dk7IjuSG01K6mGzDiM0mUrVf9wVfLqjCnfynLKtC+15qrKkOsnn81iHS0/Yb
tNAThPzgS0B0KkvwvWJbAn+nDuHw6WmiWHUjIz7Gqu2EfeaNgoFX1BTpSwfEshXRVVOaxKZLwwEU
94qADHMqNPQKX168e5wmmyx66ICqWghSEKhKvEdn8PGToSR16E/rUID+Qrl6Gl5m8LInngQIJtk5
b9eH70IDOTud0M/k8z8ltJi/MXHbM4F1pk1PKoB9e+NEYNzHT0MCxYtdKBwowrRYr+eRESPLrcVq
vSkaT/7ydEMq+S92QpE5QJ//qFKTAHTkHEHkUpGOzcqs56sXeg0fvyqrhzJ0NjAaWI8UQ4g+Ld3M
ZbxrCTUp0S3gqwaJ4XHTcfkcMELnEhNPRi3U81wSaSF7j8wu9xLv/4Eo9if3Zouw7YXHheNeamm+
DLmFwA0lcU3W8x9F5H/1Jh31ml7shH1P3HdtLw15YBh/fbbbDUvBQNYk08kjtuq+wikRqj4/wVAH
f0TxTJ7AzMkNGUKntcEeWEowf/4/GtQhQFZe8dge6f1ByqBQbRiYBX4KqBLCn3a/03STHkgQwuTl
VKw8K4LSs4yyTXub4FWfvs/UTZKGfUOHJCp9l7qnT4YmX5/e4UjyAy6VGDL6ShEwitkuU2FeJ5SO
EQFWMQxJQ2/2ZtzPGegzzDx7Z7e4fn0l6WCbA0qUHhf5Y/CWSDSa1DuHhhdDWlqjOxZCIj7b+kap
FBFz5q1/GVpnn9G/Askt+Ghx8bS+6a2KhZMHdgvxMNdE4fZpRU9m9eDOFAqm0McmPGDhsO+Q+Yl0
hc664Rif5VSNtFeuGWR3ZDftXy+4Px1EtrAxkgeUMbp7p4WHVnAYYs0T/864MAyltNdOmWmuThU/
0VXBYMFkskqegL0lkBzk6WZZGpmqgDAhisGRH6tNgIRps15qsQsuBY/JkU1QdLrmvBKKpOHwy0S6
JVwx4L/BSFEpNu+lvyVs2OAOKUs1jbqf9FYBbgGJcbOQeIf7GWOv/9abn2EVZG4NxniUjSbSGFUL
O0WEMIbb74SPwIB5Wr9DX8+XjE59WqDxll6BL8c2FY65QAxvZYdfQr5KCwvA43G/0mDwgkPfY8UP
uOClUarDSFOVBnEryTUjkh8WxMwRa1aYgxo6tT2xxrPhvGvfi18DlCfZFWMQi3QOV0acaAAJFvix
b32xw8ab/8FxV4U/bksFFb9VwtuahmiFdEKu70KouT3GJpwVKZbfIif/iTjs93MzXuRZGrQ4Lzdo
6/vPYWXoZfP2z0KInQ2txwAmDoOjY9XQ+zLBFKNJv8/YL9Q5j5621Pt9PN0LQAw4H2XdZ5oszCqx
fMOgocgHbV041qWD1JdPkZIiqIqZiMkVhXjQz5m8W+J3tT6lHbF80f8Oqm8rS7beFMU6XKs9Tf+S
HmixHWden30ky7GmvdTkTvic4rMU59PnabSd2hPyg4hB0zuem9zi5BDPxytrf6Ws/aBci8NTMgfb
M8SUeXiJ91WbX3mppTmekE1mo/yyli2qvEcx2F9QjOKCXcHDMYiGs/DzETLZMffZxveUmZJH9YyN
Xpc5W9pdD7TPo7dx+6OawwStLLWKHTtFk6NY88SDAd+u63m4Tu6ky2w6zRyvH6Rs8Ov3U2WF1M4t
J8lIqojiTkUHbjiOB7IKU/wpz6qJO5olfrqJBqztvebehxDp+m488G4sMXuIKLZZriPMB0bzHCzz
stnNlk1kFQSeHY4xBwmrZve4n/+HDxsjSwu9UUZQ1jFUk7fIugP61kNDa9QP+x4cxb3I1DRuLyuS
RmaPEQS2ycJfK8lx+VlsxzMQO9nAg2/PQmJKJiuxHUZLP6fIvmiZV0QLoqKC/jOpvNdO6ON0xYKw
ndVRkDqrcibOYh1l2H7/mKCxxRQMCgqbybrlqNKnyo7iphdmZKUr2QqBRDktK6crocwuCp6BqXJ2
obFp+Jk0gInWsHhwJ4g/+6TtW65vKucFM6kOU7wGs7FxU4mWLfx57ZgJJGQYkUz67XE2w5F1Garo
8/UOZBk3DXS72eahDjrr8xyNpWTc9AgRhfbgGpH7ETEkk0oNItBhpSmsmoqmxwyUQfQtzbAlaE1M
+yB67t4fAa4sypRNiPBoW0lyD2VRavFFhosHoRcF4j3wUg4SWOAFxDZBMC71p1OveYufa8xhLtC5
n3EBF4WiPW/x4uLja6BGPdi6XxMXejp8fbwtDO0yv07tmQVUooj3NX9rfs6ORaJHIYdzO8ZJe2VQ
n6NsWJ3SaqQOC9SfZJR2k90w2H3yoD6G+wNAKCWsM3kQPNFeyr8V0fadR3VLJh6e2iMviEozvjA+
OVY+R6Kc47/vkB880CDqBhKD9zz1fXApnPk5Vn7jhqn/vnKLfGJthN4Ubpejq+yvWG+6kbSiDPPx
vEe98pvyOd5GLBrI5cy3kqPipqrNdd3IGBwZRAAY48EXkkKmBa2KaTg8C0YAFlaUSljjYjPKa0FI
xRfQ0iLyE9giDVvFZT43edmwcF/rfPodlOQyxdpecDtOYzyHWH+anfjNu1jPV9D73u+kwyI7IgF0
VL6YpExETiQQEYf1vuQUeZKfXR1yCOIuBxH7DdAmNLOV4tih/Gevh+qqCFJsIAo8Tvtgfcxe7IuY
bHg3foYiUAwB68cY1D6GU27e2kX9PMQFLEfTtUor7vCu4NOZEfDk4rTGpwyLEg0gd4wW3UlG3Tx5
cIviG7KoiPHnsZ4oyf97pf7t0A78wFrXt7AjBUNvj46+bOM1WsoWjzg9nHkquv84NpT1s1DfBhxb
GAQ7tk+LfksSKFtvtXwffvhEqMDSFyW5AEFVorzNbG8EdUFgFShKu0GSAENT4c7gCXClkPRC6I56
9iN/0V/b+JL3tNt3UgBypKr3lIe5lugTHzPoIeZTOpW8EYpWik8Vv7lMk+tZT/kUVWVeLvxaERow
qZBcPym5MWHQjHuzTCGwzkH13WA+IyrwlxpCsGvb6kbmD0AtKBgPHkLOJV51rkvpeT1Vdj3iU7xp
nCG35wfF4suI21KZm5SpfucstbTtKKe9g1c7ulJ4/APWTKPYBh0OT1YzXAkQLd3WaUbIzHpF6aOq
yiL+jqCqffxs96RpL01pwASH6iKCt5QPHGxgUC+SHoP1JOyI+VEhW45Iw3I8meogxkFKVUH/Jnrs
2/OtgKaT31K856Dt6Jr+hJNz0kZ0NIOgExpaZLmdAgNI9IyYIhTpeGuNRT+Izk+cVOocGC5HIaVk
HvwxX7eMRj5fVuWIU5lhlGTbr7kh1yfD6DHBJAVrULxr5q0oCsqTVf6cgIg4sYGp0u8gXuaiCcEX
JkSB11Mg7kz0Pv8QqvGJq2puZvkqff9xtoHRHwiAA7dHi6YCUghdlQ+26AK5uyqsPOcESBihAiC2
sv58SN2ds9qOVOKalND/u0pKy148zugt5bEvtoQZD8aCszFb6BSusXWLb+LJB/JQhetQ2CODdy/p
1L+UGLD1TWGroy63Qq4L9doUBjOEtdjpdd0MisAv3YnU+d4N6DR8E+WTAbN/Hbje2OB3/kw5NK+b
33XRvTQQUe+9FklvZ/nuqwmYunT7K1l9ElXb/dUpXrG4ywWVIaUMZ/1GDGnXFbvuuyp1lJtEYZSP
yFmB26xwuPl2D4bivnGvn6WUSlzpcK1Tk2k+0UVkEBQaZUYM9tEww4ccmCntvVm80oV+dZG8RAdW
jMzlrj4xIg5P9I7MBhOI47woZdaBZ2mLPBIsMEsNjn/zYEGpfQuKBgYHzfcTJ70dDPduP/2mZG6q
6iuOvPVqZNpTqTj+6Az+3paffbp4+/6DT+PGoc0o4oOzxLY+5XLvX+UgMtL/6M7ILRmXkchTbDVa
2Zne1mGRdbKhOD3hZMSzURN9kfZ3OY3VzJAiHcXgWxuk8XsquijPfV4ShzfQ2Z5DMXFgKvnLqIWJ
+5hx7EJgsE6HfxE8179XYo3YA+NOeU8dNjrvKFr88DYnrpMgZ1ihm+2AE6qP5If6yAc3UcPb8hBL
7Ls57yqasNkwYC2tWM1oJNQlnCPFmxWLsnsC2h0mUsyM+E2RUXjp0l/u+3qjx6rowohXKSWIhnlR
QG2rnhAF4fQqeTUyGKVnfI0/HYcnQI2h5mwbEcfpZsqZJGjI0fQyzBtSj9xtNvxfH/nWrV3NBFES
6noOBwVDIUNGsud3dUjv3ue1tV6yT05FOBOM7CAA9HrKx+h4LgUKb3VTdzLZ5zJx1oUZNL5jojTi
+/PIwND6NxnNFTMCAvMWnVwBhIR7zZk2TSvq2rvkff5cz+DXTLGIf/scgL8tdcgCoXT/+oNcBArZ
SxEHoqqH6JoSdCgp8Euusy/xrBtLdEU+81L9Y5oCWYoM4WQUdsQm0wYNVQb9AuwR1dy0bNIOegR6
yzPhNBPhLZxwTflTLNh0rbj5fdCm2xXNjPjzDa7tn+GDuo/PbxQGkFEjBl2+kJfqqwuDSICbNPba
NqZq2KtR341Y0DTTNnzh+MpaGSZeZ+GjSaU+yCglB+XN7tfNeiQPOHPLVTrrDCtD9o+t3KMoRgln
H/9itvCb3N69T24It7SclsuUW2JKihyhNh7YnIN6T+Z6bXWsvGArFCAt2b115+pOEZFcdolBG+s2
5tOAeugN+zYCEWdWJkTKp1lkB1gHQHl9aXVayUlzRYLE0S62cK6AWLAdb6rCJQGDqbNmLaI1DCq5
KTgPe8OVhzhsEyKbPkhj4xjiLIdrADwgYmHWaiPA3JFHe2OIKLx59+jxa6hYgvWbjriPysZt3Mio
IA31pm5qQ7q/xQnRnE7F3/IHAqmsQn9IFHPX41kQqK4Y7HHRNsUuDtIRab5XUt68oG3jEfI4uhBA
SsqNmgvqUM5j0/6J0TzYD16Or8qxkC73i0NjOhJk4waqpplefPp4ZKHVlo1XxSgITaKwACpqW0qM
UeN0MfTTPgDU8Q/Yc47nfidzpy0DWrysCTPNXRga1YNYqdryCwZpCKrt2m6r0ViaG+fQi8dukMPr
LlSPUl0Xv44/oURlJ1itRprhVS2bDwBTm41CiBZEKmf9i/pwI2P6mjHnS0wX/gCtDJnE6scUCs+F
5wBMejGyVERAjpc8WBWJxvyEy0r5h7eUFPzQ6/rEdS9PpET78DOS2GT4ma0qU/g4wSVy0un34Ink
IP7uYyJL8+8aHYH4cFSQ/zaw9ZZ5vMEP/F1W6gE3N4nTs7BIroYFMTS7Wt8MG9v0nHgIlsHKzQqj
1PF/Hw2vkTaSUkXK1rdBDW4bGE1WTmyM566WWqu4cZT2hhcomFxQbENotFFIDITFFGSe9TG9Hqn+
4qX59gheLB/FdMMM0LITKd0c5doNUFIASjpknQBXuDb5m+RP6fFnDJsCv5FuFu71pMb3mwha4Tnx
nm1mRHgAVVBP/cPC19yZ1SUYXRUUB0CPOp3f07ybRphj+FdR91Im8gBK++VDFfrfkd5UELrLNuEo
QEIH7VLC6T3pZ4jwGacz/Lk9NfhQ5ghh9zHUlNv6NxsvkhTISNFtrwaOLefUdMXzY5Q7BFhLSgKt
FGC80+Ic+faQqtti19SGcLmug9YaYgf57oYq7lrUwbPLJhuWqayPcTr7gKuZpy0TddNReVIbUP3W
iK0hBIxTvTanYjRAW8mdiE1noJFVuxyaPrbxe9i3jUrvXK6jCUPAhSyNH5QU487cO7t3rTTRiD7B
vx6HqkWMR+MfgdCGWZH5PIp9Ia5mXsp/cEbtry0S74Gx6q0jrDolfDvgKZM8ai9Lw0CFtf/MnpF6
JyOJV0a2EwHT5kAjJs+LEa5NFrLAZ3rPlqADU0BDFNHHdfQg7MuGzpyvYsw7vbCj5HNm4KE0UUs+
Wsgij6THZpz4AEGOH/hWc+iklD4onD6Fw3oYdRYk6zdVjvtblrxiDV/CkefFSWBin7ZxOoN7BtkT
GWdCIv3gEwV4ex6ZZy/zTgMCioI1T+KS8HdpKIxlvICq48WUwu2wvjiu34Q8/xpsCRHlmp25woJi
n9VspZGl0xN5By0fXkQ00SzssGHrcgrSnMtefI2YBRb+E3mNkL/byul8AnLf6mZUPRAVtnKq9VFt
bWLhjD2QT65KnZwEZMEjOdpcD1+Jof5kxBxg2p4ooCsTH8KQbNraxQRfl0+fSQDIr7Ut2e8UF0kX
RABF13dl/U9xfbH8Kah7Hf3OhSTt0gCb0zA/ZpVzztCX2tGHGoPv2eUkeytkjZABN4jLYO1b1d/2
PvmOzZwTSkivCdFqpXkoWunpDZ39MEKsZSQHUlKzESxK41/L86YQPT3WIli4nELQnmgNlYoQZIfC
WFd6+SYLAxyLMRv+VBNGIsC3QJDDZt8uOLC43gc+pclSXkwlm1aXvRnfc2ZyuJ5JJLUR9dpSK7Nr
2rNmq5T5KWmbjbQb6eK6dTNAgwsfnXLKmqrwCwPhTQ89DnzAwSbP3hRWaADjVI28O+sGecj8J9N0
E+5Yh6PCY4/7Ep5e5RH8igW9Ve7o5BbWn0EjYO9NXiXnesoUp4PIWAl1TONKXAES9UoUPGG7DZAw
Nv0vAMJ8wphaut6DUs+VrYPlz85W9hx7SS+COGbhQjnK1CINfxOKK7X9MeKecedkV4SAn0311xc6
F0oZNhkavk/P6Wmtrn9yY82lhugqYeRFc31dX+vBVk98FpLPVV+aan8jny3nSItZpztpn9PIXrN7
QRL9NNBwAwknu44dRcy7y7++4JEzR68doQlBKk1Eou63rulQH6VaI/taQpTHnVQITzyNoiz9NjqM
ArjOvT0p+RvViU3cEK2KsmZA2KIqCs1wVpcCzFmJcnPpiu/RBGGDy0sywro2lPfbS8TCZH4BQpH/
OhAYHlvcUQneD/pD+xBA7gspqspj7Nwzb2j0wiGdnpZbeJ79v5PRumTcy1rJ8oxHTmcX+PnNwlRF
GN7rIxhFQP2oaP9/jdJtF9opzrkjEz9ijK3+3fgnadDq1zW43ZKOo/JJZMkO7RyOuO2Ix35Sep/z
7F+8JPEqtyzXrml80AGilfaxLpyIE8qA1hFK3jCuErsTKJrUaxzl+g8pzyrawRYjg7Buvjcg7g0T
qhrPafVmarYPUh42lkvt0u4OE4bSRwR6/sv/KakYS27xgYJQocWt5O6YLINNtFpaVxWC7E8c4Jxh
wfu+SpTlqkwf7fbv/tmxmbhR3eI/TXRFQZN+Pk4giesDaTUwb5cwU8Uw44jAYPkV//mwSB1KXEQR
GfgT4cbp6h3JPVDXuiTX9qWPSSMQ2FPr29nMNtji8MUuO5V8MuSwVWhZIo5uoGBQrCqcu3f0EOvh
ZBylI0W68NkAmaDgCy3chDMqLItFoWKOF849jn4d6PMfGEIpEbocNOZ2ct4CmblnrqUNXj6pQml/
6enLJjR8wcOoXPhKdj8FgHRn8brG0fKwrNophKV/gG159C1b81virCDjVnZ7+zbNPqKXn7/GRM2Z
r9emYcfnTSV51Q8/EwCDTyUaKg6Tl771Havz/A/mTwQrprPVu6GgwJZzCze4491nXEAVLvGA+Clm
+aLCm61lhX8DQyRGLE3kn1SY2hjwNNSjDU38t16uer7CmebX6AgnWxZYuWQe9yFiKBfgZISCrVyE
QqCXMqWzH95CKt2FYiHaS0Z3fAiCuj5tMhl7ut49nHJ/lpKB95eb8myneY0xeucEurJWpF0K1msV
kX41rxb/xNl07yeDzICqHJ21bC06vJ4rxtrsy/32RMDVBKTl9w7lq5oGuGb/+s274RgCbPQtFraP
yaNoq/j66MtQD8GocCdW7kz9PXXf6MGbhe8Ob+uhgE6eP/m5M0tAXI5ddGPIdms3ust3S/z+NUQj
MlRhnK+njxT1xLj+kkl+4AFrsGw14Pk0G8eincDfJ/dwuICMDM8+XRkoykuKvNA/EoKWMe8lobXH
OOLl+izwGSasrOgJoAnCWdzOnzK+8ol++niMclVvL+3vsmk7fZGdAWMUrP4vQr/ZNd8wELvxjmkw
gLD8gYjomkS5k+iheG54atqWDx3S27doFr2qp7tH5QSQpyx2LZpC6yMb8vbrNzlgRSY1HbWHzeVJ
MAbVrMquHdF+T7KDkr95D6Ng4aYOQODYhJiK8HCbRvl3sgJESWUPLgIeO1vH0jl2W8gaB6PjoL5/
sahhR5I42h20gnAoO49M6r2uyRUDbiDIi/bU7afug5EgOniNL/HqcSkyx6H/MfWLykgkYYzPJP21
kl/8ChhvR6OFDC4Ii3DrgWvXdR6ZgVjiIzDj1HN1WLL0uCwZzrs8M9kkdjJtBov6pPFJ0NjqQGRl
7i0qEFgcPiAYjsrPAIp/7Dx4bwWWrCmYKrCflwnOQ7izw9Z/WoiDs7RwAUDXm4iRSW9j6YGkhYmP
matHMvjlKdbVsheHfHBaXi1gWqumSDsZVepI8nX6wnvj63mGAJe29dWF49xhB6p1sWm9YIafptGZ
cPlQ9bzEBS9qsmaIO/OydfLfKxsMSERF7wbJhmAHpV3M813cYvUqgsK/4J6AYIsbaAdZXDYUaL2a
ZqB8sIE74SJNi2K9mkGA5vqTIBIgpRUgiqBXbdRMw0Rf6qPu4F25WTXWkW3FdD9OgMPFTt75ZT4i
iFzCfjCeF+1W6e0n+dzt9RufuvQDgftYEeaoKmXcd11BjF5Q4O4GdZGsxwcQixMjOo8CyKX40Vt1
911yrpni1Gok1T3wsC6YTW4fxSdS3jfJgeyrFw3MCWYFnsOHE/CigTmF2doPxg/uR8bWuKU0zXZF
jTaSQAuO075efhv3HbTx9Y3OYFt4b1r24LoRFisDOHtAXXpZqni804YDTvjB0SXvFjmCP8rOwwVX
ZmcJgDjSNeotXBmVj78IRdyvM9LW3T32yTPx4fCWy1UjDq9LwEDlZlvjqG2tWt+/C/YpgPVxqShq
9IUlh+5uVwIYNoteWgqrhdrQ/7jxsk3o1gossh9H8ub3r4jCtKxkDybvdosRlrdE7lQEknM6I651
GUkyy6WZajyMqJzL/DpLELxOxIihTVNuUIOAfjqIxs/JqB0TDOM/Wo27ambHfXyAgle4jDCjHUPG
kPe3uG7dvx4qX+RE7MhBKRZyQ3pGc7TcDtWF3HDQUfhPk2yzud+7JdhoThJEzK7kl6D5ec4czef2
5N1EYnStGE/vuS6OmguZIYoDjxMuOKWbu7xJvInLEzss/CtjFHIuAtMmiKoX+9nYLRQ9jvVhH2iT
7Oh6FAN8Ci4mrI6gM6Xbk2lNVyE//wkxiFOgjaCnnsiBia0FDoXpvFvKXzM5+STkAMUduAY+22DZ
kXD6meUznJvQ7r2wFAIG7PIbEa8IBBUmkzvgOb3FlpcZVDhQvqRl4K5RRLbTdrriuIsGQbx93Jo/
nzMo/T4d+0+EZcvVhb4MDnUn94oTHHjxkwZrWrhR6GlYm9OnWfkCJMPJ8sTgFUhWahyUXaNR1eLB
Cm3oDVVp6U6x90BTV5Zi4djDX40KlOqZWcKD8e8wpqwMjWOhFAXl1QhtgPrgJ+qmJX0Mxc6QeJy4
M1zgFEnu5B0X8eJsk1/MW5BbaIeHOX4Hgf6WFEWWaflN2OqPbBE6Wfzj7/WCUbqToqIIq7jr97cf
sO6X3uQpb0WJ6goZ9zbzmuZ02LUCN9F8rHTeC29Z7iMhj8ZCazvU4pq/CwqDBO2xhoKp2sgrvPa6
sYnPSEvQASTL9aQFUl/luozO5RwfaWuiNJ3SREv9r4MT+zZqnaXwGyZ4UA2ptcWR+6XMfOc9/Lul
ooGO60vjN3nVEneBLtd6lxOO0ErH1dqB21Wyw0pyUmsjEonbIC+OTeItc3FVlOklLOVc3eFemvUF
cnBCCLFJNDWF/sLiWZ3Iu5T8yqI69NZzzB7WxK0+stRYs6d8ShbgcSDztfCOPTfXUDLccyz7z3Ef
67OmPUUdAdMHUPzsldpePC3+KKyZlmR8wAWYnIdAHOGOF0i3H55plRFOVEiaqd7zv6abbghy5h2v
krK0fKPZV1YK9aDoqgxqOqNsG+kN+SnX0DKI0Q9I7yWi000M3kDxDOw6alBKO9zYwJjUmBHP78fV
l/h1bIeX1bM/suvC/aElv+TrCDb8RgtfViCacloRNMkdVSHSpIihCO4EiZPTxs19F2ADgNjk5+QT
xy/LwBTmkScVMhoNcYxZcG3lxhCPrEEajWl9xjZIUBuNkS08+IBe57OsnCbO9xa7BENguzio7Twz
I8wAssH5aABUsAEmmixtbIR/HA4M2IvysmF62ZEIMSN4yrN5gwiqPWXJwOGVTms0aPON8mN0pWKk
Mx0B4d4cR/3yqHgHx3J+nq7inxNea2U7BcFh/ngaj0N/9zfZSKTnx272L7tip3LsWdddQnaKpeIY
xfzHh2mwQkcNaxGkI/kIY54qkZlkMH9kDLfi8Or/QsqBRF01iBUvCXuFM+g6CS2iwe9Fwj3Gfa0/
c1uv4538UNhfT+foE/OkFxE8e0zNoEUte/QXf+0WNhRFb8gS490A3iSOzmWjINVaatMKYjeeZsaX
SBC2nRIu90693BY0uwdGAHHyFPdaeEqCEP3uHpCA2ZI/A4MpVYKygFvfh5BY3vXiJktg3vT1bPZS
YA42mN1l0Z1HWcmq2jp76MaeefgmmkINH7iwrEjHzfgDdPdjOqwP8OpZ5wAdvahkHYiI3ZuKW7HN
+4la/q64WthdonX1mbIhTOkIfu8a0WMsCRd1YVSum703CocjoYjRVZZvD3+eGE1Clo12ubQqztW3
Y4oMIKu3ZDMv+C+bvhcJFURDOdHAHJn1qH3TL8GrPQ81/KJ68DGTmNB3dI4p8Q7nSJ8wD4felCaF
0z7I+RvHU8djxwAYIITWriduLtGfeWtnNB94f817c+H8Tt80/Iw1QdJ2qDs5s3vl8xgalS5aunXr
xS6MX6XZ4HL5pIc9AUoD9nfkaLFeH35zyIAsBD11neJKt62jZNabrd/5sNKXOBcfgUkQLfZJkj7r
p4DSuGMG74O++tV7ic/YFJeBhWuo37EY1iQgu3Ul0ojHiYyYFdONTg4JX9kRUiI+7BxKAqbPgfRb
51VyoYmd/kCvSjOM5wjAYFj1cAOixXLxh5ZeapDsPyEQcpaqChuZFNOm9Q4LNi1aB6G74JkbO514
h2NwvwSRKur8fJQWgsxA5keK8YjSyvI500Htg1fL1vCWF+R/EGRvZ+vvGMGJlae6/dIHTBCRIS50
lMJK/qdoOE78Z2DGW7b2PaP4hEFDasS1Qlcifpe/YR6vvfKXypHpXcLUhkbVWba7p/RxY0oZqxa4
0X0BLv7f2FBLxqS8l/yqNYCCvYEBzGq/zqoShph/13dDNGHAWGuO4O/FCxlgASsYUoboQQIw9ion
zJNInwQMQntdAth5At+igK3E9JCvhOwk94qtk7lbo/xOLatnYGMRWRtXrDErCYkrBEWvhOQ7gOC2
JY3m+IyFRnOaD1VbvkgMcs4dAmDwAqu+1OnJoFrzRgKGeM5AiANWJvZq0AM/o82JDOiJ4leHe0FJ
XMkceB7+0eYTU6Jh++uL65QuRIY1SssRqXdQy3aXk7ngmQeQhjGQ7eEOhgAZqQfv8fQbQ/Dzmi1L
wOPMa+ymwRcP8B5ACSXoLoEk29XXaf7wWFoebgwG/CMj1pa7qJ7C+x98zobi7lW7EOktyk5RCojl
toq+6lo17NCJLczW7Vmwj35Hk4YskjDR0x6X8pZnKny5cBrNk7jrqkMq5eE+U9NU2jmQ+8lemlgX
N5l2/3IfQaK7rBZ/+CI7vknBIblzBpLCyXQcS3cfW4y8ulnRmVUSUMxRLGg3nhEfq+YhWc7GuPa1
bq/7x9CuZJPx8d2dGB21z1kka3YNEKcePoFiV1NL+2SwV1BHpM/o/+ShGIDgYSCSx6roTL4dmgcI
ZigFaZgiRSwSes2XSeSfTj95D5DF/q4gyZuEhB3TUdVcumT1iA/uA51NdV2+p5oboXD9XLIG387v
X/JqkUgbsmrZSN5yJE6CRgERJmIx1wVcXU4kyfHKnV92lJSr3zzePIwVlrSeYqPnaStletWa+dmK
1lXhKk7JG3XibEi+NBi2d6On4R4M7uwLae+bCB+yUC/POQiAPoZpU2Kt/tHUBJ74032g+pxV8oPT
uC2eXmxB116WbQQywpuKNqoAKAc6erUNzox9hgvM8gPPw9UCPE9nSuI2QCmDI2kLS4FZ509TW4Eq
QyTqstF83ULbjKeGygLT/fqp330SjfudI7WWstBlaV3X/p7QpgSMN9Ksl9VkfqbnQQ+Len76DXTU
O+zN56RJSftIGaG6iK04TM8G+Ct5GY50LDMNJFPWOZffUFNOXlRC3DMnD8hBn1MxKFEXiKkrvMle
6zs9jLlkIsS593tEB3c/P+MrgD6SNgPeR/55by7lB8XpCV39dpTTdJ3W9EpwJs1G7JlYt9D2crpJ
cVGgXl5uHY8UjI2VcEH3+hHDEaEAxgYwJ9HUoieqOWYhLOnR0VnHEN33UTjLhXuXTzpjDttspkUX
zIZZYiW6iIjXbRrCJi/w2KMAWax35AuDn28jGEnr9nP45htVxoMO3+hOvwqVZ0oOLqCNNtOqmxQE
j/EXQMiSdbvR4njOSeOg/ZFUt3tTLvUTfPTF4d9fw6sMs2moaIO0AG8ngupaqSzE/xA5u+PQ+xZI
azGnWwM/WeyFJt1Q/208yXN6L6FkwfW5+c6i4Mfs9cc9YSE0q6BvdIFewC/RLS62bk81FkNadUX6
zAp/e4dUcNluvpSR0F+8UV/HOKs2c94LrfGkPNoTpHKmwsttyPfmuoJRd2NFc+OWjDXDNkNVVyGt
Wb7IZlljoTIkTNfAraBJf/5AhyzlPdvbnPrnOOQBCE5cl8SZ1lAD3kDLx/37G0Cp9Q44WLbuh01H
nk7K/e5k9KIurpWW6Fjog95Gqlk+HBa8+8kDnSajViqFyUGVrpyfp78fWycOZLoV/+tLu4tYL+sT
Ovr6nDfQekmNFzXCF+gBpRBlx932NN9SloW5hmQAlOl2WYoA8haul7fgnPQyaOkO6decx7kJacgF
sJ/Hket9G/wUG1oIovyOLUm+13ncD8W0lJKGdb07WUJZegvMVepTlXPZT7IJoNi/bc8W83KnhfAE
JGu/fthoVnnChqwSHjXjKqkuhxe/zeTKafyQ7hC5JhmsBjSPpMGzXzVjwMiqjVvWm+vRT2IkXd82
0IFyIWfxRz1b5LsxmSlzYdALDlDhQkV5jxK8LWDEr+rFVzd3WzNrvTg5iUqu8rXTq2EPw67Q66B1
i1YT0/pKCfiOGg3NoCPS9TcM7S0OHIjymUdpsQ2km5kxKRSUg9Ao30EYrztHnJDrW6R7/n5KEajV
WirVj6PzQE7htCVOIvUz30YJaqJlsaWLr4jn5t9IoC1XvXKUNt/qYUfCGsy/oT35jevrnKl43aqs
wxm7PQhcUGd8Aco17v7KwWozlg36yDFa13lPUH8EY8h11cPm+8Cea04d3wt/4JGXfByjhTwekFYp
sK7Kf6Ufaaevl3KM+FxUOk343HX4tHrcoGnnnj2Lz9VKc10AneJpSCmYKoub31NS9KjT0qExLv+8
Dld+khGtcVVRw+WnMGECq9mYh37uW4br9mPbTc3laDmTvhXrBuXi/1mPaR6+4ElsPCmMzp1GwTID
yprbCg2d5I7KG5YBbLKsoyQkECu/ZcEwAerxJ+dAKxnrdjt1VGAmy5NG1aMXpOBVyGpau6JCDg9s
AxsW2dIRSaGlAKi9WXJL1/yL9MsVXcPRC3G56+kyt0hYnlpHAsjJ5RbQJXbqkvuwyOO/Yv5Himjm
ppJuvQ/t1eU6p2zPU8C+V+DxaUVikWaBv7uFwb4DZrJ1ivFOwjpP+dqqRGzFo23pjoCmUTC0iKrs
Mu8I2MmBdYUukbfuIh298rcha9sMvSZfsH3FSG91GuVO6tCtfFLmo9iHsYil/VgfCJlNufxL3+Iy
NGik0tJ5s7HROo2lyuBNbaW+o5k1RcjtNo805GdU1v/ANM+WIV7yDTAruKvMb1SXVIYhc2brXwvX
EJ1Vjfj7TwCYM5MZMpnxfjIPI25HPjw9AXSTqH7j1W8sHMKlz9XGd/bT5WiuaPipUZvgrztmp2RQ
ZItyH8p9l81sDxxcWSFkyOWTLyAjOoxvyv30aFC3ICoLj6zUA6NRI0sKl76ANmslWZER14IxSsaj
MX9/0qk2R1Nx2ao/ixnFGg4pKN5Ln/VLRRZu8DgaHXpejRBZRXj7OisxRUmHgOSTbuNdiVcEJd42
a4g+m8GeFrxO1ubYkxr9JjN6fPX07aDjDRZcSGfJMxBbst4Rvgh9F5BYjVjEMLm1vXNhj4Glhki2
kdVQQB8Hs2e9tzrG4kwgZ/H6aLqz/HJ1qYi40Z12i8PifjgQTLO0oSEvQiwdEkV7fQoWmOPZCOa8
u+A6+CBqYdJx1uuJ1aLh4X4Lh8sz9uXqaOHjGotCVFogwX5cr4ix/c6PS0ySTPboYhG7aOAgy2lc
4Fmy4cUO9xHWX+LmdzX0cTuoLO6KrbhanusngQiZozgZgDbN4O6KqNMKe9Y2gb7Mc93ptAokvCdW
Yn1Y3odgrZf3YS9MFBaU7WJzLh32TPk+fO/NM4IvnqgoLzuNXJgSuTrlzT8uw0i8Xlg9NfkciFwI
qujFBaAYAdXGTY13U4NeUcAl/ev+bEVU0oZToQZk9aifbsh8sIozvsmq6tmJ8vDlw6dlKS83INKH
gLjIjtcK7BW1nWbU9QACZrc+LKliPoHuXymAHc4CtHx6g2fcZberhRfOx3oQNK62d2//qgkcM18i
CfO28I7UyOXXIOVQWLWXtWTMeNrbEnaV7CGEq7pXqgpc1i2TnVKS/91zxSyb6f18+KhLvs+gyC8E
kVMiD4DeGRlppfLFDZ55/Oe9G3oP/uXY4YM1qhdIcqgGsslSDjyo1eQ5wSNtUFWb882NKr3WQ/s/
mbpbbYhmWfsk5foQ/XubmlxqA3E6ZNRuZezQ8I1So9a1urr20P/Wq/JhHByrpv991PFamgwtidWC
hCJDi1oVOq/B16p7Jb+iHhkyziWOmUcWHEmuQ1eqBgO9xe9HbjQ6HcMMSCGWublmiwKwXvH4yV/u
+J7f8JwLNGqz30ASCZc3CvkR3wfhLXkrPiuXc32VG9eZzoToymX3FVswPSpHWcWFCobIc/tBMPCz
I9ndJ8UVtiVXMdpEaTjmtYhqVvmhQhPk1Vmvuv4nkZ/pMKiN9SWGamwYJhBrser122+raVkIXl/u
4qUL0G4BurXBKO3mX309wuuUS6orBcp+hZg4i4Pb+KsR9x+YwbWAzKms7w1sZOnieYQtZMO+Ev+l
dVCg61iEmZp6qS0hCEWJ/+iC+nd9AVJLjqtrSnE5kSEjrruSsjImbZH9b/QBlZJVZbUoKpDWXLXR
3OQTsn294piEsWAPySJvcGKDO82c0vNJq0GV9TuixYo/wJ+iBEFI7Yz7/TBmSHJdY1g+5gpPLu7J
Y/wGgnryWFYL14xzv17EvwACoWDoH+p2v4Dw1npb/dygZ7jgzbrL7u/xJtsfhUReWCKNP5iO0U7h
BAZoZuyn/IDAQ9mVFkUTnZ/Qx8kB8JNQEnpnBqL9K8LmulHHWRfuKGD/E4lS8cwVnofTTs5Zvcp6
KjjQ9BOEvHzIu+stqo5SCiIfRuafNLRE8wARWpoGlisLa+qZpiJaKUqycAJ1uFlcPnkOIcpcIODH
sODuq/T46e96WPA4GSz2SMu79lGXZbLXjNKbQ+k1gSO6E5PFLPN+zGxPd2vrSoMNndi2Kr+a39Bb
30Dv6DrlPbzSOrfOtep3FrgOJNAzfBY285P7f4nF+Ykla3b/T59xFdR1Lrpb05I8ye6rl4S4yKu/
3uvdylACK+zzQM+LNMVLPrWap57z+DJhy1W6PJ3SZIxRIL6q9QKd3y9t+JkGS541TleU0lfAGwzF
mXCF7QVxjSUHJY6QSFWFWYjIUP03pjg/P0VmkshIJJFuQ3HlGf5Nyfsy6Ok6xg7PJtuo9PGY6TzY
p4NXvWhlIzhs64h4+Z/64LfWmOLFbh+8668rfY0LaPabxKmngLycEKUX9kO4u+Zx3gC5U7iUvw7T
zEXiR3IK0TQPJkMBro7kz8nipdJyeictNZp0ItmDpVfEfPGqCeQLDb1h7snV2PNYHi32Eteblh70
/3mWlsylkYIGxax2cDPEG4RU7RSkRJ3oQXQRYwoDDCGlAx9aV++RI+A3q5xjSLcEFPJPGnUE5ATh
wqYhnw/LhZ3t89e7InnoZwTR/edmWeJ0KOxdB9+aBdoZrlAv0Ss2F9DdVOwbrQJ8qKBlptexBSbk
9jtej7Vxb8Rdl3QTPK18Z8NUfNKeesX7E5xQgJw+lLuCPhEVD2PAMol1j4O1XS0MhGaTdz5RnYcI
PLlVyAugO2S/lu9SxCKYKgF7sJOGTs0MBAM4+gY1QljMkgpl8l5Luh/skhT5AXSQugx2rDuL0Vu9
FlqK9xO7cWPXAgEbaecFAnAbCbtNOBTKVf3pyO8u/yhnhlnB5NAyw9cklFLd1Gn4qvnzNRSbKUDF
kq78Te2gjst33WvJG1ofU87XDDcYHEUROvvOi/7SGztEoU9LbXS7DuVGCV4XysUOMqf9nLeUTZ0+
0uDnGXFXh2s392n5zBBdI59ifuhHMc5GlNTrUxSSLJnnHPTryO/C3YG0OrgnUSvSLWeviZMp9j27
kEHvCi0MRtFZIkewRmnE1xSkv9A7rtziycfR2lCmjvqNLLOSFEihYf/A8JrrHdL1ZrwGpUqAsnPd
4pbsknroH6U28b36YmsksBDebjTDHCGgJYTkeOewO2ehjk1EP37zE+ZeIJBSmKF+1F4wv22qiU8h
FzMYhIKuZYNW58Gqf45WZfyvqoXX4RnOf3gqWzq0foxDHYZ69C/JSmjM4g9Dt0P1lz8WKnfX2UlV
2EFeQKSdj2icFI+l9lY/DJZ2FMq3m3s2Po7USQu7scGhu85eKR2VeEkXnrRUrhQKl7zXGW0APH2W
QN46SAO0LzlYNXq7S1O1Nt7B9QqaxFpqbO5vBQcqHVkLgm76qaklGg5dwB5bNf4le1pnUZXSdKf/
y8yLdG738m4qqfsHvm9ZNcXwKyuQnXhP+LH7Qlg7Zrxoaf5G6KJ3o4s240lpMZnKPoDjUUP3r6A6
R1FKbIy2Zfl6Zq7ndFylBrlDdUxXLnSLc7iJ3aiIE7giAXEFRcqWsizeXyqYiJb46lnuhEdgYrVC
/kAFWGZQ/vxFXSuLryf9eUBa3SdLppq6l1M04ryvdkM/7eAefX1IKSTXe+GRTIQiemcY4VdenZ5v
y82QRiF61Olv5hOmZO0WSCXkEqIhicdpivfep6krRMQ1elWZ85SvryGf3McTgc2OlSvctbekyMms
dKXVukK5vT4CXjsstndxDhxwhC/NiZgW1+tdwA7+Bd8fc5a5cWsb4FLcV7RD/+ECepIPvWn5zzwi
a0spq64b3JCP8/T03z9AQKYq5jwlKlyVckrfIu7WE1P781whQBXHM5X8pSo0tdUg8mUqohC1BjhG
CIllhZ8rWRZ034LCcfV4yCG3z+q45mQgWn8DGuPWSUBDrWNC5VSCmtL3GEcwWSLVwHGQ6oB4w3wl
etw72WRAFdLXdiQw+fAdJ3C2GbgV+AfSXV7moaV/7hDTr1aX5/7FvcjHr+xjJqT6trtzuyFjgydC
xPBnyBUEHiVy3W0Lk/b6yrf6wPe3AK7IL3SFCL5j4+d78QUWMyPbFtoud8dgTUvKUta7Cnd0luOW
bN7c4R1Skk20p6s6DUof5gR3jJnk9i9b3g64E2YZNk6A/kvtIXao3Cxgkhzf5odXz1wRh43rXJTU
D5Tgh+phHClALpFrx2OgO6qSTu9kIfFQ/bDvMEcLj9LofazSeTWqgJvuVrsX7F4Oz7COELfF3L18
Nqj3LBeHeTcTOGVmqdMCaV8uCmBa1O3/ikZ+Jx5mRKLEzEeGI5ADwLaPqyWI3JCs8izhSUCwfNxe
VZz6RdRlTOnkqyJmceAjR2GdtpGVKspz5gu9w9IAS+VPoeBrdaRnmsUOMN6HqKKQ0eBmfv31VZdR
NmcxmeBf1XskmIQ9NxJRev8Xp6ZBTQYPJbVfOGgL5JmLU/rpc8nZ2jru/RG7snwdKaxbR5EYKt2y
eapvgFyy74/KEO7tj9Nbq9dO0l4+W4CJGs50va2qopunfQNZEanJa3BbiJyllj87QIQgtp91yaRn
Y/f1Jj3zkh4BnV7RMuhrb8Ch/BY5xh90jnKjopBbeJ2o5sKc3+mqExo5CumKCidtm0SnUIO0kEoB
5ficOXDFBAOcIUFsMT1RyV56AaPr7TJGPfVYdqtRIOK3RxFFj4Umbk3K8kIbAleeEjAJqleLHI/l
9U47lJWlraUF/5M+p3oP1IA1iHvScEJoTuMI1Ie1LA854enbdEpHf48tfGbCoIM54Qq8Ao/kuuQA
HFHhezRNOrh18ClfKg+38VZP//0Qeegd0SciBmwq4+O6HGbgLm44bAn+Lc3EG1M2SmRF4VlhVBxO
KNwOtz7o2Dw4tvn5IypmbvsyvY/eC9IMfg8yewHQ4c2q3IH1QqJZsZ4dcl0cGAe1yEjBDNAkXdym
zD41JLuKUNBXXY3ZeYiyQGsKxyBhwpHNdpayKv2OhXatyO2HsnSCn2+y91x/rouyHtV5is8ggv5m
j7TnpCuebVS+x6z5shgerGzAw75a0UjgJ4vggf9z0LzA4kSt2b6FliO2pNDq7j06L+u/4pScxX2w
cTAN65ITmqegN+0EgedMKe25SZwDgZneXu7IazO4iyiP1kPi8KVihJ5reytPQLocWUVOcDTBu37L
U58BRRQI+kJqt/it3k//VjJBcshT/4Zo3hAXRzGunRQWI8lIEgpyjwDi+Ze0+0EcqdkINwFrxU5n
m38r+xzef8I8dJTfQVezORhffMAW1AH1jyJ80wKKlQl6wn61mZZCOOB0za1coms4hsH80fWb/Kw3
WGuqRVWmgcGZHRGsRLj7km1cnph2MA9izh1pLLW4VA5f8HIJZSE/VnubA1WuikndYbJ1kq1EPpSW
gAh17qMyqVTIHWynqxDDC4zbPlWQDWP2Xr7JNhOKO59oglTVeUKE97ffJthG8umb2KDovJpcA/tV
vY0pDeA8a9BrO3/+3JBw7TN8InYY8VTm7SsG2IQTM8UIj/NUV9gb9JsIH0RVLBnsOrjnhFRMaFR0
BkBTk63se4IUptBVY/6COKz5s/bnkWYDkQZ/Y7+Aq1XR4JiEb790YE//M3nKprhU5FQZ97K5QKs0
T5fGauAt6l1M6faxTzKlO38pxROMqUHpuSdnjSm4GsegmvOmD+/ZIksonaYx1J3psV3MfMTKynSU
sMt4krEUSFoFQ7WMMW0WSw5t9GoOeIoSNz07s62rDqhXkYustsMUItVCR4OUvLRpcUXmVNquiEPS
iwCbfKErrW6gOQU2JLEHsNmVajm+CXeSC6gYfQo1nNiROS9at5FdDVEZtqzwWIZO4USJn6npwRG8
xVlJA+9lL3eq+b257jPH02GSL2Hfh9SdWWLA7uD9cCuzW8kteGPkWXSVmjjskiUyTMlnoCpqyPx6
E7fS2w4jca0Xy9KWj185mFkkfEENh3yOrKIdzEc6HRfH10SaN3tR4RW8t+rpDBeTbzsZsaSkWTdy
XqOeISC11EhKjx+congwOgV2HgyahIiGC2wDrJMYRdcNYI6h8aK+tyRxOKc7DlFVaHRUBQqeK+CR
GHF5ex7T9eZZJYNcI2U7/nOM6DNn9V4ZwpURp7B/5IB2SHVYi/Q2zcM/9RKxUVl4OEIr3wYhk9Lq
WVg6pD5MwrNN2DBP8JRuuTBoH1PJyzYWGsf8eAQSkNADvG8JEogJN+2CbXelPTTfO+CMhqUZzbfZ
Ayci+wOYw3JEELAD5yQje4SgG4zqlX+t6p0jyK/1ofzU9Y/CRcPtRXhW4p9/ifsXR4s3wA+IU5LR
iL0jWR0QHleJyCjYmIy+Ziy4i+Hs3unPAd9Wy3EorCcqI2/AdkGG9es40S2TjVo/uD9lD+8kA94a
4jBNNz+TQj8MRmD8T3KrxDm9skCKkj3cZuITGx0V6WzB3oxgLTf82SswUnsyLeNeIg/WuXmmNCnt
ywzBSwJCfHDlkSMDb9KWKuoSkdTR31uBeoTfDhYLwK1z0aOkWlkwLmdFr7AbklrbhZg7VgFRZcjJ
PaVRnZY9KA7FErtYS2mhkHOKuM2nAJ6DaqBh6MQ4hVn+0LnFME6gyLaXKDby3yYY0Da2AZF/Qvrp
hofLzS4SL0i+/SJKEu/LzFKM+CE8P4JJsABhKfCUuDHpV2UFmu/nddxdcJ2lHj0Cy1EaQ+6ZNnv1
5zmWtaZBoIYbBW8drXPpZTIcUvBdxg4WheofemntIfQ8OlXhBHtpMjFXHj4ZToyUGm2cYqbluogI
6sHRp+ULFog2LDCGMA3wjknCE9gI1ueJiQPmAXO4XefCKMBd9AIXgrYe6/Zz3+diSBn/3p9SD0JI
E/EH7Q3KOck4hAMfOaktIkcJzB/h92sEyIOWig6Ej50D5Pq1cJnLjotXMcnZXyKKrEDBdRZAoPS0
pLNYQ6lqMR2tRYzaA0AOtm1znzucOoIPiemSXAmErk7Ox/qvRnEdO+a+UUTnMF3iAfuaSawaXY+N
idOemoINbuNNYftyMaw3qOcdM3PPifYHGMoDWv31k1kZPYs9tHWP7q2qvm4pS91KuS519mfG3Mcs
hYUe5PV3jOVkoUv7CHRC3uyv+8ii6aEYUfmEky525joCOuBw7yWoanaPHxxt6Fdq1eza5I/2W2V/
WDzWSl+Du++bq8D8hlB/Uf77ZAEl8h2p3KvLwfXBzwLYykQKNVSl//rkyw0Qw2+fiz6TMD7q5A26
4B/uI+Qf4WFFi0IvSP2NoULed2UIHZK1c5vVlL2d7IxzESWa2m+4teQBuIVcZ1lpVwd1K/O5NFy5
dpWfSb/8yTnFjfuza7520Mr7JB+UD26AHVqoNTWCtJEdqqWsF2SKdnuJmYjegEBW2kzgeggrNusq
TohKtmSG1JFO2gGD6fMACqllwPVNwf9apQgG4jfElJYgsKY+DEDnavhLx3Cmn9s2tS35N7qfZ2b6
oIa4YoKhVI7T8WHkX3P0K4fVpkSplg3J10hP+4vTtcEvOhEWy3dr8SFptxkcmHdW2b1FgTM7xQgC
zgwHstku/dmc0pP5PoE4/P2aIH9G3zVUFqA3qG3WW7M9ebTOhPQdspesdnGjVEL7wzYf+ldmPO6/
o7x4IWaJBrVxfzWeule8ZEkPQQwDmBZ2CviYp6NfMTGODQ71W35iFyv8PXvyoSiSgEPTsglreCzb
K2eQldX7m2bVUlRMgiHHJKo4rO/ADZtDtffDxZehXya51RqUrSCs9BIdY6+8dNyzUb4c24mX9emT
ygyKWv+6k7ShuSXdhhbi1+9V1ZW+Q0AHkmGDMD4R315ooTSzFXnBeYp/DYdQe6RZhUGL2QkzjcHF
jg5Gom91IGq7R5SYj/2euEupu1gvA/3HqTZLQUKqQJr6mLU78vb7BQ0LRGaO4KkJ0JVn3J2SMhUg
Gw0klnl4UjiEbdk8N+D4Cylx7VjfTIsTRv9lkFHepQGFqasCx9ac2EwQI4kmOd4cojwOqWeHnK/U
SgHhsPdkJUJgaqPKNpSzmCcYjhWsWSZOyqBv+SB0Wgq+rp2oSJHMJIhz1gHkfXaSWNqQoIxRnygF
n4YoiIyk3n+DhbRFQzTNfCEbi/P+vAxJVP7vUIY45GLc7NrsZt8Fp06MaIGhFdAy6GJj0q6p6Uj3
t6MKeG/2G9ItTO6FWYSNp46AfBzVvl1fr0Rw9cZaIA6vh4tSF5KpURGBQkVteSTf2IEG4VzOMLoZ
LktrSyghG5aRzeZnSidGuSHqUkI+vMAbd5PAV4uVSf9QbQvK6oQZSQ+uXR2hf7TR/EXkBR9iV5kW
EdChvDeqXMJQIK3XShU7uh2Gl41fMjHWKjVwmrV47uXO72OBTq8H3iFZ7kk1Q3y0lHOX+m9zC59K
nzkXxbO57GSR8N5DlKD48LZANnsBLix3Rxuc7ExC6sfz1dj2lm3AyeBZ6hnRV0uhTTNvb6ZYDk72
4IJlWlhK4zTgv4wfrZ8go5jhiWhTc4Z+LukuxXXR8UF1YnAC3ji1dUDfyzpqs7z38RC82QbRjPDm
nxf/qhC4Gld05iWbMd2+S62s+NONzagwKrtZbDmmeLjckKQgbz8VgapQojQAq5ZGdxekk5v3lsEN
hI32QKLAAUCTuwkC6SHg8W9wTknycB2YbYCGa7kVHwCaoqqcREdk+OKYf20866GqJMD0dBDe7Iht
u4fLRMO30FsAHYpm0hgc/jAVgJlitQsRkMm5RTdLiiZo9nxkIvEZojXr7+plmD85RTkMttT1laAb
Ivg+R6Ud31AJtLcbfOzMDCFalYiQ/cR6paudW/t4Ps3hd8SmiHK4r2jDWWo3lX5bDGQeg+Md0obE
SL+nWRgHcFBW8MpMUMeEVFpTlYehPjB5eSVaHBdV31Rzjih23+FRd0qPVc2iC/FpKHEBjyzsZaBX
tpqBwjN7Kjpd34VI13PngVi2YF+ZahOi5+bUF9onB3/JKOwe3bX56/akD1yPDLDCMZS9lWex/e8J
18OqZ9FVDvP8Ya2jb0iAem48eOMqrcteDHxQSD3Aqlu67zAiwUPQ/SAZkibDAPcgBqVZhnMRVScr
mFYmncfEg08YcAuHUmCt08ozN03sHcxq2CZYGaafcn2AMOatQHnplJBizthgRcau4eaqHzvjb7Zm
dSn6KViMpmJ3R+Q9vDeMLeq2sXagIL3Q1IwEh6uqwqObIIDe5Gkvr/lgVuDz06nLZJ1DamI2hSp9
CDn0bfupLumi0fl72pA1ur4obqoamrNLi55bgc5wZSIRmtbb5E2GvY1ODLFpiqpHrhKDYwodygp6
dPK6GOX0i0FnnP60YFSJa6CD9aR7pqHJPHNmSwc/jTtdcjIu8AabZWVstwSp2t8Io8dwMK8gmDNl
XvgMCtnu7iOK+spl0/Ltu8KIFDdFnZGufNuFXoq01BXEa3r7kM9K9Qf4Ei2yw8O04cy/ViFcJ0HZ
oVS9a+eEPY0r+JDJZET9eJp/v7hNVjBSc6rrxFs3y3gEml0UzNRh7vTSN8Dv79mviKkkMhRB1wHj
wu4sxQJ7yDiTzfZGdSVtlEhkz4SdPJ8vsUHj3/6XXeEWrkXPk/beverbNeZA3GFYwcgc4yP8bWBP
Y/htWPco+YTDlh2Dt6G54r0+vBrtpHFIk1XZfGSlKBDpfh+THwvvv95f6Q53atai8DHMs0MSKLS/
A6lHlbMIgYBYR3r20rdLMwz2jPOovkTYFsvimTrLl4rAqdY1c2M3U/YoLCq5iAK9Wd67asJiX4fX
h6n5QnOfJgsO9R3laMRsGi7/w8H4aQXCVnkqxdUZRwiM7zeLc12cth62aFDBlXSdFlhMMdMOWB69
GYhxMCcrHo3pI7cSSR4u+PfR11f+cDwyLvg+ScIqCP/5QaoH65aEpUJ0tD/oKonvU/FcQLSPgVYe
7yvohCquz2AwoarEHWRkm6FxOFSONYIYApvpmpA6R5swpy8+HF2uyVckneCpO6lX79L28+Npmkmc
il1XGBkl2t6b92sGVn624/XLmnbX99l6MC4C6z6d8AMrb9Pzh2r6mPp+DVU/YD2dWKRe4phlv+lS
anNIdNXKqDguIyN6CVXJOk2SNQkKZMmZuUysw/3iP4zvaB7pZZkzUs3yB89Nr0EZUUnw3p4lAhFq
noXxcTx6O9X93LDqWQRiv8FXNchLCF2/6xw14jMSPRyvAQLmc9ySE3I5LD9pa0CW1TjaSwz7C9Mj
O7f5YRpNKv67QpCL59jBHnoRJobD00rGmQWW2Dm+EX3NLcGY7JTRwge5FxT1nLiIAilQB1Lg/ONL
pWsfcD5MYrh3yoPmh1WPu6TJCW/OcIHYEfda0Dz/4pW8xiHRloF30SrREEl9oBcdNPdo8H+p0ZLv
JvNs4WQ3gVNkWIxbuYVW8eeI97tkJybSzVn9Cz2YN6kjvXbMjl5kPfJZwXwVAwf0Sn7JWupCOrMJ
cvLNV5yFZuzX8RYDFSn3g0EyrH7EvB1oG69X6nQYq29PB7yB1EnVc8mDqrg6fw42WIs4jlDjosfa
udAPnY7nUC6bQVCbkdl+SwjcGg/ER6sVsj3neKuMeDnSkz+IT4XZ6WuyzPh+pJXELSS6lC0pl4n0
dDeXjOqKFlTihj8gxROdzPlGBxlidIR6dvGLBKFSjDO+UQtacXwVjGuk5z0LrVnxMLv1NMR9iHD8
nB7vYWmEiGB0SyjlHJhIQnQwKFD7egEXHpd7sDjTkwNxiLBxVtrwc0bo1KzyY8U7DssaW1jlq10k
geqgDUc72pb6YlKF5HfNfmAl9EUNjs/J2HPVwmWSQviPD8vUR2if0IVc8b7UbSze0CKOMGe1mqDg
qf6nWBySJHxkP4iPCH/nKKBq000fhFxkzyhm14qt5dQ1qLD9BZo9rH2JA5SrTOvZOf9YdyNifaX3
MlSLelqATzasec0QkiCZjE6cIvtlgny1snmjgTny5hGIznuBzyyrVFC+O7aJGU0mlCQNaVot8mn+
HPflGhxmN+P1eQSBqaU4Pkla06QlCtWWIn7k5B7BI9nBQIYWbWa1awBzQ6ukcCq8LC7vJv+kkb9v
5hmUlB/oXH1Aa3m7MP8R04ArTSlBkMXqhJo4YptnS1IqmRkIxT1stqOKpoKJsI7fBSO86fO3DXqw
fGe7gvTR9wWLLaeRNO7iDmV2iS2dYTIy03jReyX/1OUr+fTyPqgWNdrCZBgIgx/VIt0hTq4gyeZO
A4HeYdfYKljEmS8SWKOKHniVdbR2TJhmGRXYX5ZJL+3fz/CWRecLJOMLeriRNWqdwxNiZYpX1tmj
dqctpXUrQp5cZatMZTwIadlWxi3Gb5yEwQYmdmNsPYYFaq/2JoP2xgHw8A470JaRi4pPwSHGDp2E
wh9f+FTesZHuBrIrkX+muVwoxlz8BgtBpZxKLh9oUY9jkqcSlBoqL4HpNqvRIUFu9BZ5QbK3/iuG
DcMdMNEmeu02JRV6JA8Am+H0i48LK6+RVCPLQW0i7NPvRooKri8bvidmQKGRezWVNSRGnntm5Jxl
kdyK8HSF+xrJ+GqVSb0btEVPwAXfOA9sq5PY0usFI7hrODtzvH5hMmgMbrsoffI33csVzIGFc+4x
4/RAEYe91avt3IiHqGPBFUWdruu5KXxaTMRUkcm4hyKPqvQ+JH9PsySdzCDFpl1jjNUVor5iFO03
cnLlb33QnR0q70Si8KiY2IJNiObV2rK87B1Oc+fgmpkOFLLZhU019tz5YKFpYgmfMVY9Lo0W7Emx
BKoWEMuT8G2NqzYkA1EkTQ9kVSDm4UYA8pZaqCRgZBwV4yGC9/hQ9I6RGBvnWw8Lbjzh0wNPSNhv
Mweic7omqkQ18Ec19H47Vp2y4/zsaA/eaiDGMTx+4OCshlQqWHzqrVMVMWjGIs1ZHxCl52FCkM1m
TiPVYnlPrSHoRLHpbPabM6ptIpdB/WZRPcPh9FUFvZ10R+I3S22nSw+RJRYDHpZvx88tTdbzmO8D
EtLKNTaQKmhjaRqldeCo15s2xuPQpfFwBAez9yFlwYKdOIxtl3hZo1CuNw3UzXN0K7CDAdtvTweV
L6sMz/rSgBqnod0MlphCU+hoT1dPxwtKMXFwjlKLxIIKyYS0f1tGd4XsTzXNcOw36PMQT4P+aSco
sYv3oNZ4GZi2uVjSgguGAq7wwcEIHZe14ZERlN4h1c8NoX0XUFUVneXhJc8943XqLHA7pI+3FxwB
0CmOPL94pAs5TwxChvwiEpYw9dhaHAACQj7CVN/q8b6NEGNBTHbxms1YHBDfPBroRnI4rcZApXH6
NYmiPXClghe7lbCGHsNJ71OT0liSj1I51CLuoBBzEfARPdVdDUZiwr8v035yjJnlcepN8eC/E7JR
tfubaTEpCm6S4p2osWZhZ/YQEoBukAfLz+QbnihqDwvywYcOgiY6cOwhEweBMOQH4DpwrXutVnV1
KSLd0cvbyFth9defMKAxLM6vSkWm9TzubpOBLRThcAdeq41uQSvWglxadAYZ1PNiiMI/A1zpF/FF
VBa/2BqkTVUK/jXfqdMJy/54IYVubI5OW7lUp1/5xAgf99N0L2o0e3HQrjyRdhe+LaxxJ7mcfWJA
trsQNZMAYz3R27HO+/8k6ky+glTHKwuwrOGudNHc6O+ugDGQQYgYuS/2xI5d6gDWMZuHyuaussW7
uGoD9hBXgdNvgfg+bEOo4NtRpJJ5MhMgC5zpe/3c8cBGbQdj6+yj913La/r4iILwa0Zo6KjEj/Qz
2a/oRzwhFSWKKkovN1PmTZP3L2ZUGzsFz/9/bfTRzeCHSNzbAZpDwsZsdAXKUNhZluUHQEQzG9f2
mycjVq3aV8MiTSFoVx2DWW08Ot5G90xt9M+g2KAyQLCGHtF3ql6cli+r9ROwhRNt5osd7xKVwXzo
J4CXp+Y+TztquQlpD2MUkkwZgOFXUn1luChhtX+E8DqtG+aeV8txWGA1v/OnbH8jMdh8GUAMpb3H
WIa1+bZPdEsLt/1YlExgP6ZussefXa474C+qgewSGkb+DmTzM19Y0IrYr0YV1FhUmWuFtgkqD2RD
6Vxcn3LdrtAyW1SeVVlVuN1d/7QFcmDuWzhJq15ucmosR0tfWRh1faCUlT3H56/2b5dQOx8lWUz6
N6nt4IdknhG+C28bskHMVC50Ee+jkxXsTRpnAZ2hhDFleSyonGGjMyWS6fbXj/ZOs1ZRxieXFiDh
cIwYWL6ImsvzVS+kFZCCMhynUPXdR9RNEDxlctFrxn9sbIDINHuauNICm7JASyMGFEBhvXn6Cydv
oN82Q6mFuYvnuK662W3Ngr95f5ZNq/6b5hN993e5lrhGzOgENN6dpgMtu1jdH4tYbE65vkAtS8vZ
yXm+CmfKeOZzFh+aTexS9UjyrZnZ1rw83KprtleNXW6rUYYVViBkmOGnX0a9prKb7tqMeUaor9ul
VeljxHDDRvk0ELAy6MQopHxmplMvzYSw9mMBBoyPEtTS2aFkEcLyxz6hvmKzlQCRgY3xgIvvxXSp
D7HiQROYghekGoguEtRVqGr+QOoIZWJ2pkcvGI/fQadloWUMgzRv9p2mnFvwWW52n99Z4XuxYWqZ
U20Qn56ldeTMMKam7fqC6xXAqe/pjSn8gSkZa/bZORO/ZmOrPXaoPgQhv3O4STXb5Z9+6yXnfAb6
w0wN8tUYt/NbJ8br2ESmQU8UFOK/YpARlJuNkiNwcQyNZpGxo/noMKlrcbgbv1nqoOv7NSqG+Jvn
5Iy3mf8FSeXUei0lz+8wu3TI8uOeS2LhdXZTvJqKxlrVGS9Hq2fIHF7FcVIyYl+Vms6NreeL13aE
UGxxom5VluWGFGMg+16a03eItp3+s9R+BlmkeTLe83AB2hSBacY3bdErTSmPrnUlnODYtTTsUp81
5mNGEE4hPbBgytqOIRDkegdERRzdtjI5Us603xDTmGZcof5FmUR5OYBXXFxtXCSZz8SjXGlVfA4c
+yIeg29/8yWNEx/Dy5RLc/4PYNClmpT4Y5ptg2BDa9KcnZ6ryO4BkjHMExV0KZrRh7StsRyX78w3
47cKoo7byStVhj1u+AkUEzgbE2LuMMkdl/MjS44Kt7Kua3z2gYSfGaCcQaFdFkOhO2FbCuxjoJR4
FJY6lqz9pMUDvU1joaZH/XXWy9KFmaWc1ZPz1NVarsVfdiKrL7P7T3QYGD6Ea5B0zDtHNUsNPGfR
OvrrrOedIx5mWdTs+veCtSotQZ2GiOuFo5EBWNQWiqbyslfIhI8AtHZmSmDArlhgqRe0FrgIVDKP
2O/yGS6gBHKK/ECy+qRO32ZlqZAEbWza/C5JjwXgWzI54SGgP5abHzvrz6O2Qx0Bnsju55Q+EWJ7
yNgEPcTZdLgk2IiakzpK0SZ3n7TRA9jjbVKzjCfxkWfAgdJZVPJbH+ntiKTlEAvxKXfyACYHdmjN
1GkMd2gkR0ObO/5vcnGiOaSwy6jDnGf4wnHrharGAYMuGMOSxuiIxox3cjC3osaEOaPkz3F0rhNW
RyomGq2zZAn0fWwbZFt7zuCwJioKuWxhcJABPNfoM+VhLO8tenR81/yIMBMIaJRkR8TwKRI7JZ1c
GalDJFMGiZ/de7DITDa5yvPq593WDJeWf9qLunMDaFfKYGvVzBx8Yx/Qro7FzVpsQ4CXUg+JlC9B
0hneMc3UHvhqLHDLOTgniOd9r7UQtCe3186N6e+JAD2kII6k/+AkZyArb1ozvnW+tCc0VXfhVc0Q
ItAqjLiq8IOqE5vFGrmTwXQnB6U2V6uLoUuAup8hXSBjmKAvRa10ryEsx1Qxm3r/DBLs3QYum7EX
WN/a5oEJ1LmufcrQzwq5Qr+lFxtireIhB+p1SP5Q9el84A9or7YkcptrY8TQJ8q1eIXlgDhihjnk
75Vr1qMeDUT71102rh2NO9Ebv5JKsGK/scfPheLmFZ0z0AanO/JAmAWhtep+1HcukWZKCq2bxcnq
u83P4nxIJlcPyHDpEQWQG6iNSmcUCFFCKi0Wye017gVnIbG9RXdeals9dZg0RxoWWo7cYaUN7qy+
Wt1de+3buvI4D9hR8ZG7BFTJn4s3EkdMR0j+q+VKHKDlykgXJe0NYBH7PuK7LArFZBdcAZjpu7nh
nE59Fxh3GLzAlOUwyXOC9oeuuMFGQWOjK+tPgnLZRUTPhxrssXvyKEeanFUwKd+ODoFtzugAWtO4
ecxl5iQ+dHlPJwC7iMyhAzoZN6MkbTCgjdhp/UfseDSPNKiU4rubgzyUWPLKMvRXmUBWfZmfYh29
EzeHBXduDGUtjL7Jlkcb2vYe6h34jIWTDPEmNmWKBbJZfjlBBqUv1QEZw3/Auymu+8vzrLTibbH+
9EKOiqun7S9rTUmytn2l94a0LcVKSHZXJbZAqFw2qgeO5oKCJjyU1I+ZD6RCpZSKADotCI72AUJe
3D1JtPLHBp82AmROz5DK6kZc3EKfzU52ah7TEAO5PNU2ckxqv48o89fCBC1ORrBf9G8sD2SfTbuo
vFZirCWdtvfd0TGnVlx6hKDf0Xj1L890iiFc9+P/XpFYz2KW07vfAv1dNn/jFmWh5jmV8/1u4Ni0
d319hAzUzpijQI71wV7hMT3vNNP/xOXOd78VUGKnTSBZ5lsAfw4jZJr1JqdhLp+1FIg4PQOqvOZ1
CKowT4y1aCclwkz+AQkHKJPBRLzW7GFWSaq1ZFGCReQCDCl4YkMpVS2Gu1fmvo5/h+RMCI/EuAXn
MToO/iu7W1fjm/NwRafs6fwwAh/cRDTq/POzmPLmNHGtPogYVC8p2ZG9xKXYBWIBd8U2hpAULXfn
1rIthBNDkgWutgF45rZLT8jmP7SACoMmyCz8jGiFHLF5FdOFq/mju2ysKquOCzNM7mXz6jtqrC4X
mlqRXas4YA0tb2rIhQ2jUPy5FT3KENoHAkU/JOpTUDDpu8V+AxVV6XZYtHlhMHX8bpc6sQXrQoI4
+rPNAQAt8EceUjmR+AkK7h/0pE4lMFD54iMAeBOuVuLGVOLNx81qWn45IQzRQYCh7jtJAb1F4w/l
IR8gFGSDk6FMTrL2yJKfYGLwkfQ7zdPEZzFknHW/zX8e6PAISLLQ04o300c+iPO8XRKiVWVSp/f6
qSKF0Kk1wjScB/QO4WwKF+qRjMEST+3bUSfhCrULbH1aTjOdvivuc2L/qwOTYk4eNugDh7OagYEO
/jlLLR4Sk+u9BWKODpLFJ+ADP8P8brUPo4mIHkwIt8JpsqoeDnYUYrq6Re0HmSKzMubm9ifLSX3O
cIy91XH3AbEQJPKetlJhFO3LaS4qKDCPvdTB3uCD+AIeUO+aiOMDQy98qjbdF3pZ9XDNAMCSARoh
sSgRJYCvy0PgNOKgzjkNjF4auaGID2fDTcrpnZTbKlVkuO/mtbvXW/q6wM5MDtP/NKk3As0Mmq+o
xErNbjjBQwZTW0Tb25q1JlJAPzSEiAhFAZTOefj3ID5Nec/QjNoPHp4JS9nglL96kbxZf8n1gnxA
C1cwilbedlb0F4iYwgtwBixVfUJAihLYG0PbDmXmFrOdo+Wax/KdupzxfeTrfaVGse/jZrb9ORoN
ZfQmfSlBZmw0zBCDNqqV7wlPvPNqccWWtER4fH3r0d5gSs0WOzLceGZ8x7rYS+LsDzpTtr91OmLk
vZT531T3kJFwdH9O1djQhmf7f1r1EnNkIqVxoQ9TuCRRnzcQQq20U1y8TCRcKNnHDnijFpzvIxE8
cOKGYyaE0yU/Ay8iigE0ZF97C3vNH8ddRVV5zrluWxIdfRSaKvrQUF/e56c6A9Gm+MTP7aIiCiFx
JO1TMtrtamdt3xIomRrr2C92TwRUM9hF8vtWvgTAqWJ14YU5YHicf2RdBpNN1EiYh/MKg+Cr+0Gr
xnwK8YgQltboZZ0fOOzz+m+CQI9gVDhFvSrc93vd+4CGTMk7qf4Tc/2pSKrmMFQD9aXiTO5sbrMk
5dPdK7k8IGGz9AsdIu4uyHKx0jghi2AsWlssCFIJm7B2TC72WgyL5deSTm25EUh175XymKDYdKR4
I59EcUArKMS+AOUMsaDn4vi/LpNU9L6laWnoSXRrtyEB7PG4BNBMHjxjCh3jGoJvFyfpjE56GiWt
UmQZuCewW8BMKXDunIPUOkC82AJBQIL5kxNoXlPc9xgF0VaOkLkleYyoN+LfGqmmOUKrVHty+fKg
TwNr5SUx3eM6fHqblfA49DkyqKAUoaM/vLNNilobE7KD3KmhbN7qCTt+u/ri1BkPZzqE+uca3Zhe
89+lysS4JXSAZb5uOV05BIXmkgF5U41XirnYA9Jymrs0n1ZhRBjemj6yE1j4m6VgGsBxqu+Ki/uW
JJm2vEQoj2uzJ7ImyL8mX9UYhQrtBmta5U+2DihjpCVU4dCWhklVS0wy6ll59WKx+4Kg3TM828cb
sDhOHfLIuIK3hz/6rZf/2bBi1/nLfQWVaxmc0Nz4xUXTmk8r8SNODWjsucOx3wSODI6Bwodl8zvW
7vXfr3j30lbwQcL5yw4Vw7e7fnABmuBLSPCKPpq2wU0DEVmehGhp/IvY/5C2GMHij9V5MxhK7k6t
kyU+mgLviq/yQEgeDYR20NUMlZR+F+Br+IuULPtuhlFfgXzHAzk1MXINeEf5IsGIDRhz2uanAsS5
o4rIEa19gWq6Okvt0b6IsOyYYltFuFL1kd8jTpGbN2CJlesJnL/oiHFoiFwUkKrsiKuCexqq4fJK
g+k0dtTO3PPZmqNrSPzTfJirsqLInD1iEtb7yp56iHtX+/F3YoZoBMbDPW5PSIqsbbADYFQWKHVi
cnMDR3Dh9SJrlfzMBdner+KZx0hyly6OJ7Twx0fDKbVNVHahFgxTmOeWIJXXB15baJgsm5OyCbfH
YUseAqlB7wo+Plvf1yIKQmZKRrMG2nNLd+WxrQEkZGyI3AgI6lSDJnLDpKmn16bCN7nj3ljABpD5
tSUM3KZRm3a+N19eW5+hn7tOxrLWp3GMPlw9GmRmaiU2vH1dqdPgqqvKCz14kEyxNrBTBnr4E8nF
LT+LbqC4TsOwvDLpOZj4yoxhteUo49kcXDsTz2O0L/gvuAtHkHCEoYfWuS1I+BUVV1MXsJs4MXoW
LMJM19ClT80X3uhDxoQgdqgrx6eG0DX9/L9THUYuw4ie53pn0nOTLjISWLxhkD0mKLG7YoI0ReFU
k6nh/ac9go/cxVkvLJlgengZz9veB8m37Buu9SaiOX4Wbbjlbgy6RdANHIU+Pjq5RfizA44mUTjM
V64m5KLQ7skJmHrlSUKsqu+1Jn9WB8SPS+SRVUNLzVXvTnD8MvZCi4kcd3twyGktD2wqHStfoRLk
xhzS+YGSoB1crpFFqFFmUGD2l+ZHnFKxec/AqS/TaJ/jhCQOV4TObO/tEx5zqBZTqUMmHjZedbAu
k5dcmVzYSwdpMsn1EyHJOOY1jZANSSQwt4RxhivmCw5VqJ+Lh2jtWZZAKAQ4Wy5xBhg5nLINZ09b
t8jQ/npGgHBHsvpJKyhS7FfzoRQ4SoBB8B54fUZBizB0HRsTgCXJb8sEQJbmBbZPntWDH7CUmrtV
EM6EqiJvcnKh4du4IWnq0r9E3b+GfcJ/aErSizZiNXFB5Ffr/QKdx+f04uy45xg0aQl7vUbldNXJ
GL66JSCIq6obSFgokLTSX/H4LEBMZJdKdeHElIQhcedSodx6FCJ8cPeoi4qwXN6BGHHNbUrAuGJo
AlDDbEb3wxyWXXRbwqx2/Kdst4x7nm58Mzxl0tYvMCzdfFyf9XTaRoGNTWS0wrLb5cQJy5yenbTR
TMRrC5T+tyl55Bi69aL4QBCBtYeDVd3V1sgWWoGduRrXPUlmgZKIrXeoY0LQ5EZKtvAzb4b1h31K
RmSNGp3ny4vXgdDwG9M9yUlBts8f4Dl/3QVNfXzLEgrKt4oyZr0H/6e3pd7jtu1oy0Nsf/GiOwq6
a8kMxw4vs8UyRu7SWyVJSyo5cvqMaPOrEVYFtKI1C2HDJyNniJ4sLaE9mFawqR4Frtlz4VlsWmbF
O0XVe3QB9y1CbXCUfETGqFet8sPbqTk1XOlvJ1nAnGh53Q77Aom7swyA36NiQlfj1s00eKwOTYLC
+B5KLNYtJGmSzcOA2rEQDbk1gpvn09skqspzII9YS8rDb0ED8e+b69d+6RXhlPgYAglnfkW+fEwI
t7EcFF9BvchV0HghmZRDX5OgKAcwIH2bWMXle0yU6ljj4C2ehFmVEGnInRAAieLyHqcx33gEle9F
ah1zdejyqNr6ALJCyEZ2MrivfGh73Mb2TqdLnh06ZQPhLrABUaN3FQFboCn+400SqIvgEe74WpfU
b+Swiok1gKWKfCT5JBbby0XyP4k4ih7o/Nznp6t6cdY1sMIPNcni1+3dAyHjNl5TeyGspRAo+MCk
Oa1Xl0XupY+JxN2AytXbNbOKLzSkoMURo3wkmDo4YgUo5POjjWBcw6fN6gpsbRqM3gnhJ2rtTG5Q
hNnd55M2JYFkKj21K79MSDfP87TnXphv18CFZN9fjENQxdUd8nSNzJC/VwkIPfR+Jis6t/Yp40SN
d/qT7pRsbm4yJld3p7tp+VptavwzcFWM2NcljNGykgs3iWBaEHps+0l5W0LbQTAUtiSUzh5juBLy
avZtcRLJK8MzLpKQCftHNT0PPzWP2o+GESFtwc424f4UDKQzDScVm7zoXnym/ztPnNrcDAGfwg3q
tAlsVkmySEJv8kDLTCCdHp29x+lI5S9Ak+pG3mexiZ9SJdjcogoFrSXOtashlt+oZHqdcSCWwljr
st+CpufLUbMG9+0x/sW+OzQAnlB7uDqIOEFDit0aivaC45Ip18AdJGZ/qJzFYIeMZskCuoEONutS
h86NnYwVR8dA/oY/Itdp+SBxevYhtGp4WItUsv7SZQCQztEgObDr0D3ZB2MNj099TGhKL+CG9oLQ
9iN1iwAu4R7zOdSwPAmif+0GyFZD7XvwdMYbFfi4q68E7F/TYfakMgHwe6feI2q/ruNqTUyXF9kn
0KsEWKR4DFu3i0f7RZwACXvFaCWOHT4fYdO54g0xJtw085MK5AV2s31IJ9KmeMvNLPgY7ibIJLn/
GtaDXJJEQ/TyYmDqB2OWXiMlJknQWBeQE92JfS6tpjwvrRQ1JybJJp3WaRZCFdW1urD/7AjiGUY1
vaXq2hUcCyjEnVhvOS8cYg4x+W2OzdBTqLVh2svYmn7zyyWyRAptO0kBrxd6K0vp0qSZ6HjmuLDP
ow2yKMxOFmLTEWSjm0NNIn/0jrV90hYIvzm8SRs1BGdArOzWsTWzCSIn4uyB2l5b7zWqFK9B4x05
LKhrhDEwy9ldIWbCDm+a+gQxiMRJCSOAGCGNPWn2HYURJqLIxFuM99hH7VtOJxXuVB/WVLKnKHw/
CosePdPFMHVn3uaHVzVYnAxOHxx7HrUyK9v0xRBWVQakeSB02txa/GqCWBLnR9Q/3iz4ID2r7Hxu
lBz3pRBFwf6OI6fEGwMMe6WhWNdPUH8ScKmjxVga6taQ1wcWCQ4hrMITnJEGiYlQdAjrOQV3+N9p
/QfeUgRlimSnnrn98jlB3a886C1PM82EJ3WbPKxmam05/rF0oG/V7/DmyfVTIKw3DsJ68pxGryQe
hdJYwb0vwPGX0CTNmli7yxqTodtyGFXnWoBT/AolhGcw0VmyTkJd+M7qq1r9Ugxdl7AK2gQ0xmlE
aVb5O6fiemt4XmcG58YwouZxu0eNglGkPq8Q7WYUYO+Oue3y9uSnySgJlQSOFbAvOEicabNAawN3
8AxrsxgcmANhlys8TFYo3ofkVQ7GFhXAS33z+Lam04KZxlf7BeVARGV1v7hcyaMaH6ubxJJUGwir
tTeCZHegSj8mIhsD+2p1mF3B3FfPYMxGIEx0v5KZtKZt2WLrfL+y1tA9nn4367vz+RtC7aWBv4lc
+9A6vHK6bw2BCgnKh2iA6KutScZSTJwol1SKjS7m2Vv4+9Ppcg57UuBFI2pADDScj29DpmprhpTY
ua8oVH7Zwcr1MGryMknz0fjrzlBSrYuYJKio4xVIhANBn1LEHlnrRZ4/80WuuBQnj7XRCnIEDAaj
sDB5u+a6Aym6o9I8qEPQ+p1hEgUr5EJAWbk33sBCehHsJWraztMQ/5Wp7lAZuaCeRdFIf4HQwZv+
aZp1jsDW8fNl+I1wyCjhCx9GUDDkRh9yX8MOKq0gndDod4qIcB20gT4HIl8S9p5mgVN9lIqmEUHk
uo9C9SPEm/7VNSGXKanKh9jDn4HdC0CdI7t8Q+J2HEFvlDpHSh5D2XuxhHNa4LgvR9O848d1/JOJ
IXDryDYOiRdyRxQM0uydO6CK/LrFRuQjSuOfUUMO3pkrow2GZQMudCE/7EfsG+FotvOULlw/wTNS
8jDfctXG6Cth6BdSo6P+GyslhmUdXmckncFxu1lnaXWRntG1uQboissxenyZCkIsOC/p75Po9jdm
WEY55lvRkdYBjlZCnx64vVkUdkMea8aravgDn1mi5f2ujfBkZsi6+hEQoaOaefWYWwfYHPwshHfl
/IMvI6A35yv7HioW0Xv6GLQ8t7+pzlSM4s2QgMA6bp2f+AVT0GpydPInLS5R5TwWjByYv2gnLGkj
7Ga322LSNnbCBc+MVfkg0gIC1J0XAy9R8cj3Y0XPwXaQkRU3oMnyxiWksytxCyH1hhTUu9NMsKib
KyPVtQKGVnqoC/eyNxw9a/M7gJID9vdqLRDS21jAqBHlXnRdAPQEMS5FSDblUqy5N3xDaWBpbO0V
T9aGEXk05OuQnCSI3dFJZ1f8/w3vMrHVZgdWuIJs7NHw0DwEbmpiZLWsLrwbeHHtlV5dKIkMz9vj
L6HIEYyU6nCVMBWp2hKAmrWhDcCoKQqdKDoKDYAgxIVgVe1eXCKP0Cakhgey77NV1oBgCcV/Caha
dD45s6jObXAoKjBf9DE+qTs1IvGmdsOJu+kez+/HnRvTFA/a5qQ0AYvCGPCRvkc1B+Cv+70MtWV4
0YXysORDhP392Cg/cPBN5N/mQeQnj38wFl0elltUdsUdAJmWpAPj6nIKMlDQ+s8HW+JkjvTBqVa9
jc4cXkITUy7vu1JNmWt+FMKKXxl07kCC/Eoj8heGm3VFWyDOgCKEBgBqTsvsQbLIlTJzYxc69AxE
SG/7h1Rvclgo4MAQxAo00AQ1+FqR7nPJK8Te50ZVQN0DnNdjz9VlOZwuKnW8oQzgZVVphoNmWoot
7zPBJ5wgW8vSERahCp8e5OqJW9pH7nCD3abVPlQxmohIUN+YTFlmsdXYxc4I1zpVOzmPN7CEuYLL
aHrgM0n/3O85WV5IIA6T1T4+d12YZyU0VJKs3iRfyPNq79chFuSeGjDhSy3i5JP/aCuD1mluJRKk
BmyNTiO1lxSK+GjW7Atr9qmxsSmdX185Bk/u6snzlg4mDr65BwcWMNuO7g3EYPWR0H7kvY86rOY+
FOLwFkbrg64FLwZHYgbnupw96i04B8s6HghLvn2prmkYB9jRhO9oKNNOPIxJTv2NwpK+1LiFATHD
wnseCvgFcltO31anf4fY7dTeaa6E1fg7t1w2mVmhS/Dfw4yB4ZrpsB0oYftYcXt603P5Qc+G7wjE
mVe0o/1fdearDp8zyBxTU3HRsfJ9pvQEroxiex3ZLCHQ6QDpslbBfST2t3a+hdW9sst1XKhpteHd
4i46QvI3tLVxii5bt5lyRTj7sQs/E+EKeN1vG6UtZAht4/4jJDQVVewGeWBW123wMlEffdZ8/9/X
8C5WDr0XbDtOKEhhYEHT2vsrihoElwFPKcBbg3Nor6Lef6dzfR5fnanRW7dIbTJWTi/LDAnisEy3
870PRWtWvETkGn5hUbEhOybM8WScyphgHV/6z2DtyfxdUNldkrsZTxvmionrE8d4XrLfprcOrMsG
hD/SC1TEJIhOifKmSjCua1oCSnKLUoeKDzisbFY41/rJAawnir/b15mRvINGFZY4/C5hNewZs6Xo
xZtF+LcehTZmm94AznPYdpJbXWY3Ott0DK3IZCWPF4RCm174t5F+fjPTNX6V91uy8b5SAu9veY2Z
a2u9HgItAWjqitDXt/7zmdnzThKiKWTwYuOQB7gtBB8N99ZTGgJ0Z7trAycAaIK8ZjcaHkce3pOT
FhP04SEhYJS0tDmNA8emrwdH0athLQ3L8wY0c9O6bOgFYMMRf+xViWLyF33SRg0qJJh/gyTfuGw9
EWhU9EgheURbI2eEqSKj2oEv3Pos8bjQTFUMb/xq+wwg4TPRg/6Tw/WuOWeS4y90perPF/yI9Gh8
fcu3hBD2t37/R8nfKvGyYsQ/QdpCttG5x+VN0ghowAVoSX8n7ZVVNlt63SiqiGXitofWsZ23qrOv
FL8BGB23LHxSEaIpX45PDhSI7NTy4Q0D2/tZJBQaJn/So7FfUPSy8Jvq7P6WPGO0aX0DAMODNHT8
XksB34kKrookROIOPBm08aXeppAoQx7rO1shU85NxPjP019/eDV5bOTN88S8VkNEp1HgNf2d6VlT
GgHuvDrn3vkAZgmyEGA6egiGA2evfKEiaelf+26UTRj5rISJOo4iiknomF+1ttUrvFF95fR8Ar4n
SuPgTgbGUwSEFJxDw7gPyxrDbJR9yTsslBud30YLui7keUl0faCpIDVaO56qWzXg/ZvCTUCl7JjU
XorMPVu32uzLBv6ONwHEI8J7uhROFkZ91r+B800/Pt5nESJAyTp3nUIBeqPUu6Z1qn8CWyEk2Eh1
t6BxzPDtwMpJov73hD/2/xEj38Q/QtbmOt64O+x2eWnZ+oBmhnoXlGkUEARfz80fp+Bw5J9agW/V
Tr/JLtXUFirmvqPwbZigfofdRHvK4q7K8yEtiII3zqltLgOFbPHHx2rt1wlW8dFI4p0CJpDPlqGh
65/Zj7B3fKmYkWqllfsVGMAmKj0eioNBneL5OOvclloTwtEf5V62NpGgD11RFcBNuYrWjFb9Mnac
7kETNqmUmjSEmNnJUrDrTKa2I+Oc7dsPRTD/hJHjFFbDg//ZpQ+uBEhJsj3nzGq54k7+MiKeDPdD
FLOhnoUiB6mqRUkodECMPBJEGvj4kQKZb4jJNPBjQ4hJxhdAYEzHXkvkBCo884DFn3ffg3YCP4nQ
YuJJoSF707XMxfPsyS6+8UM2frd6/RcXu6gaXhcWwysSnCiMLHlW046r7AqwwwXRqtFSmn5KwWvu
1fZAqJ9W8QOd89IzpYaI0o4wlQ4qHojXmiPJcPrmouAFCzJ+yUjuSEToLy2ywJj/BRFinQOQ6F4q
AUio2iZ27Uv4uJRttY+NEXDqbTrfhlIcS5O8WsxVaxXgMk4ogyeVKBvJdXEuxYUGQf9FSATxd/6I
QBNLxo04VtaQEQCMt6Kkbyn09bUkV9KxzeWre43bdH9a6AouHQFMUSRGrgiSveZcXqTT/0X9KyaA
sChfhqFqn/wvIXaGgSFb3yJNto4SNnQYz94mUdDkGdzj0z+C5BEebJXERjYGGCil3CpYkhWInJPS
N6/yKO2Tfj6GsZo/3bhlJmaUsCT2UVwZDRQHHtgnCQz1rekU8qlnuW/4NYSfIGVyassKLNI9kd74
Cfy9wdFo89zh739r1NYb4rETkb2Qa/f405VZsoZNvIYbUKy/mqh8x66DcXlcmYuAb4WugbBbbovC
tRCGlKkwSBSChT2sONNHQyDAe8jCLyMx97mLD8YPdP/M2zUBvoWgarhg8QP+PBlJRj0Oh8kcm7Fd
wv+0OHKPOAOI7T0q4AFL8ljKoN8FJm/4fHcfCW6nSCSLpyRmxBCf8zDf1O8t5u41RQDCPb1EdY+w
MDMO0hRE9zASe+orIwRBxVsraVXgVU+3rQj8/EpAzLgCWo+sajniRT8FgPA58rFWQFoO9FeadhOj
0/jWONCXYm0FbRfY94G2RL2d+p8JPqQ/FDIdHOjvPlBZZI0kvJb6rlRkkQJni9+kWpp3Ji/PS71e
bVJDwPwTfw3J+MPyW6dINCccu1/q7WgXqn4PkRTEFf8k+45J4mHDz6SvOjJh3OjtknMJ7dlcKTPf
UfzUnKER2ysUSjMxJnZRpskoC13cuKK4C+0H+SFgIMqgHUsPV8V6gw9+mOdaVicLmmLbJ/lKfLj/
F5xAitNcgiI9ihq085c61FLqctp3xkubOUqiMrynYpuywvv3f7j5Y59tb11qPuJff5ubff98d+/N
2BIjLltq8c7nGSI8NP5gzWn2NLNl1g8iu4argJ2Fwb+mX4A3ft++KpIyRNwjuDxIUBCTQwtPxXPY
KMZx7UZsSNUaA3IJtUQ327CgkQR6VTzXYI2h42heSlQ9Bcu+INfUxsig76E22vdvLISI3EDDAD3t
1M0e6hbdoHE93QE5LRGRWT+SQdrz6Y+lMKx22+gMWgasyub1uXxZXdFD2I9lvDcyZPqfiFIaY5nc
ixBB5S97oTc8gQIUZ3JgNkCNdiAyFWDeKQpnPKVRB9D/bmGBXYAeJP0tgUEB2OD4dtCeV3ZbxDMx
9jVaymnkFYI0nJ0eyn/0PIaiJNwUCG73tVIIW0UEqFD+Ve9uSvwMt05bDjFHGTj28QIIPTbZb5oW
tuU/Rv/iXmvWeaZjBKzfOu2+/JYzrBqFQbcorM+o15mG+GDqkcO7ZvoCBN9dfwm8wGvY+PGPMEm+
kdQzYOJIcF+TmCUJKDn5MRnqnGuiCuMv7CTkmTjLdsekCe6Xvg0TOXLomPOMw0Fsi6nAZg8ASv67
SqakVithGy5vPaLuH+4r7zqr34cINbNfJL80Utv+4lTmoMa12paD7+1jcxAP0Jjiuh80vd/+4XjG
6xPJFbAtpigBYd/1FJuQeWIBsaGAFzyy7Ehe8+JdmgB4ar2CwM0Z//2Fuam/cng884gBT5w1rsBr
mqSG+TS7lIBpUlEo9Lsq011Gq5/XLgz54T9iWL52+ww3NnZ5KfTDtqqRKo19m4LAt3Z9UsJ4yHP6
9D5SUNlkkwFfV5teeNcNTtxq3eRpK6FjEeF9cDfL08WHPAVaeS+kqiQA1FdWlPIOWTbolbHqIDKr
l7aUfj6Wcu/L6Lbqq1X0g2Ivz/n7O52OhfdOQHK2cGD9ME4VbJyA31eqKbWUawro29TM56YA+AWu
B51R5EbcAD63OtA+DI6ugTDA0rUlWgTgrI40GdoshoGu8YtfyldPxsjcqvFMw7328g4/J2tiU4dX
JqhCAaVy7kWET1Ih6t/PW+kiO2pQRwtuHhqTuiQZjCL1Ro/+//CTyYKy7yWS3wj8o4PZzghirIZc
RqarqQ5zSXTxdEQHxH5Nmjd6JS7O1elkjuVc/bYpzhscmO+ims/nqhIUmtci5K4MSmrAQ30mXs2v
iH1opArjB5yiI6TgBZfXipiVDhCWgmEhz9+8ExX96dTpairsKzGUJn/KLaPeNXcDc4c3YhCJbV3a
jyKoDuKPrg/nrNKp+5YueULBeFuyqUirrjsAxdEQ+29zsnoWBTkB2q5/f6Qg0s0y5U05CjPubX+T
g35pzi/ptteLLDxcVOq62W3T7pF0fEXQeO0Mv7/qLm1NINTrKmzdrZoJtTPuvPwP8UJj/FlKf01v
OG9Vufh9FKYqdgLFVP+oZnxNPE5De2n9GzZP3+nH6E/SUAqk0inq1KrAd4k1gdPHTIOq1+IXh0Pn
lcb6hfZaoPcFhT07fUDi7Wy6cxgx3E5c7BQEZ1QRrEKtSzheEZ1b9F/ud3iQ2RYfm5cm3dXEKEUf
EhcuVZzqEezWRHN0HOvBHmBsHgUls1vROWEJJyHJ6Lu8y11Ef2MmJ3daNsN+vhctNvXVDMMZ/wqS
Mu4Vm1aaYi0SCY96R/tlf2pEJrPnTKUApUiS/Fkw8xKE6viTNvvUqCIUwp6acOLBzQctyOe50QTo
ghVV+e3HqGcdIhllj//0KRPcoeRzqYfRlEe8V0MkcGVDKaQWpn7spuU1j71fWaqGa6hj4UpWr/8+
D6WQE/p6V1TDnBYHiaXZnz3ZEZmbmrHqh2ibfJXS1651eczRTdfrEawqEpPQ0dQqmGrSo0BSLiO0
TfC/JxQqvGm7j58m7NjkDwbvqSwliJVOGQslBRCWWh/rdsSmte+w2HDLRgjycYjcYoC4mze3sguf
VpXDX7KQMzMi5srVRpQpX5KZTKYbMA/YSfw6Bw54q4XfIVwRAFlNxKmWUEYJCDxpSFTeaiMVFGRn
RWtng2gDE2bVqMeXO59/slBg3nnTTmqpB0xJjrinrOQeE5s3AkzkoqoTjtTgFPojqnZeL0p4jc/S
JWe0+yhIKPQydBs7rwKFLHVCXrW0pjWHWng73Lnn8NSLQSPnI51+pouGb3QRXcPmAQlk2VifPC6D
eQrzF4IMYNaCL+oDfDcWqm0eA1nksFHQdavqw3343ib96DS2ogumphe1mrraxC/ebcvJBOGNfU6o
QiVx+pqdm25FDd4+LuZ+6Y5pYkE9XFkr5q1sZcGV5jpwS4cVVt3okQLWjYp/MuMaPESrYe3CRAVh
20Q9vncucN0L1/kVqsZ0zykc6ttDLfWqTlUE81rbABepNniCuH1cvVfY1bJb8/hhQaeh9xjKLnLZ
vt9UuLKE8Yh95Y9mq3ZiXBRRgqB7JKgMXnOkITdGsZTiWox6TC8M44lXyO4XQNaWg8J/1UvAxcgq
FQ6pQCQgNuzxXnMtyZAW+ABh8XPI07aXBKb2APb/2hvmlJF+XYIYrtp0NX+sjl7OzNH+9jepDyRl
n6w3t+bw5QKOIAsIcPEa99ipK7GTHODzykj+NPW6SCssGbhK5HhbtHFSFWwSlTAlvWzkvMdawqDg
CWbTCvqJBlI88JeTYOrPb5YCTLU+YmeDcb2ihKC1V0QguDfopiIJPBKhN/mXm5o+BpHgsKwBNwSy
DOWvRAHCihIWjnWKoRhExCWlRlQ3lL6UMGCtXGoXCnGn6AUoTx8JBA0dx+c9pl3T7mx2IvmZB8vD
lmUyqm39T4AIsWZTNmiLg3IROLncVy4TKmoDyQ97hSb+7kR7OwoEAzH9sfIkL9MLpskEczirKpo/
aggUWDA54Vnudl+IEcdY6lRipIVYk31oIu5Gj/JYSqfDWZDeUViSzKVi6pFna96YSL+z/bstuVSs
sqrO58DMu5Ttu+ZA0W+1NkEa3sF7mBlxj3OI1cB4BY0/8oD3Go69B/jnxZd9BopHh1qw9vSqYEy5
6gjeO44ltCdbaa74rFNA/J6v/Y6ulf/ftoPODUxP6RlwxpyZjTkypXtlZZsTJlypW2EGZjE4b27F
xF8HvLPxhePsQuJRZ0NoXHqJbQ801NxUFUhWAghQpPrxMEiA1sqEp3dlxiH+ocUARUBePcepFDRm
Qrnfqf/lX3lCAJCkfmMG8cRb+2HptYOG05oWW3n+HIPBLn5zAYynw83Sq8AQWlGlB9JzvMdPBSB7
fUS9fE8hifUM3GIbC/7FY1RxBPgGbB63DCHmt6KNukhS5SNjgw9YJRYn/qFRLqP9v2OIa/gfJhYM
BlpUNQmykgqPadg6NfaURxEuu0xWX6D2h8nXOi7Vc5/zuilJK9Z7l54iN2uwBJVDs4ihtWy9FFsH
2/x4TAKXQMB8xtCe2BeWImzmEhdkJS36waxtW37oiT7MxxWs3lRHQgDTiWClHsa4pDy5GSJQDyQH
nrzNOfmIiIqZH1J+bzUbbxYG14pS/e9KBadnXAUTQ0xHMJO+oR6JovV7kSUXEoPM2HL3Vprz/lEu
eX42txDMh5iy4lhARECUPKGpFZlCQimJdMWfdxJ9mXzFCAKYkTWXHyeJjjmFEAYbj6/Qz5oVvg13
2W7bmpw1adPU/tR+KoZMWO6K+AnyJMP7o6Nb/8bCGgzH5akpZKoBrqc3xCuN6z+lE07DjWuuK6Cy
6HNHBwmczWWkUzZBdZsxVAV33jZuScznz4kqlGNtrZNQ+BKBRKfWgTLzsHVDnvOllhXQ4V+PS506
N1ApuaQx+DuqG66krkCk8re65UoDN255odJCwl9RvhtPvYrIX9XL+poXMvcMEHKjAU5svFyKm0ed
aLLkKMyzelRJkjbOlVgn/+/fizK0ubRq6J3RqKXWZ5UY1SWwaXd91xUwizLbtKyflb7LPs9hKnd5
8adYL3qgEasyZJmtk6GPpVz0w/J7hcIdjbmgaup5+WU8rIpKUX3KFXDu5z/t5D3N6N3dhWccokGR
JtAKDWB4nOUhxUDcSLanY9b/uD0Ji6GAt+ytRtGQAzrGr9pIK3Rn5Xi4KQyKLYLsocRDy16XzQIS
e8gPDKAC1eXv5EZNvCtCaEbJfVdGiOdpeEy9eyozilk8LdRSamNG8OWNBYBx+ekOX5FQneiYE0bp
Nb6Nd8PqO2oPyfYdAgz+gWf+cJ7E13382YYkTaa6DT9oeQ/1LGDLw2Kw1HibPsPBtayytnDUwfdw
hG5p7w/k/NLMkggiPh+USTy15tnYVuQz6d972gQXqA5Hes7D/qmvC+ewUrvs5wf6SPj6WUpkkfqp
D/kFcWUr07g8iG88wg/o8y94xd0KHS+7OkMVkDIRw+8lvxhY4lykS1xH9flLu4A/YohQygSM6pL5
qaurvoh9R7FsW7xHmw5LncOsJWxy/Lfkb3SsXnQfz01zgzVirIqX4UBdcYCoorSTygCXdQ9iVhMt
lzGxbZcmNNHmzYo6A5UWt9Kt3y96hg9pZWK+nxaKwHUPGVSKH5AnAQ9kyTJb1ADmNsMltxpY2q1t
gqbG0oExetXmCUS+nBjj3WGjhj6kjFN0d3imUVUDHm1HStu1vrJMEQbzTJhf6nW0ZL++/aSYiCsF
Ajlvuh7oAHm7cQrT/54PjXSDosT+GqeUoObDntV5J8DoK21BJjU42Pehwu9JiOsU4rC80ID3nQpD
4yQgEnJwl/MYQjN4pwL9t8jRsNJaX5c0iPCmvcoiMF5zUhOSz3oVLuCmbmd+6vMbsp8FDJdIvXys
pqY0tytVib9u+TEQFRxfrInnvRncPLI9/P5NBUg/tQn1wowRLuoQuhw1fSu2c/8PEUxghoXoFDyP
EDKQmLmDWO0wkpiNFe33eLgZ/aiBnYcAfmOh1nnVxSCRXJH25hcZGq/6iPkLxdWUe8Vu2r3pmM74
uEEQ1AUyebiQ4BQgONEEiEz3cvgy6nApmwMvVi8a0/ANflj4JXhjDSR6T11DL0CBRqUDRyIDSrjh
yFMzWk5VlyQeKpsboY2JTwxls3BdDNLJszj+igIz/HLtWFHMNTRdGwzzTZvB2YF9H69iwN/jUdRL
jJsWbfc15mkd7A01KJaVzytwvE7mMzn4eYmkakVsD3/ePwLIzupuwuXKwdSjvvFOqAB6npuJ+AkK
KyzdekleW4IZSCCUCsF23p9KXoW1lkBi+7WX9aJ2ZKX4LvypEDGeQUbmQrPkej/ca5JcgYikcCJU
PFZ4Ic6nTSGDpqlPMwRUMFZrDdp3MCADTO3MC0oluc7Neqs212GOGAZipAbxxBRDEDxBlLgRObCH
eViHlJKRTJm1SqeHF/ilUK/qOahnkmQF3ZcvGeEN6Tv1Ee+cYF/KL4dZBVZaqh7yP6jl1/dDdf0V
MJQSuPJ9vsOx23KSIKfKyU3i0Yy6kPLSdvMynSICdJQpYkhWwUN2PuyBDdJYlxSzdyL8OvYuNtQj
27BaEJPnZICYcB/U+lxeC8RauGUCDZndF8KDhBJaAlM9mbk4sV2a0De+ooXi+iVKR640qeS3AtGs
BT9zspYaOY1AMb1zFzNYimoAbeQ8N6p72JdWUjN8QvB2lGaiS1y3cnhotEVtWbeF4XT/jJEhbY/E
y4163vcG/4RtBpdyIOG+0EhEJcYJB8gRcNl2XpuuySA5WzaGvUxn+HtQhHefHDkiUJtkQ5Gs5ViZ
d1vhqu4ssScRy/EZv7FpkbsOm2YlStmTHbhnFrgpVdfmml4wDlvcb0Muk6SPUfL0mGCPJUR8Yzzi
o7hEKDe9dzQ+swsv3z5Q3DXIDGdUQDWjyFLYbtdDYZCglvuJACG/kZ6l7sEUMOohZzPgAzi/li1A
tzJ4Y+LPwetw8AYFlMjtTpLCoaYJmho1eopa4FUud0t8Ok9AyosMmSSLzwlyK7CM/VmWeqLDkSrJ
vSnteFJj54BamkkYIexyZoYX18SrdsFdKsTsiUuAuGj5XHxn0Y1rrzrDVyekZAC/TD3gVUCoXdnI
JCN1RcRXNztgckw09ljwbopiivDnWp4hEZp7ZsGNW0marOOI0XuSr+5HYIAQmLybDMOikbGCfQ32
tqw+nDBcMA0nmrcvPpTGZmF5Tf1nfKpUhvHhKHzPSJpVQRPkz2DV3Keczdf40XtSfk00dKqDKXc8
zuT5lzhAYf7VbeJmXNcqJphZDakhKGGJugOTSOgFllccInIqRZRdv5QcXAqYKt2qw5g3A9pfLkIZ
V0Iq7zn1dJ+T4UbLsZgUavfCCjZg96BZtxEUQVnIs2+xGh2GQO84PZWNmi3P9TDfLbOQkqGesV/s
ddzcxIEOPkYnbE/jmeMK6Lfl8t+HUPcKN7fJzodflqVfoCUxCNO8NvHlpJaq6DIrbaNbj47Uupe2
1A9tBBTyK+zd5Mu9HqZ4AIRrdUs6mTHFrEsc7q88cJeDBQFIgjFRSvuOSXezyIovYbfCIzSaAHSL
x+VukyxrT1Mi39KPn9C/1I/mXQqt7ahdeoHCmewIwzlcfvcj+xuIHKSAOojl6ob1ZqpPhBfSJPFq
n2NK2fx3N2NjfvoxIZVmfz7lcsycpzUkQ2MssJBwQDgsFhvpSZU04M6J2rQuiWjNRxWG43FXTDbZ
B558og3bx2jZpmws7AGZXGp1nsxEuKG5ctSyHQB/fzRyxjzHwHMuX5+sbEApSo6/zn32T8yeHImU
bQdQEAKaBsNxw4X2uVPxs7ydu3RyX/FtzA5VkqxjQVWM1IKnA1Mw+HoZesSXd9lw1s/XqvyAIv1F
RT6k4Yw0PjMZxcpdwv1pZ62P9OQ1OnFUpdQ8NhiEk5JqzQcVMe+sQsm/r9IEBDbK1rdR6zz8MjpD
wlsMTUiJ6Llr5Hbd8imSlLof8paccUjzkslrroLU98tEv+e5kzkMBetOLeUUuQgBhZvgvvcXnXIb
OPmj8Pe0ao3OYcTZVKKh5bCeC6A6cZrjcgHflubzbkW/dkwEo2+6JVZE2H2ARbhy/OscDX9aVHgG
AZQM3Edmp/fCF6j293HWQ8SignCL39Z0xXAAeoyIMBRD3F6kATqgBltZFZWmplsGXcJjFE3+oh27
ape5VzdS6d570pp0pYAQVX9UDiHNPDr52fu7EsKQvLazJ7JEV+LH6wiPIgRDGlU5odUGr4EYSV/U
0nlnE1tCLvdhSpxVMWXj1XXU4Z7kLVCLP+jVAXnHO/C/FJgEJDqawCa3UJ+/3CkAUBDwnbPa1ZzN
pFJzPom8CWzwUGpr46DTF6Ryl+1wqgA+/NYJbQ/xk7hUqt6QmhFZlenapDx/lVntTbEFEe28eWMn
hodFk5kVCE8/3hkZVQUuKZfdxmXhkWFgIUt+tbJLf2m6uLmAaXl+SrzK0lAnz3fNs1WDvgbXOf+1
QPy2WgZMEnXD0T78vMUMTsLsbz+w+s6r860GYRFfOPl4pTwYSv0Wd0rGNizlBsdskI9DyGJiPuRx
yiN1fjAivC0Gzc2cWTGwulbEVXe8IZXJ2LNRqbOI1Fi76ysRKT7r729922bf3deE7HbeZgAtgLZV
qeo63AdkHQtXyhrKMM3NDSNTr2gsE47hVnLzBWsfrC25oR6NQMfQf9tcbYSm0O7/Mxd5M60FEetW
9kyve5rAWjl48TRMGuAiCAnfnDZzUrC2sDZHQSSL2StKuZtW3AZMNScGp7b0D0Uq+jx8p95aiUiY
/tZfDZUEiAkxfEng3IBgs8vgGUIkTf8IfjyZ6l7J4VvKQaCdQaFSwgAiiWuPuMnhDHqQih/nX5eS
K9ffTzio3D/Kv5fOy+QQod04ARO6KLIPYC88smYM0SY/nOUh2UGAfwsMvpuJ5hSOd+iAtMBKmmfv
NlJYkg77LX75kEDkHmHkQ/CII7DpFFm2zct/TAJmq9bWjP8q64XMP3iMo/Z3WAjAEzf5wZuIbCvO
25jTuS3LydlWMhzybpxqDxlW//zMuzmV+QNMEDRRuzhBeO45/GsCek1+Hp+0bMBxN2zEOv/Y4lZ1
G4eoPPY1Z6SuXGl8vuTgoIW+B6lfMx9n+jeWAKAMqFhhZ9dVSh36Bo0a1+xFRaPbP4ZE43FG9y9g
h0oWAaeq7yulyfWbSpyjhf8s5z7nmv5H5fCpAgORUpSrR2dvXQh9A6S7dNZbAKz5xUSE9nMF8eW1
hK0zb4u3UHrI95aZZoxiFHJ4mCt8BAkM6e6LJ6XBOE0ZOwCmxKLKJGeX3HN/SSxH/vG1vTTbROlq
7VPgFtGV3tnqXCrLWhcbJ0ZFLe57TRprHrThz+Rf6t9VugyBPeoWn4U8YIPtfxKYIPhBGphisRDE
oMXYc1wtqMet9hxVsG938Rys95aAKLYlV7WVI0RgFN6iRwyzdSwTOHZwvQLw54B8Kvc5AXyU63ac
Ihik7BIwzFrAYXTEZWr5wt+mSlN39Fik0c494GcclInfcO8Upgo4s+ZqBszZh4dScRXYdk4yS53O
DQyPreG+DPSb/a66kwmuf9+zYNq/jStj22wpz0oZOHPztIXtTXkC3xsJI1q67KBTuTO3zR4m8CGF
Nu2PPKgP5XfcBaiMWfwypxhNWU3CNYveweVc/3xlLepKbYehiyi5olwzXETT5D4Nbd+9aYmHuf9x
+pVevYZqTPNEU1HUaUTGaKFWZYSevMU1MmCBOzcCRfxSa270wsTcMHTvwMKI+GxuJoyOsex+F+A3
pU+BnlP+GsnnZqTaq+OeV8aNv7aIvimx5ocIWq+IFwG5hHDFhQPUnZNRPmuThGJl2qU8hHab6FRh
Jsmg14sxmwgB8333y2kTd6P1Ov/xGHiT/8WVP07hVbFpRaRIfT7XnM19BoNOJ1fHF8oCnNrc3tMb
MIiUZTLtxs09vMRtlDjMlSoYdQ/6gHh40jjkwpzb/AwCQc5WRQuQ4CmhaVe6SVu6Im8h7RimEKZl
SIy2AocAjr2BD1XflGC+CK/LUWo2CMnL/10TKwqlxw78t7jHkbWpGwfIFZum5C/jIT9Bjj/XnRFJ
aRuXoSQaT4z3iGy1IzvJ9zDX6/205OD0aHw2EpLEbmKdfWjuz4YameOtXEmKPcib0EjsW1/38TyC
/haPeWsOQsW3QGijoTf/Vgo22PnuDZVmE0R/LhNWgnebuIc8HYVJXpCBdcqbkwfQdJwtNIGWe+R9
vo8pOu2NNhWvRTQK4sDGf6KIfen7bVVTH1fqKClmQ6J1OZKSJC2SMEQ+d0TNTgSdJgrAduFFYChp
ttQx5ZLYGaAALrooX2F2NFStA5P0mwyjRc92EiqeBsyVuBHmBytRljKBfgjscfMj8GdLFEVmou5n
yi2lp3NlMExBzPA7DnCBUJthjjqznllTKag6fpEKj7zbmEDFDwxELHNYLodbXPJMfjlVrsGLtNkH
/22JKIF8s9hKkWFGfg+J1aKnQHUSlUabPzlej6QQuXQ1gSnPaW/KnIkzr4O6XLTfzr/EkQm2NBq5
6hAATNUiSJsJRMLjOXr+3sgaV6c+ulmPcFT8BouQ4aJSwIGANZJ1mS7So0Th/pkwNyPjC0hPijFc
7HED5vPB5Tiz0MisDyZX0Ap0h+xKGe/JR2sxfS8mL8qZ5FxXp4Bg99kZdOq6nqezJxJ7FqKeuk3f
0q9MQ2nLXsiN5qLU/TMBzjp1vZKi2ectg+m9DiZxM2PKbdcILQJcwdGnp1U4W7OA0AE3/tOoSBcz
2nqxvGYDoO68e20EOQxLRyv4LXbhLE+UNgEvd4vgEqRKStq6HUZhARp9ONZUSb+1XNfDu90yqFQF
eCKNVnyThsGKKee4XfNz3Z0VXX9z82FzaRdGc9Ph8+I1gRuFtZi6suZbssBE7Wpj2ctP7ftol6HH
/nmCSjwF2fx5f1UdHd7L6lQxn/Wod1leNunLUyAl38SMbJSNCj2manIYO8xBIloKSfE9TqJrxCzJ
h68P01Q5BmK0CuW5Gdo86m1tGxWGxFDePMmlQAEw11krCy4UscRhIZYgkSAXXmIIQeJY15vEDwol
ktJRH6nZF9u9VpjRD8Yq699luvwr9/Q8bdHeoW+S0mqrbS74c4JgeN+5hC5YhFDNZAnFU1iwMeNU
3DHJ5+Uacebn43nA/3u58VYRxAsTLGfNqLoGki2iJLS2JSKkCbseujjo4yrVCXJ3YWKYi3pjt6GI
vkQHsH0hx4n3jVuA0jsA+REXbS9uB/T8MZDpe9wpqKQVA4rp26cekcmsmHxGRzEGeotSGX+H/1bm
ZAn+adwiWfcDNyaGMXJapGiJX3TSw3JlDG+RVxBwDOB8k4wMK4auhV59mHg115aqC8xulM4Y0vtd
LmFjzmH1LQ2KJaUnwwmNnUjzuEvqAjYuvwlltywvt6ykEQmrpTF0l6pP2WPzW4leUFFR+MFga/as
kCHMDeZgAkwC/wxSF1dZrqC3ukpp2JSaag1RaIG5V7NjZx5V5E4fmf37sHhzXgtSmS7h/v/gXbNu
ueza9PenZTXrOP6ldGnngLHGx2LErsNBKUNlCeWSHUG21AKEfxhtGDQA7Poq25JS1m41JP9taW8P
MPCg6VAYRv+WHI/4FRZAoFXoHq9oxau8MCoWBvVyE2icRyHEZ3MDgsW21k/L6gdZBaCrlEghGD/r
sHmpwOku0UNtGx2htc6pxas/ZcChOku0MRyDP1esLturo3KQdGkNqgEdaPBzNswCELNwPUmRvrBB
hX4azVl+uiaaHRe2oEY7gncD+sjbCO8gCDGxra4JIZkrV6d5mUT7JTFb+NPYbLh+cn4jHq87Cbv1
JnYxOQvPysVrAOIIGU45RmSG+lRaFxB/Bi0nGse0S3uec1IiwbBH603dTwBMvu1cV1w1n/rrG2ub
USb2l7JRNbXIRohr7NOhIHZ5uqWcA+KD7OldT1y5hAZwYV97XO7VJDuoq77qni/HJSymtDlmkMRQ
JDfn8BaZM3Z8kSzXOoZo5Rv1RV0n2DEX/lKtSKp4+ctzM8dVIVwtQ5a0brIVoIqgVL9/F2LoHdMM
Ixpj/jUcW1nGTqsYQdUwHGDhSFahRySh0x5GUBXyC5wiuXwgCNQMJTrTFZ22T1WOQiJfcDBiRvxx
yG0Gc58oeYdhhnSNfXzg0C3y/8s6+7GBpNcKMbOYVRsc2OALScQDG8CXVzZxZSNF8bfKo9Jx4am0
C/40OCXcew21TT1+Cj5WQxP/zkGbcqfBo6AfrOim1Kq3V8CjRjSXJEbfrWpPhsB6uuTYs+qw5qKo
nnfahZ0gsQsJsQ0bXkiw8qpMptaHrGBirpSKdP2aTzTunztlDvngsC+bIx+uCTxSLfFZxzgRBv5d
P/mYYnNG84qPBuZqU0xuELIApVsdUjXg+pnqA0ArlnNgHZ9gE7QzB6TBqpMaTlaIdiSAotsAprgU
/2cjuMnKpZ4nHD6XW6x1UjPUFP1A656IHSTXwu0phU4L29/uPqBuAWUJ22lCfDO5G+WW1VXgwgKY
Z+ZnjVKLUUAekE6rzSMXfVppuv5hj55cHA0jKgm0ywx+gdMD8n9/CZZkNuTRvUGOiqA0kqJ6/C2a
uRgeL3Xu7q0JVZkQWCkPEjTHjX6Y8DhJbKhXRpQWEIlJVRWF2y+/FS409woLokCl6mW39XIEHPJs
mf6cikUpFBtPeEd9eUB5buL3TiVI8pzLy/ke8VGTYvmZaoshQmYADhESwNxSsHpzihohGQyk/th7
6nEoLLFdRv1AsoXGsic0L1M5f6zYRM9UGvrCyab6deIf8d02aDSS+lNJ9nUm7Y0KDm7qqZszYKXq
DaeSf32P0uta/GauagszrmZtyvO0IeDxP8FGo5Qg/+6J9ziQzIF6px8OEdz2FdkCO4c7nMbM/G5k
wh3uq7199Puje8/BgGsdxrzQRoIMAA56MyWHPri0BF2n9b6m5VKgP5mdsicrrql6j9JZwu43+Yrb
m/4H7cae+P6E8wIDJKIbx2fzlVDcCznszMqYT4w+4NAOGMWwkjfrvqoeDZAsxy0stPoQ1YNo78hD
xU5728tRfLO0gHZxOqUqTPuAsU7BLnK1jD35zi4wO0CRxiOI9B66CVTn5aNyJm+zDJ9roWluHgR5
nuUaBuSPsCzsBKDRLGmbpDBIZN3jiIIehFIudZblqN4tuIRRR8CLlYrT0TXCGzZKmX5Zv5A7w3Yu
rnAm+0nwU6+8zB/rG5f7O1Bbcepv7NNo44W0G2BlQTjGs/SveK1cmG8zFEENPtIUPKwzRBoc8EP4
UcU93OSQaCEM/V/sF9TQLZkjpK2ejjTvFzTeruC9vUwf3hizdXN2p5iV887zl0UX8x6BZSLZ0Qv1
EY6DOg2ZdqdZe7YeLtnoeuqygc/2a5C+VFIlwI3U3+HSl8HGVFj1YMCftRZhbMx7QJ30Vd3WZYqx
njwDlAkShhmVzo/wsXadq+0Hay7aY0mXa9EGGbH/Zr2o2qJpToXHaN4H1+nP4h3uRgVPXW1XKL5w
w+tOC55JuT0vQQ0o3S6MQe9mWtKzFEd7s29U3/P4FlT1f3HSohdbiLKqqQwVvfiVeNqCJUoMITY1
lzLO9RhJGjYQqN1FsTDcoWExh4fWpy0/hhMC5+sLYnydTm+SxbS8HlY0H+F/IAg1yewLSF4v+bR2
0AZF6qtJbQZn6v+/R58Bt5pBPtrZsR+1PXZ8VkhPODfAck5s1eH1frEHkF7Cgxpr7FhsEoT8oe5V
HPlkJmwlnFYMJEUOnWI6rXgZVbDi6/5lrSC1wz3wlGJuHIkqaUJkMlg0X+uSbq/U16Hf8XvmwXtA
fXkUWpUNkjwuPvDP4bakkoDBoFL0gvHZrhRYnu0FIbAHCGuWNYPl9+zLMmXeiQuknyqSww8b+uYS
4B0QDtqhoXGrlhRtQ8oT2a3gPFms0abRjLOFl9O9HYnZnByHG+nRypSx7TNn8mqbjsiHxHbuT17E
eq9HSflwTsqKXTtFIIimFpcDCfC+kWF8WyMQ2/R8ahKRb6Hvz3d4Pqy5HDOcveKwpKQvVdjuFGge
uE0F8Vl7Z1qOprJ0JeEjYRP7y6G+93ZacUJxf1VlaVlHcUlx03jjLl4M2PFiDwBZFaxFZIpxU/zz
jlFNOulQZ5Mq6I4qhC2ty6fjaeTEGR9OQaL5dG4zhDkNC+wyndhYvkNHSxfy3Qo9sFsM+QOIMJcs
FhilzSx785OejjlfW6OLHxrFXU2jyGoLOFBLKWtrKhOAD1iHj2IPCIAmIGjxJ7dtFrgKDJf466pI
Gj5YWvwhQGUc9pnvVN4rC77kXMiIAkKi4D1x4IZpLBsG4BevptVnoQQict6i5fHYqYswpb8L5PHi
4pFYF3t4brOF+0+aznQ/grBE1iM1lD9Z4fMxr2Ljwa/lR5pN5IsRWIDkkSH/T8kIqJ8aXHONdwIH
gN0U94drSRx/E1DYY4DP/z+SxSO66+iK8jozzW4OuLG8KGJyZC0OxJJizSlLxSLrz6GaquD7c+6I
sNu4FRHRj3TRVZWEAvCOTYF2yNm9GqGQLOPAXPwv9veYt3ZfjtM81Sss6vbc58TyLld0bnyevYN0
kVMMvWwvwQ2kZw3T2do8Ey1PIbe2XA1M5bac0En7xRgmrV609WDG1c9zZntK7rdNJIvxBkfV5IEO
y8CYkY/KV1mrDuy7npfku3FwKF8Xn6Rn6Bu5657gk7XrTdwB1FTq2mhsZz/FR1lSlsCfnnOlCI+m
aO9Isd8m3b8UGDv96EtwtX4LoruSPSUz0OUzqyeKDzclR8mNUp8PN4ml58ticeEL03ORT/JF6n7L
KHT7t8prqlSms+0f5dC6IQzuSvIztezYulue4NB69QwR+s0I+e6L8yScsRWqBx8k+jxSlCuvVj5y
m7bfUGkTQPU2X50dG3BwhX9ygMZl86QV2bL4jIzHalS5Qfb4tFZWhbw4IvicwkcYKlmeS78t8KE6
cIg8cYHeRP4uUO39DYTTeILuY9Hincem9YUcFU34nRelYtnSWVfCAYDwWyZT/7v/VcLCkyQLFA2R
iAX+wsH2ODc70IWUHYTqdoq0w0B4uKpkay7S3f2p8IO+RyQeblmIH+9dZWYeMewJ2h7jf8HblS1C
Cl5I2BFKkQ5MbZwRrf1DtIUe2EXyQmlavDW9AQ/dre7NUAfXvVwpkf8Rt/B38JA/TWwmCMWBtQ7l
V2q8jP++pzvjViEk+Iz/LtW/bnJwQD4X8fnQbHe0DhnEDuHgiPpWi2cTEJCcpQk3AtGm59Mc8x08
llfFMT2oyyaV3u1pO60E2FlCqOj5MF/R0TxbdtgF1qltGaEqoSzW8WUAsl/NnVUeOxcagLvOTHHQ
2/JPLVi+JXdgA4awWDjonW7cMZcxeWsA95nNEG6ixe6agDGHv6Tfiy2O006frj7B2jzryhj8iVfL
FYoksc1EJ3lAnXCs3EaKul/O2uHBPEdScoK5Qcz7fa3/VuvcXD9UX568BqLXJfQyqFA+awWZwD09
cxwTBdJ0s4Izui1oJydVRFdD8qiEapqrC30NPBPMqbzqKFJDtX+Fe3fFzPDjteqOk9Y5JWJVWaCb
NfbW+tqgUH9C2GjVyFjc6vd0JvSxH4b47hPmxfiDV0Djx58sQoEcmceaLzIe5PtUqvFfe2reeISc
4n1x+gd/P4CEEizuGtS2Nhywf/52Dm9tyckRNegIv/ZWcKrFglkq8ufL32+L8fuMmMLi8pXWGm+G
3oshGS0PlmpGtQ3jhQT5JHVlZnz6Ri6lepokNBPYPmMe0DRW+/+xva+ewByEHZZ6CHjFq2cNYZiY
jyBDpFv8nU5RqKHOPET+wD0fUhmh59ZIU4bFnz6ilGTO7YWEt30BnV/MGrRELz4R3nxpe+/0iWTz
rf64RejKFFmenIuq2grq8NtXpSeyW9FxKCe7ssJPCqJrvqb96/TaNvqHQS57WKWAIzMKiCuZFE+z
AiGe4xhYMsmQ54NvGtKf6f1KD8MjoAsrMZR6chFce5mbEfL8lUWHRDKo2vMgpbgZFkHHAefPURGT
Jx1tFZFIpl5pV+rQNM+/oPd/qDMr8F2qT0Hhp2TxlQ7ewmkP0dkWOp/Y0EKAIaPNyTqby/haTNSR
JoHOZu5RPtccm6JcFWBtbRaWEoQtP/ll79SGK821poY5hmr5+lM1U6UCGfkEaWGXzG7Xo+aUC3kR
RYvwHaYdR6uw4fZgTFp8usOy3ujddCXaLlV59V4aV/7QCgjUakqhj5bvrx4hJlT8shkmGK6VVwEn
3sw7QqzANg6ouncDTEvC8VDlhPC6hbvaeTUGflCyk9vShMcoN8RDJcEnRr8WNxU3+oXdnbJbqkLN
Ec/6smuHgyml23NMpitnxVJzGFte0e7WWgfLxYuOHAU5K7Atp7wWZnTNJiibcKSnwlxtNeHZgxY6
D+BWkHMO4K7U0bl5gDaKtpQCgcxBhUJYZ6Jv6De5So8AZknjuKtUF9ySJqV8yWtA8B0OdjDQGynn
bezEXFtrgK5kLNBKo76lXhxtWXp9mI/bq4IgsKiBR2nsUwf5UnE/BEwbI+Mb+jkWFEcXiNF8Aula
aiyvd0CH6sK3ByruEOIpjopKGCpQkm3kTsaQlNwhTu6vSuIToQvXCnVuZG9Y5OgWrUlJBIjrf31v
VRYfnFr2yiF5NVAlpdPbkl9WxYfosC8IiV0WnNbyb2qWVlY5sgyUgpiqGcfGw/F0rdz2vQ84BGs1
EHW2dQ8D8cKkujCaEQ+JV3qOtfr9xXVzoNdFvUQF5U1g90Fxv3AdTVFvwAfGLPu+uS+UWzXcIis/
lBkqki7DIkKg0FrBnsQi2cLXvO8qG3J3dtMdY4LAQ9hLGX0E24+1vBqzehVh2gMePmSHHkTlod3F
Ps5rnD3dp/6RRunVdzhDUSv8gcp5et59OSct6tAnPrrZ/3jjxfaemC8cQb/p/gU8ysufSO0IdAS8
zi+EpLqQ5Pa3xIq7zogJaPeDZsMmmeyqDULH7nXONPz9z63Iv36LNGd0LmzBZLp2cFimqVjXv3m2
Tp0UnrRszXktcTIp4cjQhrN2X6AQ366ih5/3sptDoa8f0pBHt7s1+VuXaOWjg4vx4iLKsXlzdOIX
R1IAYDIesUx/Gwa4BspEq93yFPmS42uU6QMCUvZCnUHlBRu5/uRmQ/DqcTBHfhEAZc86pVw1/5qy
MD3z5Ce1abWoIin4+qOXs2Y+Gbw2L3gfiSY2gszN3c9WPivNANEMqcReLw7j3l+L0m/1+uCcMJ7y
nvkF8C+dQA7tbUQTKKbsRYF81TT2L3zs6sh+XVPA8biXS7190RrvspKBOez/J9DCp1/WGyDM56OH
hUyu1aq4rv13ihXOeRcVcQ+amIJQS6AKa+hcpCgtMdtcqppyzj5wrLBxE9WZDTj14LdXPepGJzBd
bjtZqP+kjiJDR6964IyyKI3eZcl/VcI7FvDxKIR/DpahYTS9baH6JLbNr8FfPlDkqQYeLtiTu9hl
FsdF+cGpakFF3PhJGCA33YhrsRnfKtOTgqz8vc+yxGaIg8KLkmL7eoBKxnkWBVdKpynaWnQbu7jo
xIdM5FhuvwS2B9DptFYSloGmyPQtra42zrJv9F0EJVVG/lhY9APRM15QU0n3UXIAFaPhJLkgG/Qh
BbqEF1qiWwb/ZL7L2vxDaPaHfrJoq1kF5DfSuUbyXiuVBESgCaZItLb7+pzLDgAGZc4nftfXm59s
0p9VfiKZ9JzLnvTkxKLx3la/7PA1GdhSOTggL833fn9bO0JMmDI6qksL0tCc8NJHz/niUtOZTeen
extG6sQyVCiR0fxnxL/iVvk2wASrLlxkkvynxY2oxrUnEKcZxA6LZcvN7doV1RCuyA64r+oCscgH
c7er2BcJFDGo0YuZ9yk8LgoX0OXIwWtaKvlGg4V73JcrYRxWCH+LtoaiELrowPYYTQJo5UPNkYEW
vJNy91AeDa6KU2QE7jgdknd76Pq4UflmzfQXBPEeg/2fE0vKkPs9YsUkj7sef5XZAG6UVGRvvQ1z
gBCkTu1khwFNADS6ZbeOQm2RGodGs+tDcYYFY88HCtmUDnS/vmQPfHA616DOATT8XLkRFctcLFVQ
95YMXqqgcGIKpKtHQ8cIDto2hURqmH1oBI94XRfTPZSmCGbRC5PZPGu3o+DAMK2+8HonQsOJlxW1
MF6HrlPYWCbBLP0zdnBVZ1uqQQcam1XLsdMs/OJ101w08Hno5Lrbq1pq6jGrM9m4nf/0fJzkoRhW
HUjs14p7egC+6BH9GpG6mJL6j5m3f21YuT/r2R/vxkN6yDQakXrfi2xHqh+0CeOIMW9sQoktG7pk
tkBAzD+CaQQpkPdORpbamq0zrbdR5ECa/cvODMtAeoMitCAN+2qeBDFqEIgQRk4pkltZ8koBZWLB
GhTWJEJ2iO+5dK0BkRyaBt6mzIQ9kK9A6gMebFa+Syfksu32lSo1xpph7/IdUSjC7qyY2KO8V0jJ
lyWjJfkywFMI9nt485gFcYEsJWmBOWi80cUD0ezQgYQik8gR4rRjdlSfDzJhYMGgAbmWpsNfRTZM
bF0tDStXDV8E0NnM4SlyHafXOQsIQMMOPoTmluIGPw0OIHGVTYI4EhxyB6XHCmVIp40BxYQZu+s0
LJFSC/xHPz/ZEs86IqBNEURSDtBiD2OcGgC5t69T3Ng2ygt2brduz4Wv9poe3EWNgXWWzhJqk1gz
7tX4EtXfmU4sXYfD1DpR+5h0R68JTjvYQPj/RdhHJZnxOZereHroqYTt8lQ6q5jMig8CDq9zeTiC
pX1f/1sSLmsgtD3fp4VWDDtAWaVP5mr1/W0h8SzTRn37FE/ID4tRq0yA34yYUwCtdNEH6XsTqQ7t
UfYjrqq/fnACEOif/w1X8u+AgU+iy6qxDTyJGJ/WiEJtM3d0Cx0gYK75nODM7VQ45TI0kRrNEtuo
AkWrwtpihVFBMAb9vnhLpie4V/vJPFc3oZ066cD03VE7aVd/EQdWYVwQNCE2GSD/GOas8rB36Uoo
ia6/LDfNwycjRL+/71um9TnLSwH1o2N+KqBZHqwJlm03tkQxPQ7CoKGK9KiO3Dx+rsdpDfGFQhvN
eDUeMa0+jIkcWceDrZ2I/K7SfqV8lmVCuT66anKy/8c8QjaAzMDzIjHz70Pllqzq1CmC2tm9C4rY
CRMpiMoR8gCJrTDnTE7QnORMHGQomYXjnkmya/l02TT22xAX3V2yeMUgZqOWt+j9ue8bdeMS2zGJ
5ox40Odo6tKbnAqqBNG6DpF8a/UQ1mNZmH+rgJadYyhVqRfPrZLOIkyYSAjNUG1sFf6HvD4VNHm9
RMTvGuYjW+Hc4Bu8nTiTweorLOVpJeXYbf6ev1sKig1jL864qcqpTkTHxV6BFe/EXNLxfg+CpBcc
GIHX0gQDcgZWBqDOelfZj7HcMR9+tJ2yk0p9Pq5e6VufMFAv6L5jR1MktRrnomIusuq8lusYHYoX
Rg9TNzTaGRH2vf2HBLF9LRUDG622VKcCisMfvHwsPA5I7CI8RrcWISzks4+N/HVHgzviUdZ6TQNE
4HlOKDgfk9vNL4HcFyRZhflcvbUC/euuiH0hHWNspkw4T6m9aayyl+k1xMYwzxRrvlDTLTuHAAAB
a7VQc95xjlwjq3fT8nLCQTjQyydhp16I4PNPvWFZHM3IjwSB5jzkLmtdN/oMLOR17DM7u9qtR8NS
sqyjmtLu794wY409gUyLgxwdEcZ4g038tHCSJ+LRCdChn8CpYnONMDioMH438UAh05+kLjmP8JHm
vye+ro85WmajgjgaDyXcEfp33NchREtrUXhDeUtHYkD8E8QGrHI85bDILeUtbebCO13WsQKvmZZa
0tuSISpxQp7M6i8/MrSsCWM0IKppuRXbz2KpwtfuPmUh8svVGpTgTmsNtumkfBTZ950iOMpemK2H
wEAvGsuGBFTrKJk7rK+il4KUKVPUSAu6BvMss0Z2fPoSORF+dn1nmpeMg9IEut92ZYNoMjvI4rzJ
5b8q1l4OR7chaRSdrydtnkeJshFhZhC42d+LmFM1fPSrEam0e4F2ldF4rNJMr/If47GPpMFeGwWR
7Dfoz8TNOp17NFzWKQsK7e+Q5AEA2HJOvFkFyQCx3D2jaZSOsl3pXO87lu5Lt76ptRUGr7tSP2UV
aJZJPFq1/xbpMsucOZT6KtdDwrjb1zCuglwZ7weP1nJ5BWx1hYwvto1wjqxh0wqBPmf/vzpO2h1/
LxU4qMk/cC7uNq9qo8Wsi4EV0VbKZzvrKy1cNNl0LufCmfoRn5I/wZGwJBu+r/2I5UUdPvybRYKn
4Ck552uzlFlUBP5sA9VxrmwZqhyHTURNbq/EMZyLFYnNw7VsSVmJlpLqqZdc9zJ+teUgGBEgOi4q
4xrU4poA5hmzysgSLBw6LOolGeSsSd74BPLkK0rxzCuMKPeTAIRQE3kvpMHJXOIaJrXGykkMAoe/
C+Fs0H/UnE7DzaBJL6g25aY3hUEzWtNp9oB1QytwrxOFl9HRhsHnLh0s2/RsT8/iAW80DUz1YH5Z
EjdJ5jwG7IbHjdVcIRoU5M53YvC+B+mg5L8vLljCy4a6xrrig7QppsIdEPKjLiPwkL6y+jQkdBAq
qfMqgVVMj0gcnvBODHfaoffcrQQINMVx+uvxQKeCvtaGfVJpkhzYbVecRQsvD10yn6Xx9g2sKFqw
vuSsWmEoWKKY4Hh9yinWNfgtYlOPV1g1m0sm7Neorrhojg1SIzkgNFZl8lVe3Ly62zT7OY7OkoCT
4D8330NyFuwLp8pV15+hEgHXSzylA60m2GWWK0eEyQw3xHCGDhkVI/n6yL7gYxFDuIOMZITHa5ZI
28XKvZyh9GfuaxMKvI5Nim+IdunEn4bdv7jkQCOvO0msFOjlFuC9c0RvFu472NBNYe5wUdUW/bzT
DfIeQCpT9zS6Wtc/8+LFh/QQYLgZy34kEV5YLyQUNuY+FaQzZWMr1+DuvV5Jy7xbA50MdEQZJsdf
GWvlxmju62GK1jlGa95T4Hs+HvXHFM4dhw+7GYLLQOmrEz+vsDnqXnUnT1GDQp99fMfg9BorNI7J
LYUBILQFPCOFjMzar6CsW/mmJVmTYN7/pDh3Q69AFXXjA59pAdoaTc496YKTRJbryZL6psWZZy5I
yOYKHAdcSnDOh4Ef+39+8GoWsLOPjEwDzPUIcxaGUCs/0xOE/kHuUhTPizm0tkoe8qZuF+ULLc2W
QUS43GLYhQGnUXIvNH14Xn6KqiKyad9+k/A8Rv+JpzzcGbp6rc40Inr2jtz1umsz9AUQh/+QLRFf
5TwH8VDwTnKLI3waTftNCeWuQp4RHHRZ/zL9HZQ0APDlwbauFD7D9jQGuO0wjAFFBhtTuZpXEnVG
AS2snCrkaasxdDfX2WjygDQwAMEavxrfygZcdakIIHNrtETn5FC4EpSs0fIIA5H7ZDS0XpQLdPd8
BzP+Y5bY9sGAh55vrD4XKxrRu/uskwXCVKy306qa4WQOGNA7I2DzVdLzw1Moy3AqmXy/3Zk0Rv1X
WMx+Vybhrxx6acL4G2FUl4nsCVPgCn1Y2vufPlh/0Anc1ySDz3jxFh9OWJw4xk7AHun4nQOeAgJ6
2tlMwDQQLEmOWkDoZ/Gq6+6EGPXHSiCPDgLr5enrosSqzjqFcxxxhZ6Fm3FAkpjL2K/bvbMQewdd
8eASpOA9niKiWlStv8pzaXULL2mX6lab2Xdrt3NudVD9L8J3O8Z2CnYXf2WIv0CwX3hz9zqyyjOW
1jZEIa68fRUOSZTcy9jr5fgr2XzEsPrfER1cJLcjIIYP9QoZFSVvHFKPGwOH/0U93XbtcHQtazvw
ubjyjuVu7mLEWFLwuMIXyISbAkeNKS0Zs+j2acwDK/EAuynovb6gbURwbWtLaZoHY1QO/pIk5cdE
0nh+tkgL0NqMfWm6tbSTKNfNp5yjA+KHUacAxr01YpU4mhK0kFUy2tTqS/lc+eF7DMbhoCxZ3N5Z
jNLxdoAd4bYmMUNVj1uOHWsJtRxMSQ/0TQcVuqtSK5OACiwVBjcNKRb/loNFka5V4uaPsw4NB8pJ
W6e8oM8JzRrIml/gHbOp0YCS8tv4bKwh/PIa3gI7gx4PUk2qgePkzEByYrr94GGPNVEV8I+ZgSwv
rtdac4y0v/NsUEYOq0kPDOdpeipPSmRAun6lEOQri8FTK+Yosv5EHx/0Oj/IZ7Wr+2SBXKVX86Hh
2X+oEfJ3ODa065RsXQnuW/DuqSQG8pT/xlHXB8w2bNfiRFYDGEnD0PF/9c8SHIiz58Y+Yh2JO0CC
kZgOdgbO+NSJgbQ4Ak2r0z2WgKoIHCb/m9u9I6O2+BrHW0TRq1oOcQTDE+WSJojJwUBrMJB4K2bw
y9gQBgKKEI17Ox/T/xxwr3Fq3gv/cSOHG0EmbEyx3Rx8AeSCcFyKeR8z0dqLFcCUBuOfEcYWg5qZ
u491JvcdUtKK2Kiji1bNgs2//8QIrIAtgfPAAVR455XEhv0u+bavA9+aIfZ0GS/TmfvgOPq9IZ6f
atDaTok5j8AQ9CTLVak1aBNgKTMQRvqbRtlSP/2Z7szAAV9r0HMkye38GTKB5zNQrzS1hgg7r5Eo
ko00j8xRL24lOGsjdEnMaazJukw3tXZYheXJNB9h45EOnED35v3650Qv4Ku0ifXqIxw7bx49x04f
ab/d5ZhYPa/knKuS58f0IsViaEwJxJe6yPgG/oFPDQHWJLsT5qDks3dyIbQ6IE4duv8Q1Wz6VdCa
9FUZWL2Bw1p0Nh/SRXgrbpw3/s71OC1B9OeeIK3tsaMT0ccgWHR5/NaCkxceN6C1BxNuZWNOER/P
CwcWOa+ZHMYEUt1tDfdAATHedkS5w87FBoYLVJp+TYY5xEqJwfgkCl0l9N8kALJuIbq86hCsf5Wj
Rniq0LiORYI3iPBB1fKQuj13IJupz9CJHA08MNx5Yk6hHdIyUPaereP4tXKcVSlOPYDD1dQ46An1
MXEC6P3r4clSJg1Hl3cGY9tmI895crcQBlUAL7hANVjdwuBd6br+4SvaiZnjWQIfy75cw3b1a49E
4lwo0tPd4kOLKr4OMOVEKqYwKzT487036tFcpykYxZqGF9OounLgyEx44VLL0jeGoHun5iSJpw1r
YJlcGCMalwoDHlvk6ot7Y164Gd9u4DEG7tgW6iVl2v1U6SzGL3SCVy2pYiEXd19aWcgCr8Dl5K0A
RfbUPdtTkLVOieGDqgMLOCD+uvhPysRoxf7oNfk1JBHfqs/yLwM5SlsROY7tueWf7kguAUgoFYmQ
jPyhxZJD47aMja6HZrfGN+0pYN0kNLbzhL3Fislts7N30eBvEDb1xBz8VyPjQH6oprw+1IkYIGRt
NJ0sYDHBfpPdUOdcwXudZJdh68FOeY+nXF76FLStP4639C3YsHAkCEipoPLielg9WwAHxv08Fkd4
J4ebYkPahix5MSfDdGVj+sYtq/FQTMC4GjLPAIMZD5khfdBvxrGdXwJLmry4nGhuE287L8tkf+QP
Ca+9du6iJMg3NbR5/mh4RRkBOBCChSdd8NJNwneg5vFfT7NjScRjCUHqvkq/E9+FMBgjAqf5lRGO
ew589SyzPUHx799vYorX1Y/cCueQgEvXvMjlMKnGY32CsUNvOSAiHW6amm35UdptMH2UCtFmd7MA
/Fj/PTYuH6vpRHO9nPBXxF34+yhET/OevWdDcqg0w6hFxDgNrN6XcwosqP1DN2A6oWajVmvGs2Ep
xXzAOPfWmis61NibptoqpA460n8Di0QE8BaoxLZXAFY1KjN/5DH6F4rBbtfKX5/6F39WbQFi8+cX
Mzlo5YQKCAzf/T+Z551LDtPyiwMFM1cD5P8LRIRN8B4dB/sTIDQv54L/HJZfFyOLbkCTT/HEfH2S
tuT2gGfqDmgY9RP0nHuZ/BA+da4GCaz8a7u2UamDSZ4G2sIQBiLpcm05WdKv9WpadL9c5uEiEbvZ
TXUFqKoAtdNUSYkv2gKGMeiHbg15XYQ4puIP2NQLomIJ71XfngpyeRQh52ya3AkCWYVhW2TQh99O
pefjh5fzU5oVGSE13z8VvjaYsayCHVrShSaQRq3gd+WBQgnCZ9P7KrOO5ubQubsgDOKdoH5GtWxZ
zH4WJp8OgkKAOIVxLTwbsBijwpS+JiftJTJWSsv9SaCm31ZwChjWy09ei833CL0zlsrfT/nQLwIj
YpcGoJaBuVGUrf81xppy3DC/pn2BE7TXq/O00vk8GOCi7S8shzJx4dhG8QFE/fpAoslxzb46hHwO
gubIAv+UeMwp2Lz90aOuHSmYRiBqoEjHRqQ8ecPsTME2DgUHcscMKnkEGfFMIi8SWHyi18Ba6Acj
xr3rQhK+XsA/ZrURiwdzs4/shyPklaiF80Swqs22oSFcEnIImh0balV1yYKBmlrEa0/qO6jaRybs
1M0JTG0Q6IFGKYZivAnHu9FfodarE9PbENHv8b4DJOIt78jhco7lRSbhRBKHsyc3BiWnTNF5D26h
pEJhMMCB7eGAX0sjLZPMZ3gonZ8TZMwe+MbyLqYUqh+gJL/vDssNY3atfoWlpf9cn9MU13gG69OB
49gS4cQ0lrOCsDj9yd8bqrqc0Df4loEkvr83AI1jonDiAWXcjj0i1nczVvM8yoa80LKcHSqMBqVj
qEMDFcbzULOl/NdskeB3q9+CxfeLzd66NKSueeIDvqwaoY1OMO1MwcWCU7oNPsc05bhBje4wUYQC
n/CHnFKmMTs32k0V1ykgI7Vb63v8yD4q1Ee+ztTERKjFgfwzmz8CmKTw4KU3723m7Lp4+0m85Gzf
yqDuB+MkYC9dP9PjLnbOh6BfjlnCcW/6iDBWa6G9AhJXaeaPZa2Px8NJtg2bWu3k7aa2xbXBsWk5
Yo4t4jx+f+HYANEZYR2u7E+ZRUJ3UoKYfPsKa1WhGwPH13og4rZqnEFb0KHZbWKd9yNXglkPZNGo
WF4otbzaaRbE0sLSvWaysRzlx2ByZFSPcAajtjP5c7M/xqRbHqHti59LHIf+jhq2nejI5hyttUym
dxUf3drY472DuULVkJCUKQqbcXcz2aEXbK7UlL+Qg2XbcR0uqWpm2z2huwsbv48Bz3DAza2VZObe
jU2CczGrLFRqwh0ergAtmBDsvJ/e+FlCnLVEqKbf+THpInJURatayQ5VPYiLts0IOj5MalgtU+gS
JG1SKM6EsU3Z5ZHzuCx27e1W5IQtjxdWBqR1u95Cn1D7+x4Po2+O12yvgPOSVUouEIzZfrH9r05W
sQICXtcBmSdeA6+HB/50iYAFSUW1C4ezGOpM9Oa+Jji4Z7EpMpwyHjwIzvna90I8TqpuLsjrPpuD
aipRQTNYaE1LTVykeOmGXn8AhxHLmdHamA+6Jtzgk1IFh7GvUIQnUHk9BDDLD5Q4duXKw5c8FOSc
nPhoikBDxUwEXs6VQP5wrXb2xK/MKB2FDklbkaJUFGQSI9MbSaCXiL57UkYGj/+w6xIVzLgn+R1M
XmsAGnpdaLb3Ua4ojl5PZTs2buMmq9xaFsv8AO6W8GJHbb6rGAEQzvEPGs7iPCuhhyKmiQOahTf/
n4lFwW2L3IBO4VkujIHP3v7jFwQEDbxmSH5QkhP5Ts/jWsjLmJ8iXCkGOPAyOikSw0qutz5RuJ+u
A9+cbMe7N3/9m4R9ReCJ7d8i423uHnkF3Tt8YU06UHqauJC313kELD8kEh3KgGGJE41+q3KuMOI6
DdZkr5OEt29NplA3UZ0zOkcszEwZggoERTSNXgxQ1RU18rs9K2WLWuglUbH9tfS9JR+Nl4M/3ObF
N3rjD+CF2Qzj8NK2n/o/0DMKiSsOJdBAbifKMXO27kqe2+Y+RQTo+yHOoK+dW2AOwVWNZFbzA9Nn
Eml5NTtlbtRBllDIKb9aoOzZJGaxuCR8yndycxYeNw0bvlYZrj7b0Wqw1Noji8zJ9M2ZI5OveXW0
ZD9DPiFphzNWjZtAcm5W6xQiHAI1p/CKOPDHQKfmkYtp9OX9UsYDOyzR/Pql70KTG69Hhxdmd0hX
gBgvr0rwwaF7tz5GRAtwfSO6AUxc+bdbnbvwzzjjd6mC2knPEds3K8NtIYM1BYWwf4qSJ4VSMGqn
aucHxbZxp5rle9PoWZXrHYBU400Ff4SFJXRSQoBOXQw86YMXVlKBllUBBu1xpTfckw7do12UU10b
dtw5riY4DsaQBorxSHnmnZdMKGBxzsKcPkX1txHDPxZBMWKPj2dSK8EycC3KQc7fNHuDMNrBbl8+
vroD66B3ZD4Sb897xul6yKW2kyF/Zeqrk8xO8W95B8BEvsfeUl6UxSFRILy5qwmnUppXbNmedytm
TpSaw6UGb018NL2SQaGdmR9xwaSgF32frIUHwraQ/BM9LZLH+UdjFZHxD84GvGCNAXYunhQ5jm3S
GtiTd5VOz+l7od2satD7jvEZ3rTV9ELfpNDf7CMD0qCQQJqnzb1yfp9f/3eCX5L6HWlU9EGo1nb5
Am6s0xAdKKfy5INHTlI8ybkO9yu+gYf0B/RPeNYMhvUqmWIbM8k3tkfDo4z6p9u0WDf9pw5nIVOW
tUXlPuA0Tuph0gVCUikxORW32v5zgbPjf21yDaJE0KrdpzAFFsOCMwOM7Fku70W0wc2p6QyqBjvB
tXolm66J3NZRItUJQNTG6IoRMGPiZKsW9uf9tzbrf8IMtnCOH1wyP0a4mkVqHw7QxlBVSiGR7qpo
/wxJR70OpIdjYSvcXDaBjQguXgGFvZP9+tuToO/iGjNftWpOxGkfquHdYtl4VgL4UmSoC4kI4b/k
JQHBAqLEcg06TFKWZmRf2OrpbFWJlF1wraD0eA6L6DAY8QqMqG7X4NUDfCcszGuybPw9dpvrHKIB
4g49LubIlMfsy0p/K1gX7ZMwQOGivaWrfpu2j0Hcjv8ihTaNJggGf68/sIl8ceSGZ8/KwE+xxvt5
8lGsKhrPKbssZFBwJH4+0Au/1NWtlv5ZKyI49FzZc0k4+61HRWbiN06P2vKmULNMGkHKmbGHYhdi
Sv3OWImjRYuF17myrOYEMAc6q4yqcq/TLahgcnfmGCkz3IYltXuUnvDLPTUH7wB+CX3vMRaqEuvZ
X9OJkouohve+siK9W8fIQkhKoU6ZqRhdrFOCQ024IusQUOMmbsHTgzGOLlItvqPfYQGDaT2vlpN/
sVznKOfEIe8TVv0jfI0dF3ljdiwWBhkIlTk7UwXfIhfugtH8LK6jhvRjOwzaEFq4SsHBdyZu/ih2
M2ZFnPgIXXDX3x5C5h39A0kCHykoWuw+b8oKYN2HHad+mpH1bPuz4KUVaMSUvRsfdmGD2jxomHX/
iSpzu8KkhpLXB8SwzdQ2NeFARHgoBon4leg+gD9cfHT6/+8IohssI4Pnr9+TcTE7Vmb8ewa5Y7zi
eV5YWfx1bj9Y7fZwPWt7GJonZ3lOGCyCkRkDw51QEO34u6hpUqStAQ9J0CwrCy0JIQmI90UJODyC
qerMLrsk0Jl/mGi9zeuV8XtNd3nBG1EokJIK9gC/M/tWpi9glwGPipU9xm8G1R5AD3VTZ2FigITk
zih/PO5KUQfpw7PpuxCH8SuS5SDotvaSK9ZnFpc0/8o/OE0MX+7/hyY7sDKPYA1qx90T2GwwRDfL
egHPBVuZnpRFqG8GPw+QKrhc7BOjIuJB4wYBC178Ci90yRN6rXZxJ/oHCRAJ33UOib8qnOjZFs1P
talypZYQS3X6U92Acw+t016uPp38UWgpS3HEvJ8ZaNOIpdBru7Ovl7yD/XjeZ0+5D0OY3jn5NWpu
Hm5vjRNpOXLh6jNFNhdjF5fvnr21rgUN2wfAPyfLgEg29SqZamKoFhc14vM60otoJ05hXGzcC7f2
aJMklusQdDRQD4r6ztqQIGfcW/N1r6G5xrrciyTKvh4vMx4kJbTXtBVyzFKSb6o/WYPofVlV93TO
QwqESfMoCNdnVGJUaw1kFx2OBU0QYR58n6pQQ2zwduUe1zxBshmpTlZFMqna7n3osSJjrsdZFBIF
yrDBjggQ+wLLihAbxjer2rS720phnZ8jWgGoUWGqqq33eoodmmEpFIVL7yojp/9xWxjuPsVJWzQF
LW8mmgURdXaPWAyrOMuKPeeOaI3PGeH/AVnYcGz0HyjbFJvLIrmQAS58hr7jAbvRBcmC3cP5ZdgE
ElGIR54cqhaqPnTs0QnWKQHjQXcsCgxPMNvy89t2/JGoD7Sf+qUnQsyTJsylFdOLv02V+qtwnfUx
m3DMZVPhtRqXuUZgcif42ONf9W06uUPctmaqBbUvl24rDph/iWCR5F1EnFafbWi1flLSNC+LQ2bE
mMtnExh0kKkEKIjHEwL9KZ7JJsBGuU6FZWHkgVEzjmb/rkCpCxEXbM8tZHQEvVWQbyG5hd+3NCJG
l4w2p+wX6mFE9YcGuqCRn2teu0VeTEXRteYLMbpAIe8mE1VULMdQq3wHjKsptLOOUVmckRgT1+Vq
nJ7bmxWJ3/OQKP468B42Ar8yDdeO3eT+lRzdwLmBx2UVchgiqh91J3SYM5+v0ojvhGIVzQSLFPu8
5wb0rUl/XTkFN+Pl3KP/Jw2BMoYJ9Po6vOxPmFTKDmnXrrFsr2UekkCAkb0x05slLptVjl07VmuK
tyl6s6fePPP196oGYtJ6qb8MITPKEtgmiEOnuHy5v6Ftf7bompDEMwlODuAHoF0CWSu59waiAZjz
5JXi79t05mqYCe+zMYscV0RqdoCOeIEx6wxGnRmQzQ+7mKLYutzXrDGbKoVn9FtXLB2dTATqmnrk
nRTIdiMZXZLq4ytZOMFJ4rAc9HnJnIH9b/wHUjekBuFENCx7nO1JL9CMfb/gTfVLiqaxt9QmVNef
pIO022elI//YznpiltktoR2Yl/FAzRQIMB/JGvduX8iF63hIpYrRb2H1KaloVDEACgGNQn15HdKK
C49kc66P2UWTzgZaJbVJ+ekphLTX9EDc1lOikjwlnfoktsBjgXdUwX5BHNuQVQKC8VJQMb7717Lq
korkMVIVkCz+yiHGKkceealok550QCZPcr/ijs/FzlQYcMeSDtFhOPvkYgHqSK/bDubqRd8tLX+o
6xC7fWpQJQluVYe0pHX57f+xGgrYllDqB62ITm7yMRMPWVXCwRcwAKezPuE01m9O2ksfGZRFr19N
ErJt8UHjlTf+gahYbNfrjyIrZ97mAlWFFAzc77pBbY7YMdNISZf8k8fi9xkdq/l8RwjWYIijdJlD
zK7cOW7a1QuVKN+uuDt9OP0utfCgIgkfdWitdslT3MBrroiwtQs0NOmFTIjL2DHRbU7LKhyHaRFL
p5UTFRnIUoMd4AOIETzT5v1ERBvU0RbvqWne/BN7mgCWZiC5Ur+7FbuP6TxLiQYBIEdXWjNbFhJI
GSqA6xUhXSqHEgDXkzW/Ifl4xcq5Yb4ujSi5RY3qF9ugHlmV1blmk5fRInK6ahWYEXkpSm9aVi7g
px8wNHPtlatJxgsznjB5c9DeOfT4EiMam1ITxzYk/DdLZrHZbItvS0WtbC7It3+YQLY8dG+DhFvZ
2Zb/yEkn0Z0PWGyxnflwbCAPonyiPUQ8LWiis3u19oBBUlVwRolc3uotpohEco73MSRp5Sbjn35Z
0RS9P4kt7PILY8FUWpMBro9cIm6bTn/rBMrZradpQvqNjJbLov+wEJ3AOkDqU8sWSdUf+aFZ6ewN
/oV7HjCBx5Mfvrn+fD9I66OnxHSVUfj1ogaHfaiQZYE0j77SAHeiWTOkmoWpNxvtboVnxiLt482N
miEurAXWPK2TYUgZk4fpR/N0fVGiET7Gv5cG2WD0sdNto2vVvijQejJqR6wJXOI8+ZGj6AHr9Z1j
crr41Xtu2YJG9EFi3PlmJwsmgdBpl7OOeaoECDoTdj7ZS++Lzqrk3OGXf2K7jxIacnYET4TvjGti
Yxjk26d//GSkPayFiV0wIgxTyOX45UAa5kyQw8v3oEM9Y7r95QXOWRO90SAJWQv6bDGYr8Mh5z8/
W9CHeSr2QAAxml2LgfriqNftGWtSg73djWzxTjOd0bxjsFP+NGEvED9u5BwHpruSaAG7bLuu9a3U
Z3ODMC16XPsiP1j0sKJ2JUXIfRzs6iUbYYvLwnqlX7UE3Ds5uFppDAoJGsb984z/UJIahbDYkJLx
9YKnKX/XYn9aHbaBozFm5yduXww3w5OuFEY+Ya49+nR8ynnFDlqV+pEgMHgR8VhCzL63eTXVxK/g
53W6/IIrjCI6DjH7TXZwVVA9LrB7UmaZu5itwMRWOSO/f4kJ/AAvoNFtS501dcGek9I5gXumvR/2
xUBCg8r5TRx081aIal6NLgpz7zBilR6wsuiq3rDZM1T/qdrCVTi5e+tazy0p3uSipTasAb2ZnxSs
vv/I5rZC1kICThZsEDJFdthYuFzoRhwXPxs7LFdSSdwsc7mWqlNqey5OaBX25r3bYkioBRZCGMB6
s95Z2L/s9xpuYduwyeim3NxnwOTwECSnEtRVwl9hYEh8SjZOM0/xeCBcuiC+mP2hQoOWv4ckj/Un
KlWMjrV2zPiJgnikJstLIpCGeita0dJBwNnNRZtCg3EJj0Mpp26Qy8KOWYCuORK3osrK1Jviz8kK
J2x8v2HzGVTnbHmeKwBrQIW7aP4bNRJbTiieAZHyM6I4B/dwQ2uL8Iu5F1awyCfOHnkOgmj6bxl9
8Z6pCx2FL0Iak2LVMHFIW7moYd/lwkBxtJgvOmJPAaq7t3dpyOQn/8Y0DY/RhoqpQaTV3FIYussZ
8mRzJlmmUtUnzRYfQxAQHC+ILwMM/NtkCd0PDQcdWPIyIIYBF8vDurVDVtojSoss8BMJenlbS3NX
8Cmk97PMRuLXKwoSNhip0nR9jA790SbYTN6F24eqNqrBHgOavEZrcGTJcnO7qmWylj2IToblfSTa
DzF9Rf4Ovkmorkd4boWRpEcKzMOr+Cw2ZBSIHFUBeM2Ht2DYSKvOhzHzMhk6+3a043Fxyef/j1xC
nyGoKNcHYFFDjUn76mxICORrQkpobjwWID0az3TH/+s0Al1Nr3qJJ1G01OGyfARV/alVb3E71V0P
bzJyT+0IqqD3EbkKrtUBVz9yTbeuV9Jj8HzmFvT/jREUDK9H+hQ51vbs1ZTZBLUMllSIOu6VoEAf
MNIfkcJsaPrwfPR63PxRamM6OojrgfHax3/dKKB4Te8oUzCYjtGAru504fUcWapoC2fJxRjZfpG6
CX+BKDE5Bn8nWvDjbB035+bf++XYwemoKPh/p88JzlJbO/l20GyfnLW1XbjWA7vPI9vxJMm6AjSK
LW3oPcs8ybiwzXu9mEd7CoZGCIDuTV1TqzSyQGCMGrQJsp2KBTXo1n1ca9XvdPjKC4WD0WeZjuYx
GuJzAV1g6AX8el1fsBwwbBhYJVkZ8fR7KNGfs+6HVwoLbSRlkeuxfsIekk+TE5AtIAiBneSpyrCx
H/9PASF5f3BH7o7wn1SgnTDFNoU3fl056A/Y3TcLli4LhsHjddt1j+jKXf7NKRwJV7K5ycFgJwpu
gXhj+6PBuo9SQ+cRxDTFa+HeyGsD+GqKV4Qn2aoOWvXwdq9KB3dXnPKx/k7blguSLqeBZTX0YYA+
DaAich287bPfpX1pmX8UPeRb/p6N01fillBIwGOmx1cNq3v7gTN2T9qlmLoXLdx7Bif6WLGlrelc
bLfJf8qrMQiY4Xtzdb2iU094nsDQOSQ+saIDt6CFLPP9c8apwy2iPRhJr3iojkdSZ+B80F+7l7O+
gFLAxEuDZU1c6Fy0VB8ozjl/0i2OK5AOZIBeMXe/3hUxd+xqtaKvn2jBOOJ0NvW7Lwk+W3CcURjJ
eggnlvr81fb08wUEpbeagBkxymkOELtsVjWW6cTWXg7RJR8hQb2YMtJjw4J6rMWXTE+5ftljJEqc
G7BX/iJeLk0s3y3JKK8J+Auz8q4hFPDWSDwhNXaQtfOP9rUXI4YaQDi41cxfdI8ooabCiIyj8jnn
GWWo+GP4n8rln/mXkfGsIZhnThk9/VFZiQWFsGFzz8SCZlUKLyB6pdgJZQ47qLZm4ftycvsSlOK4
kqH8LYGB8ojET6l0WjKnbsgM+9z/cutt810S/FL5xX/upkrDcNe5wifboaoewdioK+M9Um9ejXC8
HmBEod9INxo7g0H/bO6w36qEdOl4WBV3qYwW8e29kKNE3V0WpYqy5h18fNh15aeuYmYkB62Pf5Ue
Hwc6/cBOyofvQSRNKt2XXwMPJ1iYUFZaV4LzZ3UItXVLGCTceFiCc4icDnXFMX4+psO8jibMv43F
NsEz8VXhqwy3MzO6CwfCHP8WDT/+vEiBxIAkbAlIJkIY6dc6Hc+rrj5h5m/rdDNfdK9SPl4EPIaa
7+Y7QitOXO4kcRVnJH6j+zdxKVxYD5+hf46Tf4YyBmbLBZm+AqIZUvW0F9138ANKxXfyR9xHJQys
nSu3YqpavtsUGCsbVDYxTNwhvUJuz/E3CBNio83dWrn4mzLXPUV2RtnFSG/ZWSj4tHwDFH+jINj9
OCUhiQn2SU29Xee/m8Ip1a+xBzTwpFeyMdjXJJLF2REghylv/0imTtICE1nkDNWaU979MtBrjiQh
6OASD8fvVYsoV2l6LoZEve1lNNvEjN5ahtJFnU6ITuuVtGTncaW5MH6zg5aLsZwaJ+3wwaRlANvW
KXnIbN5QFp4xYQPsk4ddwxTFE0oaTRMOBHe7WS5L5RJW/wEby+km2UPOw+4BHTuu/annJbDs33Ib
ZPhmPZRqdDMB1biU90op9AbViBvaUG8naotvAS4UTbLf6I1pZducgyUG6thhSYc2FGzpGrSdjR/x
kWg2VfOvM9zb19YmPj2xTM+5d/IK+cgDIlLoq+RQSnCSM4pnMzM1BXe2d3qs5jjS9AUtw5nB60I3
qWLBh35/APK37zhaVpVeZuURW2Em8xZpH3raGi6tNvqkQJjnZZbFdvgccpjkoHv38ObPSrovgFem
QAyNZbYcZY0wDoAt+YDBCYyDxJ4HgA98yPRvGsWtqGxMr8S0h0Qn0Hv7cR8ST+ayqsmveOL3VnNk
l62V17Jh6eiEKXiF0+2N9QMgWvHMSNSpXekjlqyDeONItXVIuPPPVQj2ATRjLHwHvE36AfqCuz6h
gc84yMII+MC4+U78IBQw3PH2nxJ3H8zAGfJtVEAitaDNEoy3JbCHGDgIeKOBARSbjboz2xx7DXoT
MsXPOCKuMXiC+sKbAdGVvbxjpC898m1cfoEwniech5zkK13o35qc8Py3CCDdaktSHRlxGx1f1Zck
MWxi0yFmiUjytc7gtiQJRf2ofkuFP5+3GLS03ELo8q7zJXsbDqUIMEHqgfMG6tJiGpEyCG3WhEJo
pCRuMoh2lfV++twIoQAaLSWVVijW5DNyRyw8kQZXhEege1TvrkqpENmEPf2zjjIeOn2x+GoQe9it
mKVcQ6QGVcZw2SJoYvqIU3fFPN1i0uM1N7Rs2DLTJTOx6kmhjmn+H90PO94G4J+z15lD7jpmGVqB
Yjmp8iCUAY9MfwLm89cNGv1pc5KeKkfuyKhaRwS747HOvvdSeF4ZRNbA0WLgo7vPCSpz6M9kg7CD
rpMmcjS7353vvNQVBY/tpmkEFhQbA/l+WeIdLehJO/RfXd9Eev70LCtiNtYB4RBs9oeXrPpiM3GH
cQLQxWdqe8DVh/MEC5in/DM9URRz2b944y4xBLXCa/8/LQe4Xh2z25YVT33HH51l2/H20+4TZCVA
xOWkFmPpHYyFAgT/MR071/GYzJp9wR3+bs6IIOXMgnA/oSJ2t9DUFCeyaKeOyG8PnhrYs81/1o14
iYQSH5vE8R6AT6dgk01CcmL9ItuGKTF5ll/7uX7/fFLwsPUL3JyWeYmu41mWQgV4alhT5uLjumgB
Vjh9lUdGHCgatU6Sh+8m9FF2tX0AC9F4MnHiWEyu0SSdT+Rk5KCJBvK4roEt7MqGvqxCJ2JYoSFy
+euqL1Cpq+Sj298LUu9yG0r55zlbgGi15fNSPGn9sGx/Cb3kulEwCQU0orUk7FgfZOyGoPeFYBJD
DChneGJ+QzWs4ZszMZI7UL+uZ64U7+H7LeAX0SYsR/XbZV1GoQw0YkG7nHdboQgQreJ3fn3KaHoi
INwuHNiz11HI/exQyHebTpLBOZKAHcOjNqHAtEgJT+jMXKiMppUOAQWjEDSIBubn0YM1U6DH2Dbf
ceiWJGj00iltzsmWT6gpFWlwVenaYYCXavQGNyHrUV4JQOr8KHaCGYN5lp1e6SondpGGO0vm4CvJ
tKLnIKZ7NTHD1G/X2cIxaW4U21ViSI+Ttg0D1+zITCr0ecEBHVlyHTNEqZd5aU9GX1J0WCc+Xp6q
pwnE70MHqTzycAzWoZm9gvOVW4z10uFtke0H3T4Vn89vG9zlvo+1IYsb7DGIBjEa/NZ1IKHGBuf6
VDNsM4NRd26hnOAongRvvBONksnD2qhG5Owomekvk0N0+HLHrAAUqzWUILGgUMeuN4RTBHKJzKiY
SmnpSY1egpuIgC3Eha27CibUGRureWEHftDekz/RjZmAhv5D1Xxj5oAZhznXF+NGXqh8DOc5drLM
M0o6VC8KuyIrz0aGlygbVF/iH1gwd+MLXB9lcCfi4g9i5X33iM71/99tEB4FirUlEVBbgJtLCqWY
dWs4uldzZHniojgXmi33C7rvzPvm69/Jn2ZUiQabZBpLW+OeeRuxjnX2jqC85AnyIokfih4zDktq
kMZvTMsv4DvexPUE/lKARUcy2zkVyOyp0S2kCbUsQjvQZCHARgUFJgAAYqChI5FacnreZJut4qEK
K9O5NZxaxuQix22QGOVl0RPGR+Rn4pkw5Pe5/Wu14V6mVXurwsXfkexqZw/xULkxFvwVJsCI5T5r
gBlf+Bkr9EQcRP4quCamWP2YLMzy7UAiE4/MJITyZ6+POCVir2O1cuQwFDw0nzXRsmmc9WBmA97V
2fjyWq8QirLS+OaSpuUukXEAswn6eg2vp6yeH38AXDm1MwM+Y1NjPVAJqG+IPagKhayPr8G2qDCs
60a2UIQuUB1whDJyWZzr4wQKOKiD34MhJMcbcAWSahAPWtBpMHoUnZjleYEZXh3QpzceJM3ud423
X2c9PEHh+EFwN7I3pttaeK47VdkvBRlV6xVcJi0ReowJYUhVtM1pM0J3F5n8X2ayJ9COrMBPzTAG
ScxBu3AStsONPTGUxgjA0u8ml9B6i5bhhFutQ6Qb+xSPk3PXdLSgmnuc9tDhehb+99xNODiHhF7Y
BxaFNwYrmrHL4GLEc08F86uqt590DzMe8ZED8ij8/vutqLM8cq0jIWzT+HAn2xhPjmdYzCyJCBjk
atfwlLc4ojeduUoungr3JWOnOVHH1BeUi1Gt1uUbxKpqGcDLWUNYux261I95OmcBxM2ESd4JOC5n
r7VpRQaZgv1DpSziDeY1evgQXX0x83I5Zj58x5ZDnYcGaptlAv1JkCuOfw7H/QgJkzzXN8SSCnOH
Fi3cEysgjtW3fCKRWNwANce7qgzP71/uV9a98PeNgVBPxnwbggNBwQzTj1u9CWHdzZIzcNDnpPX7
dxvxWXBOc7VNaKX4Vk2ky+qGnFxRY8wPHCIEoTxjAupstR0JGr4Eu0IyGFJhJtdYuSFy86zuGasP
8djR9LUXimQ6vfjkMBc04iJGfv+PqTCs+vPriJt1Mt4KyBUyYBnS5Lt8qTIDhpwKAXBmxmKQkapw
SgRRXoMWFX8UqoeOwD5WUMN9diHi4ZTMX1hiBC8pnLeVKUJK0GwjPeoMe58DM4Yyou3wjv5hHbJn
ND0ccpv/ImziV6FQV5H1D7Gsv1NoGcSLiu7Vogvjy7Nif8Y8L9wEhxxnVtyciGqBbQeWGdOKy2PO
w5TLGO5ydslZ4FXCYjjaTE1h2WL69FLm3UlxlBHmiZTDRUuH43A81uk5CREWPVaXurpbQk5RBzwj
fm4+oZ8KRCUimjD+9QwXjK1lYl5SVq3n0ag5m4Dby7TMVELmTlWOvHGFkr2R85BhqFzSEQoQt0mI
uUhMehCAaUYjCb15ZF8q5/UuGKR7Dge0ooZcnagPiQLddaUFPbcMPOQYRytQ/GG2/MyjcONG9GOy
ArN83+IT/0fmfGYjlz7UGoOqgD/3IlPG5700eM9UVcbbi1bHkEzg9fuyim0nKMNdupYw8xdzfDRY
FMej2imEsR+OooYoE4QlTumlBDEL8EyGTb1ZxT+rko5P2OQZ0KOvfiqGqKwIZK8FIM0KNdx+dd14
ngIr31mytd0n8Kmth5i5Eo9tvcO8+WmGeQhXZH76rlnz72xX4jCNeJuVB/0szSq35vadFRL2kdwC
+/XriUKyzJG6Ex+ZVo6XZQG7zTQaxdSgfyQilUwdGjVYph3gqtPgv0yvqD64h2BTt9vXssyI/z+w
vVatUAhG7fH3NZcOEbgn7Hfxy9pzmFm1tHwLvNQO7t5y1ybUOobcT5r9wCAwzaGNVi4iV67F5FX7
p3bTx7nrZturyD3F7cV9kWlefbP+uteToCTOQfh841ZfVckO6azpR3Oc4WyXJ9nNZZTlnlRzLvbP
nzkC05cbACu6piVrmRkTDHdh+KzF5yq+kb0/VC6hPXghQyPesuzmhxS7uS6NPSwH5+/i/5OEBNWa
TOq++6FXZ6m5T4rq+DCuCMH3+10SUR7y+q0LepDM8htD1u5RENLL4ulqpJMUEmRAtk+yTzmwC0a+
N9UfGjB/VQ6dZDVWQ22ih51tgcpsLDmwzjuBxKBCQkOdEITc9uHimpU8Pmu6a4j2BsgcPsCQYMD0
LKI9u2tiykIuM6M181uJkf4hB8SVrWYJYkSx+do9svOd1JOiakglVPijZbGaMi4juIj4tOAuvgqE
lvgDPmKq1F4hwghj9z6Stxhh1Qa17CoBh2QjiyqKVqIFngO3aZMmX9DkzUJ1aHKbAEe1DwBITUAo
zf3f/jZm+mYSUoTh6W0xkLxUvvRQTGLNlvNMueTaMfUCR1hcej5drGCKHET+Up/PxFH+LdS3oHMT
7MntqQSROrWIE5Hgd1LjJCmlBlLNNvZC3hroPAzxDFze6uTYH/uduN68USNuQztgIvFpcYH6hhOz
9Z14YAkCtZUFU97Q58qSuvXeBz+xLi1v3+V+T/toHTxqB8z+b8cdEy++aRmTJGRMBvfEsoS84s03
gPx7fw75NuMlFY6Qr6Ga0X5Ynb/1EcXqI/9dTCPPMDNrwaU4j6U/hsJPl4fT9NCXdyTxQrF5cR1Q
H3sRAP2pL3D3mFqVwatxyM2GHeWZTLCjs9Tip26FRss9H7aCtrLNvh7jAC264AItsmEM9MK9RK7y
Vxqa0svqr1FjfDyjlAElBjl2fqPP9KPuP1VL8mLtKqOdqS9KeB9KgfeZ93rNuF96gboMdtornnue
FvRHWLWMfqb879oHV3D0KgfcCWHmxKMY6t91b3Q/MnyaQXyGDWRUKFWvM/ROjNOG84GNnporVa3W
Yr1h4mMGukYjN0/chrSkXphfHiznh1ui/168qMuwawH7K6zTk+NmYwQKZfT6JYaNgLAoQl6KhGjD
9fmUIta6sPMcpZ3zlenYP8nVbm6u/FhzewM5XB2hh2HfcrNHuYGGNLuLaRVOBJFXmYVM5T4haYOH
9BNVwDqhCb1cqkPk0pbTIqNn4VnUJi+sHBFzRv2kJ4mGTyqKpFHQk4pcqRFqhJ+N17NgQ0GrRdi3
Dl4GzK+2/RQ3F8hCMvaGAXKjuhj8yAVP2Hr+W/jpGJhK8ebHDiDdfhd9gglFv6SVtkdu4ojo6StO
MQpkMMcFcvHPt0xpC80axiz57mm581w9Usw76iSSsuaagTG0JaMdw5Jt+V7B/9CA94FKwVUSgftq
t+lwRhClITdccnM3Rzm2azgj78ZMExbcWCZo3H/grgOcsMTO6TH40EwQLsh9HBlvdg2huda1xpA4
/AFj3KIialQDnq6aR/WmeNcm+RDWFo7A1KA7iqBmclL8ydoqZoX4rhIDM2xfwmFRnLg0AfwbbpCV
n0mGS9T3aUHZ3JfLCMjP8YPwF4aTth8SyWkHO3cARR7bjcZ/X956NTHtwprTLRJzGn3YSWkH5Fhw
YJoWlpm2yMpPO72VzW1oeJV0bHFF8nquM8dGRlZMe7wHXpDw7Yi828gsqc5vF5D2dkocyg3+CJKr
RmyLtZQEjspva3o1BPYH8SYI3vtAtMcLyi6r6WTMRS5K1hmVEfBfJvfOWrUmtgWZad3Shxuo+XUB
R9IsQ/JlB8IuyOE3QpM6kCP4gimPyS4MNeRazS+kAl+QPm/KRYCW75Jgwq7Kg3qkezQTOvuH13FK
m/9AFM+1QRj43JWLDFzwTcmIraRGOT2jwOx7H3dnh4RIDWWnOgx6nA9u2f2zED2Hc8TVbT+NYUTt
nUezHLkYYaFCnx6t2iqVJmSEIIXartwRy0M/+pvYh9KVUf2Os1m3xilhwOXPpW5ulWZH4Z3cUxrH
ysG9bBFe/PM3A3N20mMYwV/f0nq0+mOQPoJxuWIBl+GDNd+75LZAlpNkobzITALd/QMEq1rEKceZ
ZNeHVwDZfz0q0oZMq7cgadZnOB+HZlUZyXO03DDTp3pbZcVWpPG+/kMl+aUYTpAtF3ehgiSuiX1q
qgePFYlllJJtkutyEynDR0hxOSUqY5p/VLQKyDOfynf5dDU7AFEWsZy5JlMJ+qXU66eG5A5XT9zs
MfvHjgnx2RAHvH7PpkVG1Ixz1e0qtuDBNfswcW46N1ibV3AZthqSm8qKCq/EO4O4EWeZNLl+aqG9
ixQta1AEfLh/c6dbIOU+x1F9YQZ7JDYFVD3CgcZWjyB1z2KPG9dTorg3hE9Kgy9C25c8euz4aIa6
SSbXaIBhwGpiVjplhWiz791JLmvWzqcppJBRivZHpiVUTzsznpeTieiuCIJFIIwOxNr+70LWnFOq
wlZiH3+1kqFbqnv+J9fI5o8LjRVrcojVhqcU7LMxeu8gq1avLR/raXUsnihDravVhzRdfvChb2av
gLsA0shObZF7vBSg98Bcf262El7KybdBevOmBmx6+zTyt4KsuFYkDOUMdVpOUzbPrsvfZ80cwCtF
79dznIq5REhLKzqjbzd8HSawtELn4kRmnAQEpxb/S5g4rngbkeYVcNYTPIyBA9/onKsXPaMAUtsA
l2Covo7zZ+X4QNnhHeWHjYHak7qVeG+lXWXo3oehSVurpr1T+D7bEBt+/uRko5GaoRYHnH2JU99T
8zS7zV5sYqNo4K+27EcFFOGQuDL6a/76TC/P082yfH62DsjyUwEl5u9IZzxaD1IRaujFyE0p3K/1
alc3M5+eeSFlsDtjjdXBAMVldT2Q8vSQ5AmaF9RBPhvzmVDP+J9k/NW9NhCr6cds73R+VRUtMW7z
CCe7q0hnqrfb08d/dP4RtdTx9sFnkivDJGaQ0g9QXD3gLnybBgpFIctmJPSLHhCBbNCxAM23cHjr
gi0e1Z6utRFEDxr5JDmqY9aItZqUw8Kul6+vfxkToYc+af5InSOj1jLcN91JWwHZR3Y7Iw72Ho5g
JfW3OYGJhqx0QGbrUahIt4lr9bMHnwE237Tvx58dtjx7PkS9b57Xu6RF6LJLu6XSICGwUmjq9r5R
fmrsRkF5GBzwYGNYcASYX62YdClz6Nh7/iGP+T5D+VIdpYp35rC9pUqhnWjOwDwPf72xVWY9QI50
U6zKIpHNnqD8O6gdMt4eqUC0jk2kYCVvsdceDw9Ja5jTaalMbs96aJgt+e8LJHT5jRCSVIj/21+2
lhZzQNYUoM2RkofHZuvwXeEsRkhnAbeRL2ALuToMZ46kC0KU+lnTbycbYsG2YH+lmMe+xeLlAnV+
PZSnUHWaVAtyd6QNm+uuf2oxIo5kZTq8oXhNdJbXHUhRufk1S5rfG9VyRaZf+30VhczIELBH2jV4
7pWrllbpvI8EG3B2CSipwh1D5uMVGqGNGYLuHnAQGqAdtcvRq+avLdgTSup5yB2v2T16mU0EihrB
R7TuWuF55TRydQTSjJngClsy1/GcPQTqDSQvBvkizzNXOGv5lK1bsLJ9N6OCedStAbsJe/9Ci9Jt
3fRrJB0O8ZJ3armo+rWcv9QoAMGEiXx9sMdkldpkpNwsPXSQm9hK4U5DpQrobUI/w8GXP7VgKgny
CXpLd8TzzXcDUIswNF4xazhuMX1vJlMsq1rK50nW4T9K8EacdGBYFeXFoXHTNYm0mz1y6cQulQVc
rRM3Ij8jG2W+absNjte1ITX18m9qREsjFQGrFxUIa0yU9BlZ77e+1YH8NjSxtw8f3lAl9S6GDxgY
zLN+WVZM2UjzKPQGkqZUxfWu4OGkLdqoNW4BW39vEEm8DHSuLrhvujwMIt9G1F83YPpGXA00ZV7v
YIoa+1bd6YfZySFofQhXIUgwBh07/RU0wW0zSeW8I0gIQWXtEw1wL9FzS2rhLOzAuXJ1rNCKUhsH
svck9SMtTKik7dOCOZYZI6wT3zKvXHzFr+ww4JLjqBf4++QLu6mWLxG/A9k1DK9BWTA+JgTglxCP
HZYIP6zB7gyxpPu3KmHKzo8x/xj5qFGwBtetULaUIEuTErDIck/zbM40qJEQmBogJRIirfQtDL5p
Idvt5zHJoStZAFPz3zaQfXpJn7pN014nFdOkOL+qys4N6N9KBksDMEwNzs1QIA/gVnJ2qsO7ItRU
1FtSDtAIROh2bFUsrD4iehKTFdwxctHLemGOPUbf9BCqId+4gJgTocOf8jmUyarz93J+EXZOWBvd
QvYXrMMRDIqyKrd/ypdQoN7fDod3/Z6/69GLtlT4YraiPaBkHnjjI1SpApSclCoXCQzp/AUokc8I
oyyOELuZzmqM44oPc9siFW/mQO9uWP6JKk2NAQpN5jORc+YPiIMeuIKas3vUaIwXhwoySSF+/dc4
GX+2bSBOhL4696ZexyjlmAhoJbCho2VtBd9OjraxstXt3JYmbAOWe9yn1xDH4euel4JFAtSSSALH
6j37v20M5+PO2jAJSpLBH2ltjiS4CAl7s/WpiMnDPC7ChQSFoUnwPDLtsb8OrHPglH4+9Es1ViLw
tihbf2fRwfIKgwyOC5Yqy+GNuuENBGjJhqYS22+UrAwaL7mt+UZMI54v1q+Su40MkrFxZv6DuTUO
WzQ5bSFDIhhDdhygr0VYcC5xGcjXcw36BLlr12If8SlZOLNbLw95ZHPC9la4cKYsJ9E2ibGzdkjH
rWsbImxenRvB3Xt83JH7kfyqW3+haecy0u9URYJDONKa+PNA8uh6WaRwWKVsSmVqdW70FyJy9R+n
0BQYLreLKUTWXJZkZUsGQAwVlKaP+6PVWoRU8fLMPWWvE1GR2zS9+R060U8aiA5EjgVRVZllUBqQ
fsJ+14B+NQtZ5k/y/hmemxPFNmp9evpGAcXP6WJ7+t/x82fZCZsOVRQCWWxz//qgJNxcIkgcWuO8
Lskxjc4ij7A7sil4+KJzQJR1FkvZ7darVKhKfx52K9kKPqANrP0QymF2WCpz136jw3X6labcG1bW
blHrCakhigSzfY8ADZO48S+trkPDZmlpYLwthqHClyP01EOZNdOsVSY3pQzU0kZm9CZEfG9ujCjC
xOsd2V9htu6pZ9R/v6TcMW3kOImgb0WnGLNDxTONvS52P470xwUqSyF6ai0u/9QlKyQVQGqS5t3j
nG1vALDg2TYgbMuaWLFcuW+CZDcIfvvR2B0LzNyPF3qKeMNFn/Z5urfk5V1pD61CJ7GEvFV2W/1U
1KXS/Id04pcd6Io47Kctky1G3a8FheLZrOY/QGWFgLVyjkBhFBhrZxZEwqwp6Xvbdqxl4AQpqrb2
fqDAyfywRke04eCv7HN1E8FY5V8z1VTCQNXNoP0izWG87Xb5ovc3N+JmYS/MZR5lMdkD62GREaTr
yz28UYbrVNIQdw8OxzMRAfZX8jXT2nPN9IxwDsPXKNxwXVSQhtukaeluK3ZEiKegLyTQuZ+wnQSU
AOgk/bnwYnmw+CNyPF9gXq7pFE7tmvQyrGpbNmV8deNIISFxMVRdagh2N65XDqaLkt2MV82XkAv6
NAVJ08CO/4Ci6fbhV5/5DqZ6qVrRVwetdq9RXFz7LcBidmXV4rH7Papg1RNRn4PJDyiA43dWn3g1
L7oUf9S9i53VTNba8b0+LUshHmnBnrn+5k1hSEBOvVT0JNlBtosO/91pDGp039MxuOh9xyzRZFsO
xpHqC4oDY3hg+05fRJsqPyXePuSyFXVP1a9wGDQr91OTBH/46l6JdM/I+O9UEPTi7kdKwSDHY6NI
9EN6Vqw3T5IBq9tj8ASz9HJ8KDnds7/4Q5Toeso58swYMhn7e8LMpGC71hjlXXNjFDt156+4gCgq
XRfdxv2N4AxvcwXyxq26bT2YRFN+WNh8oXstYCluxTVzg2GreXLxE++Zvy8xZjSQQZ3Zro8XqkfN
5NSa1/mbUz3g42hzsEIyW8FA0ru6M65+BOvA1710PBwDAVCBcBojd5hS6qBvhBQAleE9p7H9r9h3
/ghyGwiwLfEjWK6yWLV2r23jRyB5+q45Oi1IMrvNYIcwiDLklxy/cJxn+swlaJyBiHT/YL5QDg2t
brOBfXBokFk3T6G3xtyQ2fs0v8CqI1fD/Hh3wnydViL9p264BN5TicgjPzb/hMVKVBGX3w2s1vZM
8zz3C6Qd/qqxuNM5yGK2iBZKFeFxV5MBBfGQPSVO5rSq500w8HWss5VlzbcEzD+NLAF+1oRDpc1I
I6cMfExQ3lBh7Awo5Del2plh0GfcRUBdnnAdIyJLXfqe9CgUV0pX1ATsrevbF3wmtZDOJwHljFOH
nivt5AaCBxWQKzZwz6yF3xTGtZ7Se2UfVX/RJz5OVnSjfD1Bgq4+a/pcj13dyGLkpCkZfHt+/2S8
BmzeusggYtxFQ50bHwZjPTdz59MO4RGGeNZrKWJ2SlL8Yj+6pzN+xKWRD4/JhLY9tUmqtfRoyV65
B+ANHTgItsyPEx6TGQUsycOMyFkuqANaevEj0X0gUOnpLpOhTw9VkbnlXjjD5ooyIIB8VCQ3lKWH
givSZ0fM8XpcpDu2gPzncZb/Uld4mUCfXrE7O6QMRxfK/iWP3V5qSSbveutFSc3VdPkmu5tqhV4p
jM6emFAtPpZSHB8iXedowAV0oFqnJuL7+sqJMObwABEujTHjC8MTaFAxbejeJZw1E+eYO2tov2Bf
piycbARAIEsy7BWGXNIQwFIGD2w8Q6IZ6nSH9SzVLhN/XUsxuq4CdykeXGqlBRsOpKWVgE+aXejj
XgN4m03S+bIJwSYRtXWNEYyTS2UOJ89lxEYkd26Aa5cfQ3vxFsjzSN5LDul14cIWBVYqCfJitkRi
c8D1o2EqYOIORDl6Kj8v0oLByW3uk4cp2aKUp2xBrJlzQCUxcsrC/ziZwxIw6eHrcZwPpWGsD9Ys
Mhl+U9bkyDBJYRCYdMs3ltsd+iK36pNqDhdvW6T1Dxrbg03Hum3oHd69njo15KvzSC1IMStz7dBM
h1H+6jYJ1Df5yOOcfW0FJZf60gZ51PS8w+qhUqpyD3+jJE2oj4yjR7M+VvjrUbw8f2SOJMYKmuP4
xvFT2RcL5ahZ4gjhcT7XO0CD0t8r7aSnVjX2vD1ymbCM3hH0/nPxevq/h/RVz4KrJagyAFJkpUZp
K/kU33KCxOSWMKbwvEpBvL2sftRiAmcsbkB2lbgysMMmwG41oedx609gCWgT+q5UuZhtQSDJXeV9
q+hfh+nxO3xf6H9NXeS4Llq6ef3N/Wv6bN1lWdXgtipRrQpwggemW6XwXJ/p1DVRpihnko5MUeo6
N85xKAW6lPCC3C6pvUgv9twKkg4MsLAMkwtGpfotSKkTiXcF5H51US/erRF5W6bqiXNVoNqzhack
RJPPCc4DpdikNwMHHpnfgUGhXyOvnxcnMsw1XCye25rnGcaVWBDwCb9J811VtIkNlkdBxkl0ngxP
QfPb4h2yHsTK9Ov5n/62WyC3jEqU3KGe7SmKbkcRjKin9XOenQmtJkSkKs2zt/WQx9q2UTmSCR7f
xea8fB4Y4ziSk4bJdKboWrGsC0vMXfNBg8wxY4z+k6JUiqqbm4xT9RvpjuhqQIc3KmFe+al/zN1y
KyV1H3tTghlWAryjPmHw54BahLEx/sKzgEC/R8k/JakEVTDZkeyArRBvZOL2cA+lpzkYQA3fB/Du
LkmOUJygNNGE1KreYtg6wbg+/sU4aTUmjgAvZ4RmYyv4n2VhIQVq+YmoVni4O2mDbmmRQ2nqZqls
2E7QuyCzo2LT1cmpW4gy/5g3XElTqapLf7i3ZyHd7e21VpmPFN7MOQfOj72pYfepHvF3RDjXDifK
MiJXiivz2ak2c2UTPHURK6fStTciCZYbObMlAT9Ocen8gmwBSjZKeMjqPXxUiDy9U84A0Nigpyoi
S4/T7qX2gNeZEcRjJtK9qpHEJ8tW127EysrFcBHFvKZxouYZ7yG4HXI33OtCtzbxO4t+jQ+QCk7y
IVbXGn1erBA93+sPyPbvUxLCMiq08c0AAwpwxpA3Q0lT6bC9pKuDWTzOfNeNpeu+2SavAtR/gx6X
SdhW8yAzwb0T2Wu1upMbk4TRqZNUd5ummVBN+bNh/FpIsx6C+1unufsneDxmO78X4KLSgdmM5WFG
Sd3sAQegmaDYv8pjKzE/HvSNHvGrjWdcze7NYbOuFdd1VlM0WMOA1joxUDDiLB2AjcKJu0yvhQ4B
5D6YjeJUXHGQzuQ92/PzudFYwZv6H1dHEJxcEzrySvOoWkrPybTfGzRHU2VPxOy3sDxHEvjjvc3K
sxxO0xBKm7TJY0r0SLVAWVa6efaj4NgPh16wfqXxTlnCwvQejFnovydFzekzr/K2TjwHPA9GMUA0
LoYvufnJn35yLoXoM66zZ9qzYvSRKw324ua16+ERpZ6NqJfHQ8OXfTcwNiVF5Wvm48BDzfsnIivs
8/QU5T6lP4v4T9bLUGi2BjXtSkywPxxbqlq6VkiEcVq7GcCh6v9GaaPkD3oJcidZLk49c6fTV0wM
T07oJWOcTkQC5enrsqkL77ek9ry+hkJQn4BP0X2JDSKUgt2Ah7gHH+TqJ6Xu40WGQiy6LYuI1jhe
zqBKyIjmGXJb2h51AqU5TeXittyU/tMQPGxpOeM5Xdh4tXbvZ3PMURs88Q4qKKhEKCytDQ1JS2bE
UxJCU5tby3Vk588tSXY7jix1uJMp0a/pi+/71hyrFIgeqO0bWgNyfbL0IcXDmoiDWVGVRWS5Zkjw
D4kOq8iC4gs/To3AQP7N17quL1Dz2/IwLZXGMMo1xSwuPEN0oqgGRRqOT6RkK/m2JlfooRqh40z2
iuMuaIX46+M88oVNl0PozvuKjxbz4erIu/zsMH6W+Y5DV9F1UqpYPqaZRpLC172puxPPsYWUS4bo
uwThzO0HkX0gup+vFkxaLIg5N0Snnjl5o69M95nFYRAyeHo5iMdZUVbm2Vya0UkWuqbHAPM8XtfO
TjZy/qZj68mHgjWnLGwNbY/TaXDJhzGXIiYXLLH17ay7gz4A5XGRW5iJqNu09FRmmPaNH/tFb8N4
U+MJxbmLd12eLJp7OWhlvuCEqvGv0xE60wbJpr6yUCgz5QLg/NkIARMbBzmPfSeh2JM9VNrGreav
+67oHiJZCQBI+Pt6BdZkk38tT9KsyFM2DR8KajFA7BJXAcbXthXYVZj2RA5y2cb6JUxhxOhoXd7s
PanlJRXyniRyxXYkToAKGezhLOrtUQZnBxG4xgloaBHMRvf/v2zgIYDZsdE7onPYJPO6BwdhIKLQ
EkuG3ICy6RhAKLJh27jL6V4kBphtROG02L5iFDRie6l2+JtEDx1kzFSJ/K902efQurHE7y6Xjw6w
fDNyC4f8ouKpXy8+ltO4g+iW0rtPe4SPdFkJsiQOmt1et2MMs+JzEfN/myU9YBuDEEm5jCmr6t+A
vEtHH1+CVZIDwoJfvUi1QSUfczbleJGL00IyKlUp+nUv0/usSpPgfDilV6jcF3SVmWE5IPo/v4A5
iubJyVAsXv67mO7WlWQD/8EpO21YeAKvFu+hxv4mE3givvpefRITMT3Y76CtAbpe+Cgvnb9JZcEO
BE4wvNhwrFjnDnqhNxbdayPRa8BZqUH9YYbbgAbEH67KS+brZde6NrvnNI5U9xLBXW6qGW3NecNu
gNLXcqEn3X9bGyNIXQPrkzSrzf7XpJgVQdCxEUYE3GeHac02/eoRxtT/3ljGgoLovplWL9N9eA4i
ZHbFcRRRkM5xIPWFJd/UmV6NO6U7q0saE1yah0v6rPyiOI09tHcPMvfUy06q5S4IaihUrMh1wDiM
7qY5U9vczC/KJD/tyhkOAixTCqk2I0HRCoTatCYzgeDl5DvHgIPQedEpP6V8GiOey65tl9omVQkN
cKz2/3UVJVL9TNvX0NIND14iu7dNompv/1b3aKQFq2z/QoEDXKaei7l5lmEyGOZBgla5r5yietVO
A58BVt+bvHp9OdSF4FJ6cK8+SoEc7w8i5zRnbjCQhIMsiuh9Xb7wYJJWAz96lIbEhu6DPoekkSK6
gIrk0cCBYJbFH9WinvxnEPcsi305TYAdOXI+kT2ZoJnLDQmJFZjSpPJm5n9OEKdS0Aovw/ARC+b2
+WkMoCOS3Zp4RSHolGIuwBW4xx3TA4B18sES5UXecC14wm4WxdsL1Te/BdgNcYvtiE+sNatYZF7+
a2hyJKxm9SoY4NgBvDL6VdWSjCDtjMESFmq8Z+DhYfx7/g59atM2sQqdk2ARTBNMz6A+UKGL7DWU
QRX9Rob73RsCWOmcYGpQ7mQw+VYynK6VI09oYcbz69ySXg/1fmusk9y/T5wwffekFn9GaSNTdoWh
QkiFXJpDyPhjoZ+ljFwzHB5WCVCMdw7+4Kn9UL9DQ03ni14zGm9hI/udBPjJEeLOu3sPRDGu3nHb
KTkBkNbn5V2/bGVfn9+ew523qg7V+7adjf7PSDdSjnzEdlv3d9SypGgIWf0GxZpFZyMV91IwW0IP
rJZwP1A8k9H3Gm6Ps7oKi3DdBEuZwQ98NyILKeXLaIQy6Z0kHw4PzemYU33ZrUrxbjpOiYYxXpJQ
Yd0y8Fjyv/9bZ1sEkfj+nJVrq168UNlhSje1CNjlsgI6gSwRtTDq32helxZ5PprMY9WTNN2Ek3Ux
mVtvPbdn2WgvaEuQRiH0T0dT+hw2ERCSFqrz9LfwS7VZLz5UzGaZ51vKYTHvfZzBEMnXbNm7644N
SSLpi4JhRYJ2zPdiBT9dnWyGOTeykF1xTW+HvDDMf3ueqharqbjhQPCX5sOklUj9l2S6ZP6dDnZU
lkorBMk5MzyOLn+JPkC0A31CJ3Pg2dlCqARQCBNmjkc60YhpW1MhFcCple5V3IDqux5sIuzgGju4
JBZ0fYEWS7YPlxx/DLnCjARyeTPGuL5XjCXl5lyF8Tb6zxuHsM3t+qsgQyi9J/7aLYHOZMS/6wbq
SGhlFbcGmE48Zdn0v3oc6LFqR2RuRt303o3m6gcpe9UIBju5QFQLRdcqP/oAgitLIP3MoDBAnQcU
MESezp4bdv4ynbdAlzr/m5mmKbElcWcK8dqJpcqUHKIGLEy8UWizARDwZgMivjWPkPss5AKW7csm
1J+xSpj57HAiM0B3iE+CcrWDzt9L/bCDNc9XS8/E2OarbfSgc0seMeNU8em5udl5W9ncBptDyhKC
tBB6RE7k1p4yCJ82x+xrFaa+qVnXwyUxVuEWKiDuDEZCMuXEzcPGG0tvH/89rKxtNfxEWJEmpShN
WAuOAp80Jf6kBiVXcgZikVUEqZ7AC3mMf1KWm2TDWMPXKJRgScutxDFBciNMM1UII3Zk6gdlxtGm
bdlb/pCyXgijGb6NcDDje24mEOP4miawuxOMFfeoFzRnwipghW2AX3QehiqzUmavkcRDUZ6ocvYc
IHyDfzdVSb1EWOJoc4y54YhSL1t3gWA6yqPVF2fLYapX9lUEigAWHQkjcSaD1StJUlAWYrtlfgG6
CpVE8SZDWFZhagZrSHgN7HrK+CbUSNEOBAWvL5Lcn1OptrUus4lu6WB4n4wMVJPgNs0pw/L2/cVn
BPWAvJbRcMj5Md+iJLwKKzq2iQWPHzVu074QI3oYgp59Bkr6iOJNxxeACvnSPX6GgDw9YUO2Xgga
jX70aoE4wI6fRMwceC4IZlZ+qXhlMgZMxUQhgI2iQaL72NJZ2AaJq9ZU2a3X6E6G0idfjhLw9ylo
qv3Re+EpkAON4Tbga7cHnhn1Zs2uvoglJXX/JHQxvF7uiN/rfy6hhe53YeAf+4CtyZR/LP/kaZjm
DyRprxB4CG7vScRU7x3qYacmG7CtAd/nkHl2InVG8fXYoOcp1FnzBT0MCqB2pPbtkckSsucsGV6m
luko24v4bby3SQOm+wVToF4qlsQzaditrG8Ihnw0T47UiIvmhArDSg9tfDfa42O+A7gw+/dHB6jj
OBKMpVNaEj85alWl+glReb5SNSlRD3bFMsF1QpHv66IjYdS+321MzNt1KpsSYRlbUzlv7b/6bD1w
4ooOynzjPK8hyXFucs899NprU8HIboi05jgfFBBaEhUjoQljMGQWR+inGCkFHQOlHXLCpqnG/Zhc
/OZ8XjjG9uODvdJ2dR32JORqfShc0RQoPghKDUbUB7VPYznwkv93BOZ92wnNojfliShfRq47PiKW
2j6COzCaxY8C+TL7jUKOYkmXPcw2BfanmRhUnffq5Mcx2m7sSRRNAvOtU0Ap1Dl5ChgnXRo4Qovf
yyQuU5dWqgWpGixRcQUe354Xr3q2PXOldpSCvQKKQBW6AlqF4ZTaoQGP782ARG3QLNn35tFYWn7O
PV9W7t2BAsGkehPRJ8+9/HjVrrIOH7Xdp1ImK9+ltWVcpM6v0YK1PY6T3v1iXaO4OcUTHAaaJWNi
76K3qSReuaHe/zYoF6ChCdfkFfANA6Nk/4Qy4UFgQIsqJBQyaUDbQYK14fAdfljSykJ6S4FsY5KB
8Fvv5rMv5YaSdhlzdLEuwMBP0cIf81Z4bA214dKhkcnC45scSfYM0WaCgb947wrqUDBwv0plgeUl
8Rr7LwyJBkgk1ZtQRd38qR9KngrIQF6jcQNyay1/JMmqjxl6LNstY/+l7+XeqM1sfaRx139BANeH
XaZrsBbHuj8abCU9b7+GcduPY4AfsNyRG/1G/m3fNOoZGFmW3ebVnNFyIvBN2OP7i5WMlG7DhAe6
nYj9uEPNuM3DppIHgIqFOXhuRZQ68dG++ZXqgsnJMChL6Omgb+MDQGTnCFxwdy9waV+JzNVELQbO
LFGSSW+wGje3ndvMZRkfGTDGLJ+v0YUB28b+kUfcKYVEP3/dj8MTK466WtqZKoeZuIx/B/x62C0Y
8cUKWLOd6Hg1UEk8o7HWPJr/xGp2aSfYfSTyqmzxdHld2byq7XNalL4/XbNFfhCWuTH5GzhnJGQG
BpruuRxh42mUHUX3k27DH6nvTCMW2wG3hZKS38VMdXohVWk+RQHgr1hDGnS/pDc1/frylfET7abk
ZtvR5+grBcNT6bXmh3a9FnZXqs18rsqMRPec3OmJdzp9Rp0HoTt3n8nGgLS3qRJyp7K5sZY49DqP
JTjErWDRjPg2PZlWrGt2/nWVqy0Qb5ktrEEuTCZZWfDGJTeX18JL8arkJT9MwuEc2MSiDaTHpc84
iNYjmqXW+K3FOMl4M/0esRY/i2XgYvyM2dqU6vC25BblWdNS0vuyZXJOsqcxt/DWXBkNjRwtmM2N
SxuRSu0Dris6z9mNrpHS/dxIRcXw5pbc4w+fcTSEQGrS2tuM4HbXDC5ht+5YXSuVXgpym+EmMhU4
/fnc7fWJlNBiqvpLyqDr2jPcBzFYiYhq50JMG43ZLsPEdaWAX9JgMR/7GCVuCMLVVtIMa8FT/i+F
aCv50ne1qaQcuqm3CmNbgnx3aujQHfMAlyzs+1y6JfhtCfyrpEs4w4z+lLo8QHmaWnRVpVtgat7S
koJBTzXOKByVLF2Ld1P7YHxnLg0WX69XVu7UEoYZdjBzTiCnwWV73VbipDclLXeV+fti9SgbHYAY
K2hTjuSZ1aaUFZGp00hVjtBp0Keq1rQd7Z0Ptb0AalIF3+JhKw3uYecJfqrW2cq+QCRAXKvIq1j1
4CeYr4PKLi23GKPNuMsJtjWrtcS/vMOjCHInZDIvh3hFa6qKs38W48EbJLtDqJ0B4vt/Qu/k8vu3
iNaP2JL9FhYFb2KB00hzuut0UuHvxof6IW8l6JtHaOSOIl09h7B/zLYW+7nu6bx5xaoBaWmVqT4w
YFrsZTeCuKdxL8AKnYE4ve4/r3VgnutDKv16HI19pnJYOaau18G8ZjojVWl/VGrR/R0FSeWQNE16
Vp6ncXgkJwdEbarJIC8uM9AfpLYVhREoG26ofG1vt0AOBF6FGBYcGGvGUUAFp9n18WuL/K0yg8xZ
edpJ7YridQ1QaWdowbeBrDMU7ULhWQkgOuHzOOhScOUL0cxazEGsQuOMQn6u8znLEqxi9zUtuiAX
aWWd0W93peWZGVRUdzOaGcb1zXurpdiI2srKi/Z2DCV5mo5e3bnJ7FC9Mj3lc+bDpzpuwFMY11k1
0Y8EsNqfYpJchHniVd8Xg8LygQpUaM/lq7FVwAD5xCeaoQAwCuhZu4TcV91pyAbSrMxfcOrh6x3w
nLRqwrMw+OdbeKrYGxY2/XiowLDNHIt7hBnQQI2cqJpkKbL4c4mDGCn29vquyOvdiaGO0wMytcDQ
syXUk/b9d3qix7R7zAuwzHQResRVhis5ecFvAg1n9+ISvNEZyS8KcmfgSs5//KItK4RvqBDzVkr1
ukNejzYxGtdej/5DHfD/qOEbZ0Mtpg4wmaekdxbpLqNhZIc/PnUKT7Aot7rxhQy0EyLc8gjdIKqS
squswI8cbcLux8dGN2t4jADQcqYA2bXf8uG8mvVxA9bl0dfh8zUgaURHexS2Cjx3sNYb1Pz6cc3P
+tZuzH6vFW9j0r0Z+oH67Z/zaAMBSTyKxiapvSBKOGGwZUXhlRf+pUovrQqJNf4z8zwPU4z4Gybb
poc7O0DFWDU0T0W8uuZPnue+JPTjh7SauUeygyas5oZYj9+MYoO5+oKxgjto37veY74q/ewEUCba
j9zi50G5r7jfDIbmEYv52PJGN4kmVLSqnbkN2VlA686OBedHFK46+e+npi7WqoWKHBQAUcNOUVTV
EyWYPPexxpMoSIRWop1ojudUc1h5k5aDOob8h7AEQR53mG1hQlxGgtvrfmsBY9F5Tjvbh7K85T1K
hpD+zoxCMm+35ryfUux4Afn0wTQOSaq+FHN1wHL3mkl8fEHgkifNhj2XpIBgbt7g27d4HE28bsXB
dzKzXvz/IhSYpqKE8/Q4eNvvrZo8rEbaHGflp/++ET4UAxdSDxigVeouT4+bfBr5rIuY/zyiV5cE
XE3TUh5XoE4VR1UTGxyDMi+fEAqtqt1/WGNCKPAkdbtAfNHy5UoopN48aQ7X6skyclldabRD3mU8
7MCK/k0Br9Y05KRQmaIzNvA2nhHqx6y3TEfQkiTEuCYt3+cJKwtq8oOQ3AbmmoxBxfhZzrbbphNw
rq2d0qUf5KujXmqS/ZAPEf2qrxz68/A2WlLMt7rSPwY3Rn0leIYO0nWAIeyHOLr/6P0Uim0OOqJF
pr1AllbrwwqzcYgilc38xcA/ssiDVssFdFWLcW5RYMk4Yf09D1kyLIhIHdTYQhpfchK62zyf3Pt0
hTXSvCoq8i1drWh3vyqbDgWpVkbYL96HiJUG/ftYrEeUFXSBH+DATT7mYe22JXduJqxF9yy4eY46
aoaVJqM2amg9gfLjq2HzbHtXk2qq/3b+2GqQ/HPKMuLZqGz4/YTre6s0YmRDStvtdihtxvra73Ug
+5GPWsSYpMDoy8MP/m+nVEsm/UGKJAKrYVnzsXmXbqJXDBBZdp9wc/lQQ8rndMlEo75xyujrx/Mo
izccF4l5x+Jos3tr2oltQ39BluCvg4eEazJQq1E2sCbw1Iw+4W7Tw2mlEaFu/tGQ8dKEd27wNWK6
YIKUf56KbolkneMPK/Uf3eOAFQLhbEoITDOWcdCDPd2eMN4F+F+2/958WA6ZUXW7yKoSx1BFIhAF
cDA1lp0R6VPANilIJkKcI2ZV797MBdELBi9BFotDk9sAh0oPWGAZJCmcHtnELgB8pwMNhwHUY/zP
5OqtmHMjVGkgU3vr2h7RWsgBYD0vVHUpCCMQ2uAP8jxveVNsKb23EiuvTFGlFmHPr7AG/EvY5wvs
fITIjik0MmIZKBT12B6Q8L/nVaOuo1UCPV6isO8k9TiIEBGVAnOY6ab9iy8OCJr9X1xkdjXT2C0Z
Xz7x/2FSbGevX9of5xMgoa5/KCDGF4jEsYbfrRfxZeVO/3w0FJanIT2PN/pZuu+GGymIpJUMeCEs
AZwLufR2eaWRsWUr3IEoTjZulvgDKpE3JU/I2NpDo5XHE12HybvVrc1zHtzun3T0XMI1EET0SULX
8zQ+euTfXxKbdLVhpeyaRM7fQoSZ/VzdS8NP1y3kP86fGVjx5bRpp7c8q458IfQ+Wrij3+49NVEq
PiKVXUvoBFebDj6T1fqTyw1pySa2DhclM3pTbOJmpm9pAVXYKFP5Y/FBC5rAB5lw/Nu7z6nHxvjV
TNo8JQ38TkZvjPLaa4VUA8SO4F3hxW9TtW5ZoVliR5mund2OWS/QLGGHqF7CHruAVY2r0gRnL8//
oEo1oOX7eeB0zH3UgAm5iP/m9mhiGoXkIGOcf1UP+0OKUXbLtpRh2mr5G0IzS/FyiBejLanNr9ks
Xegp6gq9EpB2OK4rSjdwpwnK/zFO88X5m7M+aLrsRIAgNld/Gy/RedK2xHpJCMiDhnnPblbC0zBh
Y4MxNr74HyulUhAqi0CZXAW22Af9pRghcA34peI8PRYB7JHn4if51v78MssoFR6Cwd0mAKmx/5hP
Io18m4OnckjWpTLJUrVVLYUm4C6QT7zzUP4GgMTxVDqcOI7S0HkZtCjXpOUO3mB++U/8/dwXughB
4MgZZXEitnpZWkBeOBN3IwLJFZs+9E/QsjgQkyYp8Y9nvWaRZKQyQKapvbDl6YCwG/Ps4Kv6QMCt
bIo+2JfNYM/EK97Q6HzSED+DBcAVJjA93gPUSohnGYfMMKwWsjj1YToD4twjwdBLHALX04YSFd4P
d1xgeiZYbQ1a3UoN+4Mu5yE0A1GJmWLui4WusMJR9b7ae6WKAT1yDP6jYGVag27j2BHrZCYGBt2i
dO/afrbVge7fixY/MQWVhzd5/nblC1y0ANcr8ucGwJtYYnVvkTSWRUWKsOFrWrQOPFSws+o9aLwr
0PejprfillgMETcwnzPO+dKZzRPH5w+5Fy9GWAM8FZST5qm3jPrhj0vH3MTXhPG62nlY06xnOOVV
2S5FQwIHtT8t0AM5bmod1HFLPlB+sshAYZK3eyuoflxeKt29TBSEuxAiMuXPLzsCP1R+GEtP3D7J
KuT92noFWPI8fPdL3D121g9iZZxnvn7nH0zCj/CnVtvmDUqdVAZxK5ZD6fTw/zszquRg+yQQhmWl
awDKbYd+6kMnYryiBZLo4gIw8kSygRSTqL30/079yNYBdM6zlXYSL9I194MII8CNGLdC7o9znYdy
jlzHEkjW2K3RLG7ubyWYQNfjKoZ/roUTDIVMaXUbGX6W6eaYfRfdGdhBov55T029Z8NihCzn58Eb
ZN3U6NtiHJR1XhomAxVIB7WnBqvXyhJr1M9zdqdHoGOGp3Nt9M0gScBovTDqmXnoBoCF8EuZebwT
WUW1/+rgIx1S5lZW6s7GcFYq6fbIxkWQ81B8y96JJ3u5vi+HcFIxdUDiuv8QrtYxWysIsYOnI9a4
0X3CTu0WrnucnyRPJLlWUUixofoAKSPMQsHj6NhzMSHiStVCA7TVfVsByy0SU3mJtgR7TblDsp8W
ScRUcZu67jJHvWXGIhbFl6Ti3xs3t6IWOiVF1DxHCJzLBJ1tocTmLFG/EpPgJ0knZWDaESkhoBrK
8uJe87hbWze05VYoVXz+RfgXcx7KNHGStR+/D59EIG2fMzz3ozVqHGV0+aKmLzBCEM/L15iGVvh+
kA4EFxvo538idU90idLCNVcPmRnXEWnB/c6dErL057AEC4hJZeGGb0tofb6dEl3JLOd6OfVbYa55
0AWEXXQieru0yDfwquUaCiq8UGUEEx4JmdGYgbd82U7mX/3lp2cCO8D0HyA3Ob9GA2PUpQGDox8e
vJiPNkMOZ0FqB4ZMe3XDHfT87AqfAOoHpyiSgi5fBk7LKCsMG5Gr/IfcKb75W95bBNbgLxcFR47f
EGzlWV5CgqG7noc6pxFOC8Z3iEIKeoPq5x2mwtktvoFbEsEWQ1Y06V8vFr+TcglR+TogCYS1wwZM
ZyHatRe/+hfi3ktn8GR/KBmZmpBbH+HlWoCZS9OBkKEr+amKLQc+9JJBZbaZn7u0wVoChhRDOAAj
f1jvI6Roq7cAROqhPCdEYR71067VG0YZOXnz/w4cjoCufeExPFaOYFd/LAH//at3xjiamoFXqRZS
Xlq0Fu1ehOeo0rdhP3XfobKTAZ2GSPYwmt1q2y2VGJCHIW4ge/bV2LJDjh55PBjuqlStaleZm7HE
qmpLLrZa5p+gJ3wIpAV1nU6iQrZjkiEI2PKTHqEXWBrV9B44ERTyScaqEqUBqXWQbS5YVdX9aYeD
UnQtZSNNn7p9TFFTuUsk2c2OPG7b0tcRZAXr2T5VvfEZSKLIfBCqKIqskeZZ/vkIJPOEQ89bnI+R
rx/fJzgVMCJhdArDLkuuLahnPxYNM+mdxUne1876+dvPAsShD+/Q86vkunHe8IqtHfGFHOcLZj9m
KzM8RsAnCLBwKhLIqHV6OStA+sFm6QVnbxvMNST06jTOC/eZ9I2OYdxVi4Pa1nvwoEtUBnQp3So1
tcuyjk2rdKQXVPiI1Cp76LiiHxODGTELFU7ove+Qp4gHfCSLkEG4oumlVQ9qs/m0rp6Rouc5MUZa
a530zTV2q4ZACnFeudkvYFWTd8fvJMDgnRwYWhriGD72CAHtEr42wNgDG1mGZIxujD2n6mUjib3H
Rh+Nx/HGoXw9jMQB3J3nqKBanKl7UAniNZWUnzJrRrzLEvzwfG09/usKkG5VqlnNhQDn3jyIlux2
qwYjtUP8GzwGI+4bYMPiNRdBvCKUmcHDoYTNNqhpAjZ2BnEDsuvewV4UaKWDfsUsB+1PM4nif/qj
MXGIy2sFerrnWtIt+AAy5K0BdGUxwz+TUIKapRUZ+F37oM7B/1BHA5Au8LPDZyVmedAbd4ooWINu
UR7LwOayeEtK6GFYFpR3/YYEHdxu3xZZPga1U8WI9KbOXJPIeZAB+JLv5SJM7lwfNHaDXQfGtrkV
g9JTNXKBrQnotiDw8UV6G77JpqvKYFwxgDElhmL8tuuBqMjfDG3r7OJUBK/piRwnQE5JWzZVNJeb
uMG3JwY4cj+k1Wo8+pfcdWbsd5CRfGGM3Vk03eY2az4zlGL+Ak6EOJiC0o6sw/il349rXOkSF1Sl
d/VlzSoFzurmnw8EnYPOJREu7x2TZWlNm9TuoJS7cAKSPRZ7P8r3OwUHSwS83LmrJDA20i9Kshn/
32SHAvNatyz3dRm3o1RD/ENlVYAsDz4MYX2VWzYMNEmrGcU94yUu4h0idkUaNzbHU3bgpcKPYwoy
1SomnymBZKpE35GN/+VZnxf6X+frf+fiAwWf5iXXy9EjZjkx/46RMjGi6feq3Go2PMcEStasGpJg
0uJdASRFzAVcE3zsR50/HbFPJ+cPOEwG8S+PD3ByWgf/akAurRoY+Lwi0C2NuIgO2e+X4WHpjMlK
zir4Q7Dos/w9hwghRsPHjEimEOeU9r20FTUNrliF85idknmcaP+YvUi2ISU9k52bMr/PLE5iElGt
x+F9p2+5Vrd7r+zKyWc7v1m++h3o+P9rR8NIUARGxT2ypfv9pIu/5VoVZE3RW5FOe7Llvq53ewcl
GjL1gIZO4FH69bdO2QoaGIWR7YrjauJIxlna5VNJAohpjboyOKwG7iE9iPV0EIeFrbVq1+vEUBXY
UYMKQG+VOzy9GVMEui1/9PjPRNaxlYArGCvR8bJAQtU4umEDK94bydFDxozbJOqrZpuMoe2HMRpq
hwIprG2a1QCp58oNqYgjQbE687r/7Ado76M/EbZRBNt5fCeAijANZRjpp6HCX2X0OmPDywQOO3zT
ASyaahadep2JmAh6XMyD2Meq85c78pSX3oWbZ+rKY6zX/kXFWRbWYf5LH2HpkJZlbF7U9wbXIFeL
faWbAAcMWTRs/U/xJ7oeAIcQp1eRAIbEv14SUI652A2ZsxPrTG+1nksp0MtTOtwR/anRaRApwxgX
v9nQJOpkfTmQBwfD5Ca6SvnxzV9yPoJsLY0L/BdQet2zzKQfuiORFSZ+0AoXAjtPNTVk2BajdwkM
j65Yr6h3V4CowLmeVK8d5F6+izY5zhfX7X1jWK3mSgFJCZx9KJzqDTGbgiyFp5qYHKgWvRJ20sDN
U6ABBDyS3sladIacuqNwHdNuC1p4yRvkUmqNeydh97gQZvSTVnfeBnAKTE5O5Wcd1fDWUx6IRzFL
WgBvhbqU8hTbe2AUy4796BUYha/5J2IszrNsYB1P9dE1RHkLMclsXPNQCbi3HwhtsficIP7QNIHT
8sUEf1sQq/LuW6mpEmJa0bwFhl9qXOMoy0HNtbgJ6T/41Nzxe/9Yqd7SrbVkritvg/U0ZkXIPY3z
EemxHJnXs+7mb1sMi3LaewjAE5UvC4VSgzkW7KXrpSNbRjJIrDJDXByVVD9p2HSpOpzmViOVPxER
BCgDqeSpXuCJJC18BmXQ3bFzbBKFwKb3IpGcpXzHd3fEyw4uxkzxvL1MffPh4XFUemTenre/KOOb
F1+jzECMS6guslmrm+1sX7JsD7HD3asaU4lYofSiU8BM482/G1Z/lLzBFbz6ksbuUZ/u711h7BNC
KlU7Vvhux6iDzlV0wvQPjM8WmNHD+jZkN4AGtX0fPBhcHpoQL65kDB7sv+krlOvWs6q0OUjrAI4Z
lmDVXC0TzsIS9kMawp8+1Gsn3/SAuXn739hcBDNEE8NhBFXa2Z4E3GjH3EEWMWoRhMQ4xh2sjSlo
tZ/kTTJ9GEmS7as7ekTVN8mOYSL4TNo7veO/9mnEHD+8UDPT9RUepC5NZJHifATuk4zAqqh4otmW
WkPsQ1FNKlwIHDw7Z6D2i3RL1eRiepWmcbAnaY8ZlufhqmfzqnPkvVRKbwhxkCWOLqe91NULKyIl
HEyPXAXWBhM+mXdpTq1tczRnJz4D/AXCnRafVGVs0QaB/HZwNfhy1jK0PTA9biy25Di2vMMmwfyR
HkeOmW1JQbBxZv5yL+Qeu6COEUOl9TORGSVw6pR8v+6vIZ/tSdLw8f7ZHlVMN5ps+SDwrZLdmfZ8
a4GHN+Et0L6U38kRoLqqTTgIgeY/+8CSt1YDW/T3ENMeMpEBz7dO6tbJm/H/kYjthgbCO1ZFay3G
x/2/Cev5nW3wOUvNqIoS6/UuAaD8orT3ux1VU6bWRT6dDlGULfbugf3XeRj4MNsXIgBkWArmwd8Y
vkQU9DuY77ZZQd9EQUp1GqlK0wfTe9lWBvGnktFlTx+x/cBgN+XKh9YhKHR7ovQtxDp/CHBdcacK
al0tv3NmtFqcrtbkzoxA5oWAklgVN9UQRhHanHH9Orlp6fcmjF7ftW17O7QBou9kRvB1LfhWUa85
wpo1sPcqv7/CWc12S2QbGpN9u65BhDOD86hLffdLXgbCsoHahIrA7Itlwc8Es4+ke4wzekAZi/JV
hBI0PSyPCt8t3KVzrqAKiLcM27q9YzZL5ulYbRnilAmyLgqdVqSvNsWMo39i2MPh/ZNRML05s5tV
XEEqxxVQJneJQnY69CiOXvOYJnTHI32urt6MPFj8hdaseM4PP3Wm99kI99i1UH+uh54k8QVDsvr/
WouEuVyH4lETiDztBOUzLh2ce8UwrefLavo6Swb1DhIAuN4srXmeQAT5xvz3CR9x18aRe6VvFuTl
yP/a1Ewdx3CtpicAUOPFFxVV/VNreWZs4IaT82Gh+qvRDZYcNpFMAoBhNjXEGBFiRpjby0ixzV/6
Dks8j+vYif3ep+rUtYCvjB0SZeLKObG6czpqjJNJhxMPQM/CvrD+vw6AMlzLQ5gUGqkEJQ/sEkSS
t2lNUavPBiHWF3MbrVnUd4+zT2EQitH1bX+GA3LpS+3agHL92hQwbT9+IZEB1uZUzUDH8Pgj5P3x
HBxjcrF3D3fsKIx7/KoLc8KNOH2Qww2U2XIwvWWPg7d+AFNDH6HFVMnKcT9uy/PuDSpYdeVjm7MQ
s7E+X/CcW19QMrihblVG2o1hjlv0JCJ3SDr36YRV8LkarPAHGqJqOP5uFkp9tZmbZzACq+igDZ1D
2dZYSmianPqLuSNMuZJM7Gze26BaztTNl4a19cSrPt0+11yvci4ZyZ7ronRbMACeJOaEXgMzIdrs
30dkxBEQ2VGyvXhChGADIMA09e2dsNORUEUd+zuFyrslH0sp1kB/dcy7xtle4lX5Z4rdmWB9vT16
dyRb77U01oErsRbZZ0iR2/TdDK3BHFCu7fI91mmp+m3NyvJd7wXyFnHnaHj5i/RhirqoV6Hs93Ae
ci1mA3WkG6qUBaFMe1aE3DMY9zKJzw8w++CISud4spPk08HWEqVTPm2UdQNBjbSg+LmvyUDIAFgm
hEY+7ttbDTH9nISXnlHfl0x/BdmOMZSC+xHOMRljPVV9kCYHoCAzgH+WWC8HkctoXbz+5u1WE0y/
dvnfjY/H7ZGHMzszE3HQE3rwuG4EcZxb5jcKxNwspG1n3hPEWlGimqVBwnL88+T9g47DIWGAtvvP
kfqtj/LesVYLgpB5GMGillqAF0G4sJW5Wj0Z049l7d9eVc3t4p498ZQrQjFX+KO/9dL14KdeJLXu
kcw4BxJXnBryIcwxPTiM5brajmuH+YFTirZYdaKco8lkZVCKjbWIkYtRFdRSRkqxRBEaEscWvmEi
ovgKsbYIRKcEJYmaD76Eg4rbcocVIsOcGVgxhwI7wYULLZJTJ2gvUspQtkfmCUh99rZAogeFC9e7
gt3l3ly+7CVjANWRKsFevvWomny+uH+W3Wh7zC+3srW9xwTbwXkh9iSWctW40JYlZ/nC10ARO2la
zPLvolboQUBpgOdHDRRVVVvnuFWhkjACOZa7Qf6V504SKpXa5e++lws4aWWYWYbEXAgOlqQI24am
7/e4DGoMJxnciqeuV1oW4M8itBafOVXkKghOYoAcYAqd+DzT7xMvsPrPBmdjYEKNfwdxCZdgKUg3
rrg4FkH8AmDZBxLcco7hz1WUA8FuBSbCOaMBWsY627hdADGMLiMw5wGOelsx6bbdowkopqWLU1+0
yLC8KyYz9WjTxWjE7pV3JsauybVTy1FvlU6hpiJfMyzJfuDpV75hDFtRoehQA+YNNy1O00DF7b9E
j2UtUwDEj8Yt9YdIL1R+8ldjSWt0RtxSe5iGybeyUIuNx8sYm7m8zNOUq5ne9tl7huRHpkT3UpEB
102kYruBXcaDqQbLUoMceqqd97zjy3IGNyXD7J3Z7JxFsAY7YGWo+iGzy/tj8QncsxMsJg2l0KD6
t1DlGTQR5ncTWVnjPS0gKBHt8xp9gBMlQe0txKSRDSjam/lB4bgNC8a8WagNuMQFKiDMi4PfVjJT
j6Nqrlkg7F/vpsFQqPWYchswHkuW/qINLrF5RPlyLF+kTfBvDbtEoHdr5Uz3JmCOcCZ29qKHvsnA
rENBHfBoOeNfq58n09rIajeR0yzhr3mZKWHa6BDIoR0UBOs6D+4CSs7RPwwByrU+w7T5viYXTong
kH9Cs+FEoWKq9PFGVUJ5Q5bywHQZi1tK7ifTO5kEDmTYaqesUwbJUG+XShKwFjUSM1Q8pwliB7Rg
RqFA3vcHapFB+joJ7271i5OMN6I6uxopdnNiynVjJ6nsw3FRXw/riXAs8661X3i/5yA4KGPjEuFa
0xe2susJDub4t3DvCS5TXgUIyBCbtVYog/v0jnfnNEz3ZP//VipRICy/g0RYi77tfxYZedUOPSqb
qy9MpEdTJPNr66uofSSAgpMTKTBAssYdryuqgVwuENlYweFAQuElpahTUiprEjUjrYY4dVG0M/mx
wFANqRKuRA9IxWh2/b38pqwJJMYC7yu8tMo0WWzw+VTEysC8CX40t1riS757eYsbg4cx0qG4SGm/
39TKk9oJVnN9X/vsDf3VRlUSsjCLn8ptTrBAyk6nQej8tegPtiLijp0CIxQW0awUwfPvdA5yIQg0
s4dTWi5NvDK/ip0e/M/hRIKcswlkOQ/8KYaqlB7d0d7/MPmg4r/zN47Hdy6fZlP7XH5MvbZKBywn
G7jysQE3eCoEA23vsbL/7xwBXOKaAvYVLU5oi7uR7dtAVWO+rXYn2LvsY0hq9TFtheHeOU6SPl+z
kEONpzQS8YCSlcX81iUExYvaPmOx4NTrmD+n3Zx9s/K6ZDlM/sZwqU2V2LVDkbaW2uYkyGorEr6I
bV+bL36NemK7IQNWOo+Qx5+vUo5SdvpCuusPl1LAYqQsYljh62Awuhepe4wNh+cgWCfocJE5pqyq
yB0zfchpdsr5MSisdcyyrFqMUdPpoN+FJXdhGQFzOlIA2dsAhaQ/ehDNgxKIQKRZva595N9sEmwD
gyqL+2fVQKIPDTqKHeHUUPEMeCZA6LdRCs9SWDWxNXTlMKiTZ8IbDtJ3CIlynfkNpdSdVUIshRfn
mfSz+xVcv+MUeCil/miMdq4cJRL6xu59e+74kIPqxkh90bdB3mCZa1SnJ6dlyYS2US77NYv8gxe1
lTdHSTa9K6yK033gcqBuYHRlkMqT9MZRO2g0cDm9wSu5mASGfE/MmX4MB34DWV1ZHxP9MIxf6Qmu
+sHjeyQBMNv+2a7xggH8V5KT58GQAsnJLUFCzoM7atZ3+cTtotdVI1hGf+/EFzH2fVZLtRe723wo
NrcbzrQUBsdkAdNdZ0QnuLbQ+YO3l1N14UUT0eHmB1md5AzfTxTrAPD9/S6cbjK6M369BIl73hHp
8ZBrcCJKiYKFPqrNlFiPMiGw/cHENH85/vsceyperT2F40VXV784dLPE65D/BeYtYwOzDEASm8z/
Aet56voU5ldR1S2B335zya+oDMHxCGzIW4IzZTCdt+CUdpp6mplMMro79nBbRm0F1tcJyuQTh0MG
Y0CTCJZx9d/2K/Npklw5L0y0A1iRubmrbYoWn6ZeXWvIjAKHYNBK5lqwFNBIHLCUItkVFeTI6X7T
OKs+E8hYOrSEefVzAy/lUMrqKieqL77EM2mD+v0NTL7mVhiQwUKz7cTSKFx2A7EanjH+vNabtPay
XoL+eTnnZFVoGbYg5e9BI8TQtxoWpYzxaY7CaC5E/rGvFEZ9RWQz0hsObgzGOQgVhSJE0yN1GQgx
PCYh75OmF0SRMKOyVWLmBcotXB6tTVxwhmkhyR12SUC7613NBuJI7AJTgISJaq6B6RAs7wCs+tI2
bJjp7ioDXRnaJxC7h1QeZ1chnR8z62+rsuGMWpf2S/8t56eRVnQIiEXI2W6756tZhwmIG2bKi8MZ
NbjnnNk1BFDgfS4ZFeJeHkpHRiZSXGTBZfMfa9iFkyF+xV0KEwLwA8xT+C7USUgjIKvL2NI/BuIA
g+SVKP4bSFCDaN7E7Ek6iGF0cO9AQdj8UlP0KYKb7HgNJwm6LNPeUyIHg63xXFK53xp5Gg5aZ4aS
1cHEvkgC+couRSVlM/ICp9b/yhQifSKXhAGZh5de2FM5uGUOzbMpBDmDpe5pVAKYjCy7mpiBxkJi
GuUEU4Ox3B2M3DSjpIBWPgw4jbJ30MTxgHKtbHZNh7vOaoTy4n6N+iJUdmHVAhrSwv00HSoNZdPj
p4YsJjFbiX8+1cJoPO+Z9Wn7ouBvoT1ehsCcRcNG8iLqXj20CYqcps0a3OnAPWq+ylAgGX3ztaHr
NSvts83kplIZ2sypG7Ds1hHbMuJImZdxnhasVI868HwkMOBKI6iZJhspcJQ+fkifcPVHYBFu1Qt0
4kcIGF4nr9JgiAElA1CYOqEjQCuakzV9hQZ3ImAv4jkZT2n5O6RopOeWaAN3muuQawS6jV4KA/Z9
MpCD2w0RALLwpgW8MtZaJX39ZgMntO68dfw+QpjuiPgxLoNWx87K9sjw9e0pWriG50WM6/bIOYqI
SD0HVHwQQwpujtvyJAxw4VOwSgl1/ZdXjodnDSugVGRIL3dYM/pGfYBxhKNdmzHH6ayhLgkolUTv
nlQFl13IX0QlrEyB5wnMFXWkPDzISiaNpNvUfHb8+DqjPrFxRkjXa1l2n2sf9jEnqGBSuDLUqhxs
rWIOAny4BpBjHU+DDZsdSffaNDivstx9RCw8JreW8NngIehCqMXuVicNZhvtZvyuygUk5FZU4adx
A6P+9qWqYD8IZmQbKFbrMjh1gAhg/3bnBBtthmDNZB5wlGbDv6gVPpu52djiCUh3nAJYjedI8/SC
W7CCj81dWre6sIK+aMmqIi0/iae+UbPDuS9P3NOXIx/uabT5BMdJRzwmxo9KV33sArEfoQLZDz/t
dldoAQIXuhBFS7hlFVLykk1N75B0H5u3VT6ve0ZXFpNx0vRyPa4UJAzVYY9H9n3PpIBYv4saRYvB
TyEaDOU4A1v5sXYWrRwHgDDnXLDjgd9u+nLm4rgoqHhSg46ZeU334wnQVaTIERXLqzAXzHsN2yQY
gFEnayW1Z4DfDjZLeFk2uPazHsiXBOBkpOL3iKvegqBlt6GdXOrLRbHkecn3kxAVGD6k/Axpto0l
dN9neElha8kTylZ0udAExmemSpSWh03RhzUgKb2tFF6yFYD2PgaemJViC4WO+vSq1kmjWz28ZFVj
x6sPJUhU/K+Jmtq1/HMwciOIqwPXM7zmhX2PX6IMzGnCCcADp9lMvCfnvJ+5wnxjwUXsNlvC+yH2
t+LDKd3H3iM8yTW3Tq6Obz6WMCu2RnHI/mOln4uy1bjs4O0Wyl8FvibI73QMzhdqN5SY5Bfn+uu+
I4AN3KVxpHYPiM3/Dpei0k3x7uy/Dsy6bPf7HrhMlMb1tNt13NCzILex85yBFQSSWIvgo9mnZ/OW
2kZacY9X1aEQKlA4hbUB6kwXAgEFElf75Mi5c+G6D8s8oYcE0T2fKfJTG2mKl8cUBDwbDkyrhb78
b6iU1OjeXDccVY1Ycjgt528jEUuisYyRzudro+N/K36pypYDAXHBzqtjE17sxhsbOP80u9nZIrID
o90Afud8x+3gjsmus1yFsYgWxGo8DFUVTCxH3CU45s4LdejV8M0PLsAGQP4wGxBJ4ue7alxR7MH2
0x1xp17dVRIB6pDgnlx1DJkVHqryPrc0BZGc6tqS4TxbNJVucbuE+x3NWsy2OszYDrc8hYGRLLni
+4dUEHszRrG2oKID21WssKREs/1IDSa993VRrwdfY91MuZ4KB9bRYhz4rlIyEoIyEJLJC9xin5J9
BcawSKmHLRAGW90/eZybI2rCuLjO/oUdY4/YqQ4N1My2cLCAsomdTMVaSvhnAuT+Y0m4si5XI7pL
NcIAQ3UVNpgyoALN+dsfd0cvJ9V3qKvUEdiCrozpE9uD3Y1RVg+2ReFEXlIte7CWZejCYmI/pd0Z
oBr0D5SLvvjcKNoYoJPjtEXlUuylXGORE0fxeA7pypqwXI+E3bYNZnEH4D65GwTtxig2XE7/OL7s
uqPHWyl5Z2LLvyga9m9FN2YjamT8QzZGbKebGLRFOUf4bl4upfRoOk5ENbNVdjUA+tNSKJj+cLj1
TQMv40M0IqYc1fLH1WTz9y+mIKQl54psdFXs7139/mMaF9UQWAuR57/sdrcbjHg5/AhlOJsw5i5Y
TJbUXDs6vSXTlhLDe0C2+TA/XkLHpQGqTwtv8YVemft4rYOnmorTm2NElijLdx6HCRVx2/cZeoO/
Aq4IArGSdt8RIKBFNa1hRCVGQEK/0lrM3oW24/F2IOdBkq/PpNLBF4cM2mTzAcNe+1KjGFXTe+C4
rVY1Z6agUZnGlDoNsidUR9Hh6Gg1dPeT3xGMeG/4fLwZxBaT3ZvCTPCs1M1iIENSw6X+H3A8YfKU
aayhQ77+IV5VYLEaiOQWyHFN8sSsi6ekUKh3SLralvbopUeIoPOrGT+z8R1I9PBaZP+nM33a51bZ
sQbFgxkm1UaDfoC4Sbh2pgPZKyf4xcTtwqeCBpqQiqU/LRbc79X0i4i3dEvNYvia/Px6mqA3axxt
BjYjLy78BDESOmOrRi6CzZ8wTs3gi0azyT1udofIdspzHkMrFYiaZTAkT7kVKhk7cvjgvHo2Cm36
9P1Ky2UQw9wX/2PuXq0XjVI8y2MrXa8MKi1nCqIviMYmpVJYkVUPDUdwMFvrzkRPEKMAcdLqfN5w
BXaviGuGiLHgnAsEztLeDE75YOKIkOf2S8gQNuvojeDfEr4e2tTJ/NnI2nU4QB3rkL8Sj09SmAyn
eop0AdqkC9CBUrol9x5sajjH9pduYEdbLvaDlahyfDjgVaGcfARIxarKb7zPw1XfBzH9Q8tqSZDs
V6fVv+1DDNFKc/xtpAl+Cb5ugKK07xFe4y95V5JXNr3HLnUKg96nChefWW4u/tlVu8VE8hDaPnLW
HUvpBy/9o9ssG2un0W4DFXGRHbufsNFuppicGaKC/id1060UWDFwcWj0LEl+5PvZtwygOZJ2F2cD
3OhthC2g9ygRmL0Lg1jS9VGcucKmi+M8jT6uQfVunzeZg2Ia/dxRVSznDw8bJnljvIRTbcaeYBY+
lymc+/vG0aqLAtAba7gHOXK96LQbCBXGzg5HsDI+9VUF8r3DUEOlt9OnQ2aJURMGufnstz0h6cke
lp1x40P7IXTzuOQIpOil8zkYBJZfG0SbfX3IcemdpR2oFlmy5/uzx6GcIblRo+Er6cfoE6VZYFpG
3TR8SWGcO+KI5yMQZFa9r/PFWttlRs/LjSNoVzJx3KOk3o42gV3jA3ZlAEOr6pmgxt6I+nMae/Ut
080cbgqozNBRzJvJNBS7D4WVnanr03ilBbdbamLdyIs04F0Llx1sEi7tSINn3GD3o1fdS+OCSlAm
Y6BKHwDvjJGbrg9C0nBAMBd5InYp0i24fS82VOk46NZwKu2ZnrSSJ4dfu3GXx8h8U6aNePh+ERSe
OZHZ/x+r9FaBqWEbmmEJMuyrALVS/LY1GWAGEvH6e6XXW8CLkvYP9Df2MZxBsz61c2UELpzKBcPn
7kFsSN/7WjslTh1H8C1F/lPowkDV+97YGW1hcZJDbiT26uYSSX46OcVZ3ixjxTVpF3hFCa1wC4DK
Xcyw9qJAsO+gga28tLODXaUZmD8EwaAv+tDCdhRLnDCGdA62ebkyTXL3QCePuL4QMkMnH+WMzKX0
EmdlBi6n6HmGOAcvdgU6YkXX9xMpClcCuz5UBAKiUOf4Oq7DFtwa4AA3eTopdUa7qp4fz611U5AV
APcPrV4BVNUG/qGRKh/rYiGcf7xqQsEO2N01zC0k50zQfwQF0aazmNEaiUP+qeaux6R7TDNkE/f/
8XNBq5dk1YPAp+U9PNXuKsVgT3SgF4rE066aE/67/umbtoXcXpgJyiK2uvIdJXn4fAI9bRctq+a+
rZ/mHf40Caumh70lF2eDGIEEyETEABJ8M09CTmIdrk/J+GT9ZMU9wF4mah78o18H9rDODXqMQfc1
t5EaUMX1QXxc3vY9Je2/MXe9iJtlsMTz7M7YnTg0625QxiMUe0y4D6dHuVMXSJV8UNQRN9AfpQUJ
FiPVcswesazPZwMamLmOtl+8rmUoOu8vK+35tDxqMWGcXHfNiyYMV4jkcqUUCFNVGx8XEhPPkeV3
iAawVMrZrdW/wI974X9I/9f2yoVrsiqV/njdXIRjxOCe2BCyxijjALEXvjV/18H4N0bP5OPglXjw
/PQfOjuP34e6+nWvfm6EvYMKnIc3pRwPXqTkS1r+7IdULLo8Ga31753nwmKlgqQXMWcB3gsf1uSG
CcmwQUoltKne8A5ZJdpdbOdHcJr2RVuxNL71rN15mG/MUDqAMFBBl2RynBmFH4u/ye0u/uR1FiZr
dPBzFyz2FesgQIKJxIoDBYmwzXq9D4daoCu3hv8Yh6RrF05Nuxb4RZQIZGYcbGXXivmErd+uhKWA
KbEs9ZcqWVhuogXeqEyWtzLWWgk8pxBao8nmWcf7LuDYU9k1nw2SBYYR3qWRe/ypuzP2anHKErHa
bRgtxSVdDyeJtd1hRQZCEKOTI+KLiHkZ2npZ71GUiMSF5Rzp397XllfH0w0l0/KtF8w/53+ZYdGC
b4L0PrjgJi0nU3eSOX/0HEJ1/5+LBrtZkjlClarT1AIrRIFWbeMG8PXRy+26yV/z3wpjBCic3ynG
vGoERgYCJ6osJSEweE277PpWUXI59C4ZLlMmb3R0JXJ0XTP3oj6/Nth5M7xLXN5Pgg77dCDILUi6
T0bwnkFFu3U28JhkLef1s9t8k4THw68PQ4chrfjdQiD9lr+B183xtu48Y58dYCSsF1/LCaFx465W
mj5yZ63pCyk41i/SkB8wd4WjiZWT2HjNuczbKkTm4VACVkA37cPZXbqYG1F30n9pZeRfdnuQ648e
IsIqHZXyNiELubaNPdbeYvBXaho3WfBjlZ1bCu1k9x3rrH1j0fP/SeBQ3Gz2Zxyiaidt3NQHBBaB
ixaQ69XZxAuXE9gbqcPSM2430DFTAIqb2TVVPbsPv8/RvSCD7zM2HCd1CJFpgiokwFJj8gN5dcMR
rV9/W/dg1GEtP11T6RmA4xd/MYTS+hISjtgI+lakpDM1xLMnrom/Nlc6oEwMAMi2/1S+AYMvoNMa
nwoAOiwZTYK0PO+idmHtHsL9Dd3tt/7V8EPAp3pCqa7+mLv5cjqEq+C1NxPnIzD3lPoU7wkgTaqG
Jq5gtLCVdPOO1YWYiAgHzpWJ4VYH63cg5BAaJFM7HkStweYVKDdMpN31U8ANxngKZoGym4cxtwUq
pWZ8OhN2/MOXUUJxSPIifOn0DmEGJzOwKtkmHAGPoL5STW7liDlei78f3DN0ol6CC1+2t0Rt4GTB
u/Lb3lddUXwgB7u12NAXiwLvIEcXSeTVIIYKrk3TVLiBkWKCh6r6ujZzz+qI3EMgwbMq0eyWp/zb
1Gmv0GdxJw7KH+ngZDbRuL7/sx+HkdN2HHnprWtiyGNTTFKbnb2vp1LndUsaePyP5VmKCNiSKKNB
zIsU9ILjmTXQfkq1gKEPViBmBCb3coAQNyYmGkZM+IGlhtm36EZUguATdvCIPaCVlj7yi2PB+ebP
AAxz8rMlcESxMJEfcvDPDwKHUJhSfZ/VsWRKzLjM1mHHcTYTcFi/zqEUU5eRPCYz3XMKgY0YSuPr
mcGtb148lilZWhD+17ci4pKaAn7dLIZObtzdm1pR2Z4sGS7u6fBuJCi7e54jOIcXmEASlrGSVEE2
RNVg0QsnVCvco7hHBRqySy8TWdBzfCtShJmcsxihe1fVLSCYyMi1KtIq8EiGh6lt9I4w1bTz2rBV
krFLJdnn2KXLzu/KUrN7wuuurbDG+cVVz+KeVbtRVoJEpU5Lwra8QAneJAceAbUl+akkBQfDY4vn
1K6zZdkDhxSIn6STTkoUSa3Londas4oEafad80xlZF5mMTpcd3BW14ZMdE/PTOMu/4R5LoL1EoH1
jPgDzIHTvgrUThF/y04lBTcAPE9qNfzopJvk78F+YuEFmNdl9Q+eWO9a6io0EgbPvE4ciD7Urfk2
gqDJfHowCEakUluMeU/ZLhA383nASx1bFzNnf8Rp7gw/qwAwOjxn295BFkCs9TYFEIuc1vl8CPli
bxVnseYJ4crgvE9SEz/CeuzJzt9I/zB+//MdGQhAy+kme7lU+2LozFdXyJ/6WdnoSIUk9BIXgyP7
pHwnsCHBtkusF6giDzbdccJr7dmDmGn3+yPy5nI6UKoZ1285px/oNWic4EpT0yXYM3AjeTy9HCXa
4k0wdOWq1nQZB5Lv5x1zEQPFBQHuCFLKfGY/TlGExq9rptakbsYDFD9NhPlFmAlp0qm1+CFXff/G
IRkF1sZNu0Fzemy5MD+nczbCnwGtdCU3tcXr3Bl8vVbUxjxbiUGPwIzU5IRX8tr+/AaxwYjfPk1t
hT0ifq1PaFO/ssvExMu17DgR/T3uo/lSbQWO1HPUGsYYrO7dKOw/rz8A6MWIrm4N2HNbd03/O3jF
XL+yVRvxTT+ubQDuCdAareVZBZ/kFT/4jEQ0A1COkybHDQ5kOFCdYD9uqBZBGATOLhiUopg84IVj
1BPFwejSzSYYN5UF6tM3prnPT7WnTzjlvN6J7c42oRLLfWrTnyZVLFDuKcub+622+/HNwwGZAtom
fXQf8Upsh6zeefepgViyjPqnv4wnxGIOZrGc0SNSDcinwiqsPPi0n2SGAjdc09NP2jrPHkGNpBJI
QzkC4JNlDX+pv+vHH1i8ofTnRbgKPa3hKGgJkHY3EbXNPRdp/UyLU0RqbzP7kPiwQYt5ttT21jMy
rhywKkpLM7EV8We17sgduA60WkguIQYNV89QqAC0BuRlHgdGxtvNE/gK/FPqFwY20a29Egy/EkwB
W1pvtrhIlcFd2Dm3+cPwITw8i4n0j6F+TbR1YL830jyZdyZL7c9fLrEOvcEHcOc5OfZnhnCKM5dL
x30shfH0pPNwt8O797qUH52QpFM2pjta9czHRoRAo8BTsF9AKoXTM9k4fHtK0cMj/gSkPV59zVHz
6ag+/W3I+Z+NbFNJzeAFHWwtJbv0jbr6en37rW23M583B8D5Blae0yRqry0bS1CB3m8P01oDKBsX
bPlPbCj4DMjfO3Id8PH/uhBxLrlCsKnhp5s6z/mVJCervwnPg8BgZYSKaHURl2kADQkfe6W3xk/+
gU+XOW0alewCWSnsoc2ThBRb6BJ3k1KDCR1nmJLwQT+lhBLwcc1QDYM+i30YDGNYcwDCA9JNtjtu
at9E2tvkpZ1bwH1mvx22+TKBr3EH2Z4Xbsr1sbXLiLsCOl3sWV3Kiduc4mCVFShG4f+sa3QZNPvn
zEw/thtyrqW6AiGQW06iaxWknrMPhZfSqr8Raq1ddlWAHeCXUxS+P34AT7yK0sPx5lXBfCs5Ci+c
C8w9kYHL2emr6fOBJkv62OAg09Qq41InWwExmjgsWtqBt5KP6CLvYtQGAfk2Ws11ldHsCy8Nj984
hwHzrhFfYnt9NwM964FYYD27dxtKW23zyTpffS+gM/LISRoZO/rGAKM1ay7WmtRp7nQp6KI2EKc1
UhunuuJphkQxcGyJGCkH5FZMdjfVLandHCJtudESQcqL0n5BYVPG+s7y0Pu6Y1AB4VppLAgTFuyV
BK1Na1U0KC3z/QamB8cjzCHLWqj63chY9WXKjINJhpcP0W1kS9xunRcc1iOmHI2eug+mcLI+Trod
Lh4PmVxFwtkdkKFdn55hsDKtVydry3kNNTdDUxCIQV5rMYlbdnrKiWYpX+z8QPb36h3Flaac1LFW
ejQuGk7zzUswEHGcMa4JmfwpX6ihvQNtf44sRsJHCX81zyI0lheFaKnzd+59Qn4P9mCKizudOyJo
CAsXVcXnzoLZxjXkF2qnZo5LZkF63Juqx8Wmz6Bx4ot+6J0CuwH5nJf4Yu3DMHZc2Wl3PUtoHNV5
85kNByrlxOgD8inyB8Ymjsh6RhMVk87pcFBM6Un+Wqv2Nmyquxr7GD2RDExSBSIAIxANdhtgdlVF
iOWJuwLcxnm9gPmIzdvpMjG5uWkkt3VNoIlzxJnMRwlL4JzO+QMnp9CuY7ZOV7qNx1SPC/payOd1
cHrVs90QlFi80GBL2L8eEkhfQZzCZGLG7j+snHNozMuL/xFUH4EoFBPIZr9qMyN4+VmuVyqWBpdC
wM1Xm1ijUy1J9tMaFOUnYD+eNGGZIc6XvOhOpmJZP+9QFDiWVZ4Duwt8iC045gmqObrymcaaPdUw
bI3mZXF0CbiH+U0l9O5MEHFLTJQsoyjhT9gGdoI2OlTD6I+YdOKN5lFNrzVPs2Uw/4e0bgLVRiL6
HFavdm8mkI/K/tHehx32oY7JqNjjOMbsY6f0+oKy/v0jbRZ4PlqjyFo7j97uFZSWzvP8NTKjdXDS
boac//zS9BxIDkRize0W0P6sDW8ThLKDgMqBrM0QFxHtBF0m7wNX/0EnixAjj5Lg7nz7jKnnZUyK
aT2tgOmWgff611VqLMMOxohC0tTDmaGRK7eyUYXhpfz83zvY2cSsxLUMLhjGHkqUBLx8MYFRz68l
dUd0/r5nrerzU3IUrVC07MC1DlHjcYPzYle2bPLts8NmDADvNE0pRIeRVFI+sS3XEF8YNaJy5uzW
4qcJ+vFG0y2k8mOAgg4H9Gapz+lWlL2v+vt78PlwYCY+N2IboyDGO5CDKNIVmIo3/msHBghK3HLw
UEtoWybyt342QXpbMNoWaIg3sCjnkKQc4vh6qRNwT7aPWzjz4jrNF3nmEgTHo9wEvUbHLhL3xY2O
K7La5derFnrQC0afJZe5HEVeB7icsDvYpf8nBBhPCOQKS2vf7Sbs8cqraXk517iIjIsmi0TAt8DT
qo0lrFgmk5YmJ+xNVBvCixCqXac8jSWxvWZn56T/Ex57K4evwZmUwURBrED0SXBXrfJwXx36OLgA
Z2Kznh03bMY2GBYyYj9Lwp5vcgS1Ow1IrcXKcOzHBO7zdGSwtflqxNCtuJbw377uVdWUF2vXTfIT
QBQKv9N/uTbgD5OauEcfcbO4ax5ksrhM+wdMaUfpSYN/nizFH8rsGeN5xpQB+hfq9B1pNvN8NCMT
R+38f+Iqxu7HQji/iq/8fOUaWTnhg8zKttlb9/NMNJKV6J5xXiVve+MbeM0TRq/fserN26QHag5R
2JwAN+71gVDy7UAf6Br8W/izczOI7ChHpaXU+VFS1HnXKIJobKiuIGwVE0F+fGZEcEY/0TFECN6X
go3x/S+fhortEmv0iWzBwHnebgYLjnKhlF84ZjK/wX1JW4xeU9j3L2q01sbiJS+Ao0NzXgyGixeI
OHgwes6jQEspdchJg9mByYnDjfloiRzU0nFLVxt3IxWpSNsXlR0h6FYFRTX+KGsGmCQlIMTcxAoK
1jyV2yneHVMnMVzCj2DVQE/jAhCNrb96DROgQyoCbruOWrgX9cffZL3vF5fUIZe+lRhrLT5nyXu0
nR5ozxTI25HKLEdcykwaxUQ3ZicVBrC6XNow+RAn9efTW601PqlhvNhkQo9K+XUIq8mTRtJXGLlD
UrAdC7bSlM8gYMjj7YiQ23zl0n01aBoQ2UvTiKuNJ4HWp6wF8VYYZHPq/zCiCaKvEAmai6p6wy9v
iEZLhZwJ+O0OxhBJETa8VS1brpTiG8Tbj9U/c0BDeaIp1Z6WYEKjzUboz2gGhNOImEnaszAR1eOh
Qi00s/JIG/SWF39hCSjmnLMDwBWiJtesXe/5drN94zJw+eJjrhFze2xZ1Ey1knaXuESecp5DwCNF
GLHDU21a/5Gc3D7k0i+ZuLp5JIWocK0eDajFz1Y/FmLptnHqoNpV2aqV3fUmPiKwGjkn4C8Wb+/i
wHemk1lapUxr9VRkSLjaT6MPTCw7+956ZaKmv6umZoYUjoQwR4jYcjlzeGjSeSbxl6BbxrX1wLmU
OMZHCrmq/QiitS/UHSPld/Gw107OR9LOH5e3naBZUftCCWEL8srQbwhOU72zXSIMnS5SiX+sc9O1
CGiqhJdvc78UwgoGbmowGu9TgVrPdMew1T7xQzOPaq9Jv53yBs2gxRA7Pq3NrItbu2isFrm4SU5d
jC5hxenV4PPwB/PMqFwRznE1nTLTSciEb5c5MgHWN34ovMCLg2pywYnNPaXh90VNC+fSzJ8aRXuC
O0TirBVMqMkDX46rn+a7RW8lr+Hesk73uvBttQlrOIaIuDrhpscmE+ifxO40RXxQIb4qVl1BYIN+
rgOMJSfhhpz9J1DVrwoWlm7eBAkzZaSx2mfbvxyGZ83n4UXsUIdPk/OqM5XPukOrnsAnKvfyvYmm
tyPpVMyjKlRKF4p2ixvNF7HrEr0v4pU26JHKebAR04pl4yD4cPDWVMUmRywhYgZaTC508uhjLB9K
ilkYsHbbzVtfksehUF66nViyAVRJmqMnC3xWReup4u3fKexJ7Lx5t8XjCmFwx6zqBoJXo/2Ju86m
HduBetD7kA10Y6thKe9pbMZPX7urMcEIZ0MLceBc+gwTt8xWdccDKSwuJVkXjDDFRNfjekQXHJCt
6ECUcDqRwGKttetX1K5BAL4D1TdB00Z8TEQNChPPGPmQxzE6GvlXSFQ5kW08xm/qX7WIp0oHBHRR
4T8dnsdY7IG6mReng4aP/WvNZAUTS2fz0myUSeIbz0QNMtKNHOlKIXW4zRWGBq0eXxV+25TiEdEk
/eJpA01fexbRX1hgMxHOjrQPnp2Qevt7cHF+DSE1e6E06gEai1SpkM+UrAKYqNi3biHIU2Zac9X0
BTKduLZtbSUTvs6zYxnx5o4EfMbp2J+4enq3DTtGYh2IQt2zVPGiqR5k0r33w3csauWNv78mIFef
U2Tmgu8tSdbKFQgKgAnB8NvYJep1T6wiu5XMUCEE3/o1flSOD98udx+m/GdQr5fw8LJSJ9szHU6D
sl1oZDKS6S3uJdx6Kl+ujgTm+joCcyH4WvFTeZkF2qtHf5U/vfKIaT3r1h7v1iABTzwOMyB2evzB
6XNIngu2oLHJNO6vp7oKxeqqBliPXkJHpKCIETBv6SFuvGQO7hOndNuyVGAnYOQbyeJ/yH4pHuqm
y/u7txsSo6EsKWDWlH5m44rhMZe4qjwGzLUeeEokpXgbN5cLaP5Jo11YaeoPbvie0TuzBbmkq/Ew
MA/Ow4dLywzuyGx+7n3BMVYQeaNJiiR9dHJDwTvhtd4LoHBd77Vs0RB41AZFcKO0kqA5zAF5n2F8
LPHHtVEUPdIpkq2aOVz7qCe0PXjYtgHv8YlE80yUFAkj4UIq3uDP/h7q+Ux7TzRaa+llk97R7nPG
XT4SQEEB62b9CeT7oaK0SO2m6ohIGFyHSC9FWXmI0qRy9Lq6bWrYjkWtvzOjjEaNp72OyxtEsxPA
pFiUy/yS5ae65Hz2DuAhF9FMHBABBQ6taPjUFkk3oYi6M4n/boroei7wiOIKqnXag+dtZnRBHOAM
kyeqJfxxbBhXsFcImD5ZURGrT6iXM36SlvVmClzq54yy2cnIpUgfy663vSS8o4IxkMwdJ74Dms72
zld1Vr08z6lguCR0j9GKstf+cdwpejQeFqS2oMPZkchGknaOZbQGQYfx9QQv6dUKSxcQ4gWCuieX
wFcsU8mp5L1rYg3YYC6KwZRXDdJ94JDFPWUr09zmFwA4Z2zJGPaCHrPGvV+3bh6VHznsMy3+otTP
wa4ciqodMhnD6KBgzjHnNxtr/1Ue2X/uATA+Z1mgyU+sXJofCwgT2Qb9BBisZ/rLSudv4RGsXEja
aXFXZoGqnFXTHgGAvdoUkQd1IT7aWkiNK9hyvYpIZ4skYdZXFf8WPukvCY28hFT2qy23yKFwNXGy
5c0m+bMQWI84MeTf0eX7KZS21nz0xQA2OZTpy3/ScVd/+Azl1tq8btCjfei1dpp8/p46Wm5L75SJ
WeY4QQLaStdstAUBkP6qXBen493D9y1ihXwB/T6nRDm4M1Nw8om4nVDcWeT1nkx6ZVqTay9ea7p+
OOPAMo7PaMYWF9ygU+/llQBsc/wPrwAcnzBNfofoFezCm+io+8/hGbd89i050duOVgqPcO/GR2dv
VmFsLS7FgxjOLZlSJ9ynl1hp7ExEl3hanOgEmP3o/QxF05YvMhRy5AFyIv6LSBetjqqrn9sKqWC1
Smz4V3ZYg5dxBYJI1OMjZEE18qMrmxuV6dv+3jeW9mQuTgYVg5JSYsZnUynx8y43DMBLxjiZ6Rep
xFg5Q5o1ljmlN0hWZbn4OocId1LNPHJQFSG1pPIzYFORO6PS+kDzOXBKEkP4P5d3leafTYEXROwL
VxeV911e1JHEJ5rGcA1s3JnRZd14oXYHE9Tl0Whsm5GdMdE62uMgutdpcDI/0xlGgTvp6MVLYiyG
Q1QjgJDzBCYEotkpyeGu03XDluBySklODlJCkF1gTDwpIU7I79wZkICEReeCpCqfmdW5vov0Vtti
Sou4TJOpR0Gvpg0FOAeAFiUmVtmhtAxVXkZjZuhkdBX9ci7l2QnAVsklVVHy7OozqwLIzieb7307
jH7sAdi1w47XWen2sfAl2jMlEmJfEUjBLgix99koKdH/PRQM39vhTYEHNM+u+LgIk/V3yDCJBKNN
AZdalmF9AkVyeljzoD6wHmN98Nmt3CiuP03/l/TulWJEziP/XH0fTPmjxVM1Or86Xrupgcrl+KyQ
scOl3sODDEVpHMjzyIEITlfkMlEFyuXkBy2LDA4nr4aJG1acD85dvDxMkzzhfxgJ+BkHrcbfWHDG
9/UTc50vcAu/Ez0q4gaBZVgsonZGmQlepruCksTfgI8Zu6G5NFFOCq3S+iLvqEbwXM6mkSbVQCyQ
lFliXXEDaQssDd05NbJhpU6vX+dAJApN+NgcXl8om1qyP0Xv7i6baCvHerh7vq9OdsXLYiLcIMv6
2dTZb0tD1WoGcOtxgVYJXKg1U1rMbz+noTpRX2pqTseLkumUP6dXp2hHOLwMgIgFGZUQAnb7pqe3
wCIQP9u+V4+3Goqmp3zoFQZ7CKuSRTdUEbcVgsuw36rSk77oNnoDSDlV16KgWzaZovFCLSUXp+5W
Vxvxi47GoRxLIWO15qucTzRqZwQhi9YhROcMEA+3e+xUuF8gWbSSxqTyYevMY6xjpjgJQ7CH54MP
T+1V3FdidJh2a4bJKtmbQN2GnqNl85E0tT62SS171ZTHEyBtvkEylFt8B8d3vGQ/hRHvLMQghc8R
TFTQZuH1IwYDe3ddLGRgOJgtNbBw390gUaZ70DHxynC7jWVRkes0K+3oaL4tGTHo4Z5Gnqay8HG0
1IupxDpUWZwqiEqbpUtDlvacfsvXQjdsypF90LorZAy3mS/cQhQ2RkDLt6wCEuDTIzRz8vqGGbH+
8wLF1hy1suGbyKPD1B5Q46YhYLwsDFMMb6HUTxNOKUL9CQQKgf76qeDlX7BgGxVoJnU6pyXRJT/h
guopCek2QrWDYgD/jv7KgL3WPDKbBSRJw6ah9AdZAPJSgntGi9x6VEjYv3DyqslQaIszK9WK8iDv
SJ9mEUCihe1ATn/bdjvmXUDC/T6v1JbO4MWvpUvl+0yRBnHw323uq3s1xVecxvDUuvXgYr3nuK6M
Lf4nhvFEdWmgYkQuDgpUwvcKw7rjmmEO+s8MC2uQ5au+FRafTZip7CFAZARxa4x74y0Ndt9oSM7X
G3fbB/0AoWoMEagQkZMNVg3gUu7MQsb39aDco/YCJu0mkrGREO3ZElw9SPwW7XCsc4ZQ9vRpNZlu
sJcxAXFbnHrM9WTKpwHTjAW+TfwrbtlwXCI8l4rpjGQfyl9n6F8WfQgElAbK1hjfgL94wN/4dMXY
oCFYTJ/4apXywwdKb38z430PIYSHRifFaUIkl0wOUOBpHLycZJ8VTr6K31jS5uSLhkqdhzWcgtwX
dIridTr6As5q2dLKDErtFxAsyfMX+FWXrFy/S0TWkVV15FvXjlq4GATBmdhtwS6OMYxM1FzuDfqK
aBxLsbfDBMpYVoOWCBwXA/RRCsW3TYhfCBEP7Lodaw59RuAy6BrCCjVdfHLOu0l7z13fk8221+vH
/y3x16cTLpyg3kIGtR3sTiaNKNlkHHxCGNzcYhXAO9RHg23BYkEJvZnCXMuRWW2fMN4xZX4tqF0q
f/Os9+lm94i10ht0Zyl+953/Bljc1g7rqm+iiQ5kdtJc+Ena33cO2RXQx140DzVp8wMKvX6RAWZP
HRwVs548imo462hzvfveomGdFRG9x7LuNu4P0glQlKqwXWbbg43Fl8TCxsYPsH3M3V+ZelXeKpOw
yQWredBLyB2BrMVfEleBIkF8cM55XYXX0aMocnRvx+OdAXbc+Wd6hquYBq1zRcHEt99Mb1j97jdL
7om5N3OsGtAAR0Pc8/UGDDsJv3a59IuKjxOcRgakHEA39wE7V8A8OhENCfV8axISUPsloccNn2pa
Fuc+zjWsnWFAYinUmORQzQNGcztLJ7VY97QQttaDwME7eUpeCjZesHbtqJMXVA2VbD0uw73W9yFN
ldbbSUXNXVacfa9ozBaWKYcLyjQXF2Bh1pAyCp1sglHwKD0AmCUV81jUXpuibTDODf+LxQ2PnvNp
nM+AJzNCza2pxnWwMthH4OPDJLPnVCWiQtBQbn85Qfn84Qb1n4V2uVyplCOQYzIKCif1QXYkc3Ku
vnfaYhuSeue03vPXCnfyBnrRwvcNNAp+OJODRqHFP9GsLU+QpjiHDyNmvA47Df9xVfouLnsMTw1A
PeHt8rOvykEnaJNwmMpSjWrmedDmm/RcPCjeWOpsamV/NXk7iT4ArAq3toP47ulIkvf/NEQ+y4zh
UE2x+xLIhoWE8WrUFX1TNZ6aBXe6Vx6I5RHSl9lZpbX9dInXSz95yEu1AgsDAX0sA7DVafU82s06
Xz7wJhFrsvgB0OtRybf9tzMOtV4AVV9sbpnZ/eQvznWSSeiSrTZhSOjrEC4MBBryVxCKn6wTkNp7
MCkXgeRHjj97hdGvtG2M3y8hmdGPr4+GxNQM3wXvOSzZRrSAsWW7w57AuDz5wXsmSXmXKMtmifx6
ZaAcJ85+PfXMXbMPZcOGq9+/mSzmhyUIL9hCzzpc0lwlr+GmK+g+g0nLJdhmKyTXGZuzxMIZr0/I
kaqLcG0bJ2XEKFA0mi1phMyijHAST8JqVV8kG9V6VR0LDNt9gkXogbEwdHIQYfccx2GeJw9/+TkK
e+3iArUGcPf9jJR5LK3b1CnsXurYgv/XMMGfFxM8y603o9t1Byj/TFeCIZU0Yp5HBfvC0GEV+5fu
ju3q7TUQEb7vOkXS9AIZvzMZ/SYXtCN+r/FvVEPNJs7etNNuhwggn+pL75OXiNeEZZOXZ8KNTKqM
A89RiybEkxIQavVnSb8CMXukj3BDTt4t4uW/Sc1omragAUnHvm1GE7cOHiwT3Gt17qYGWzf6kZ8u
MjuWfcTXCpIgcS6UQzNDbNUNA33wnJlUY5efs2q4crjRITAcb9ZeXoP2H77kDwvGqm9fO52pf8jT
aWlFDzhZKQ6FKcto7gjXgH5Ldf8z6NR6KhOg/6vRthwBc2PPniDR6se6ASbJrV6FwUlfvlYQB0A6
N1etaxusEHrKbsopgBE4T4UuUteXChr59i1+j+9x6IWNbrvkakjWnoiabI2cuUjf4QLyadweySGe
g/7fqXjXp+LBzsI7vuIC46mjlJoVMn91xjShvSgU+1c9wFY4ykcVTKkFkGCZtKSjYOYp2RQpXDWG
LANE+1SY542LGwOomXmZoU5tcubxYVca12p4SaLvflWGp5qm6snAEqZTxsjUetePe18qA7DwERMG
I319vsnIrhRGo13x5XuA4jIRPGPNcITEsJkSkaTRaO4dO5DpIJEAsQqBjFfDPMSv/xvQMc6ROFcD
1yOKDhErYlUho76GvHxl0aB1S1FUTbGdUtSBxldhZMSGZBv56eVEY6dW19tQWeaSfDmJLiLvEWV/
tCFmZHX5/P9AMqVahyt35Va8jzYI4rE9nuSYzlFjgSc0rorvAz9/xLABEX2Ia14OtJ17tgbhQgOv
ppRNikaCbhD+05N9lZ/EI6PmPN+ynIDh9svUmvgTSZiig6xSVTiQtJzoxa2FVdLjET5TcvUuWt14
xFPn5drvIGOFuowjSk1EQxnb7lPH8iqNR5J3u0O/ba7fJx9Pnk6uClbFUDgMpHeVtj3srm3aZVZ8
5rzcgLt2zM8uxAtINoTypX75XGRmqhgmOU6RuJGadknMx7kDT62egQSt6CKeCwrDg+Vdv6lOjuVd
2rAoFf3HCbUKLAsjUWS9WQ7LlQ2cqeVT3YOuZnlXDGF1WRgaOHsCLVgVF1WAGQ52hNEw5v1WuwUD
xDSb0GiN1MNz66MeAP7piTxYVjZ8ZBSvFPLQUx/lyqZHICESShthnlPfOiZDMsv4GRSWtdwFGglG
ni9ouDEwVxPURj1zUt3/IIl5b9YFomjfP/DhgcAKVMZtLfwg3Ib6q0sDwwcyr4rMZ2w/EHs4jfBe
uMiDZPzuCBE5rAzGRp2h1H8Bk6j/DueBVmOwWeKcAVXJO7JJgI3tJq7ZVnenXHHC+5IO5E2Pzv8j
Uv4rgYSpU4tde3JD2oeFHVzEnzpDbwNeWiqCbvnr6MRBrIR1GqdieOTM9+fRw891zA3w9BkRSJYA
XY47AvpwyFRVtbEJEGzuubLhCNCTtCc5mgBO07Pcyg2bVJn8lnqH0M3/NyoVtnLpMT125wXkVFp1
SN9JSv36x6+aREgeuGXxO/FTlS+dY+TFYFINUigHyhzoZaKYC9pWmo4lVSvYjdO6JBqLUDScMKQb
UF8BXTZDqYLIKvc2tiHK/64VJLIlOCqlv9pSVfks9XOHbzvCOuujqvavSpXP7nKiO7RD2qgBIOJX
8m1Qtw+F4on7MMrWz+DhSdQGvaycsMW/UKGIcLNzWSm1L/orOifzwVp/WTVbkrMIXiwdgVV+WTbO
qaIuqS2musvuz6q/7TerkKYAbzC7ftfSVCoZbJDCmgMDuGOfu7u2RTD22h/WSzv5uF986sF2Ywak
9KTBhLum9jla9Za5SgHwGqkFOKDvkmSiCAM9vFMGnZJF7lujPNwHWQ1yGxpoIBWTW+PpH89D1cEI
bHTQSzCsX8gBzJYm3pJqryQcfmvLvg8s9fgP022T1tCDyzGBtRKuVos/XeYHjHAghytuLEWwAtQw
RN5O0LEjxuSiPDZV3NXXwbHGKXnov2HgTtDkdQzvQP+ZMynFkFjJzyW5i6nRsqxycc85lbbWkpNx
93WSsNiOtNDVMyf7r5sCwunnWeNMclcfIdlWZFNljCbTmVGiGpw6+GAOh3i/jGSmOX2FkfcN/ptW
0GFFZWaEeD8ZDczZCDu1LPjZus73gVvgLnZzAu08kmBK9akx98yNf3IAUjXp5qcAOlMaPr72PC0x
bnWG3mWD8onkR22jkyfzEGV93WqXf/gdeEJ+caOxRWsvkpZ278O5G4FpraoKA1tGJI/f0fWts561
bIsftk4jM5q2Pm2X2HDkQ9IEVHsUyzzqGb1DzVEyj5J4o/6U/OfUUBSaWdJZ/CAHDIYZYlpQUQVC
yLyidQGLpITAwE9x0r3eeQmF/+grbxqVdZnFl3adHYKCpq9G9xD4d5G2gtRjLMYeTbjRJOEbEpQX
aqjVJTSM9wFwSRK/cWNcfwJXA6mp0IKf1IVazQUP1w/VDQG+kZ9FsyIzft5COrn/2YAk/Pj9P9dD
wVBXcBBblB4HWNdAoVLxNCZTBD30f0n7jGScJBjmaDmpk7IT2bZkrjvi9h3x6+TFsHZA5DpOy2Oj
tVSZUv7TkmqXFxE67kbmxnCV2QZhU44WDrAbW2iDLxhQmRaKzX4iINuh6ZrIXdphHBfT/2Rq7Ofu
ewn6Q/9maQ6iElPqJ8dFZO2pPmXMYnImtFnifvr3kquKj7srvK0bp5UsBEXNKf00X4fZKZXSdfxK
vEI2mDMdHl54gvDl2sn9ukJEutTV3UEcw5qYTNowudzw1RQO95WHnUfRBhFHT/QyMgL7NfSCW1HD
Tlv1bkZTgl9VrPcKJEmO6u0vz1TrN2ldFuacohkfh9NhWXJZVlotzxVHRUAXC3BE5n52ia7ZLRHd
V3z7+A+84C/c03qCSm0vOs1f+aNSiCyaORjIy6FTfS3/A3KnFEf5flsy8ADd7OJjH+hFC7lJ2m/1
1yo0zxMMG1CqOvtecO7b9pRIdOPtEXzoeCwKQ+wHplSTMKYwsXM9MFJPVt23wVWi25AXQXV/jj6C
DW3hDWHN3URoylQeGta8VqVPPRYJrv+VMagMQZxW7G3Nbb6hkAKeprQxbV/0r3mfMcQt5kVrOLhc
3qpC4OMXrRK9sDOxUTPa3wnHipOzSLjAo2BtoYsY/TH1f59BtX6pHnS0IyqZKoqG2ERv+gj8980p
MTaVUztlfBa/WMGu3VqFPYMAyUGSCoXRY1mxE4ommIGPtQkfxLLPnqt5vpGm+JIM3bdylEutNceG
jpJ/DXbMpjwYsg/YlL+KUSbhqKLfFLR0mQjgHMryJ67dF6FakRe7kPYWJInPeBiknjzrqhaYuZbT
1tDq/6LQpyaVguN31edzTE4jGAgDg/ABY6k16fNvJtal4Oo0/4jF8EQgGYFtPnY4/9i38x9Wiycv
HXVcA7KItkU09GQ6xUtnac5ENX0XRX4/IX4HHTxJBq8ItpIhBw06S58PBknSZtJFG7R84XYtqdSy
Q1cbxo4MSzh3QjARtv2eie/aseZ/29pz421PkT6eh1l0LCuNPvoNceB9MAlDFZ5iOZr8CTJA9Zhq
OYWjwAHHxpv9Aft/mliJUYHBNGV12/11QxJKhKU8YUbmpwnELDeI8HK+xTnVsExebWvCbsj3zHn4
aXBnzHBoPZCPmot3y5uhXkBe8HUGdwLgyHVQmlSE4Poj2kz6G9UFuxKzqbuLCHl+lktTuBjToOv6
IUj7X7gVfEngC9f/XjRorw0yQa5zASHewaXDKh6IrHVbNJdQaA513CcnczZ8UqY1uP9AbYTYcu4A
ymnRp7W+mXsyT62pTlUFf/WToziCva28vflgPRaiItnlnqfXxHKZ+i6ybBjKm4YNYXKwTCdijz63
k4RtHV477uuYAd4DZg1q3qj01mgYmH1dGKcQoKbx6PIBRy5NjfLM8lY6nC3YkLdRdG4tWKEvfrkg
2xzlJU7p/OvZ6zIBBeLyEXL1K7hW85NwPqYWvIhLWi8CCiktjav8xLuRKXoxmPuLI0lCT6mfu6EK
YEyfdg24N6DuBaTFxu93r1K5/LxWW85oi9j3R/1aHqhuIGV6JXggUTNS8MmPkvraQ2shEbqdcKLG
7saMrX+sl/d4uZWdYosfWca1DyfjmT5Xgv7yxffFMi7oRoBMzGCt23osngP9psaRP+udcw9Lc7Dr
w/+NwM6ex3kdlWLs/Pe30EJcehFOepLdluOkl8LSGobIkhOZnFusy/EN3UE1aPAsKEj6ElcbUwzn
gUcQXXB6mg2ghGG8BnSHdZJO+iAfMQK0gpA3E/gm6T2vVJSmxYaXCWKb8GfSxYOS7rmx+o/ijTzN
5bur4vBsx8Ra1Sp/d8v1io6DWCO1lOamrlLPgpRI2kqGHRxdOXRM3fzg9Qn/8yPG+RrCNOBe8vc9
yXdRazOtzFY2ccJoGARpnYtFrsZDXZ3FhTP4aI23dyqj/EE6LOvi0/udBAAfOsz2QvfG4T5Snses
vOHPRronLYKeekXl3Poy99+BTKlH4dy7ymUZ6Y0BVAcbtft5C3IxhwhOD5yeX9cCxhmaggDMG9RP
EXoipbtvNQj/8yDguAXn1K5L36ZZ9szfW+POOfSDOUZP9g4dymNW8Ip9Kxo5KpVuHDcioOI97a5V
GGTv4JYSnHDtggqqo5XdvmvQDDPl7UCuSfojYPphd+R5FFY4p6xGSJHpJkDanYGWJ2QXdAj/HCqw
Kor5hHfMPvEvw+Sn6OHiQmfctVFgmL8QhvTWAsaE8s0+IKrc+NCvko6OfSCIg4TVrUfptgYeaWoH
oSaFbVBve/F2J1h/QRN2NE6Wd3B4ZEIyHVjIEyg+VTXNPuMxGmEzwK2nYmEqup1gMfX/DEgtjBw+
km5wWZb9vTKWEgEycUEVtVTcLRR7Q6OsMU3ImLEcedElc6ID30vzNNvwVxZEmUBczKA1s8bNJeJd
gjjKpTXA1irWABAQMexzR6bb0vF3RKiuuNsHNfD9ZVYJJWqDPBKcxWAcmEn8PuSx3ueYS8yVKf2M
1JRAEPCYduVKPNUpmHETQybPQkXpLtSPfPDCO6Ft7m34p7SgSHLY/6dIXn+8YgvJuLnjS0XtSi7x
kDIHcHqqnUYUJUsLraHC3x7VvdqDO3S2aVx5qYov9Xv/uxPGfDiEXwbPJpvE2+w6mWoDIfMGWDAs
/IXDVY4C3YJ+/N17EAkHsBifO9gwFpzwzA6lyfpdu3AzFvIgOezjq+hdpCstJJMCT9hASC0I6aJB
Toc56l3MtDcl6opqDM9M5t5MJJ0t65XzPg+iGqg2aP4A+DcM6bSPkCfLXaSJw2D92sLEiClQ+zX7
RplaXZq/sxbZaaTOP0PSnL9TrLNvgHKMBSr8ya/uBbuulfiErM7QQtfU811XHcR36UMXb2hAmWDf
grZ9W93DsLQF5pNVlhlMzLNVVgvcMD7cvnYjFXTPbIGLV2onZvt3yfDLzQ/mirCEjG02TPWBUTQn
h0XcgwqJnJMLqr73KaoGnwFMafBSe/zBNLiCr9yIvaNoOkDAtgmmfmmTMfFoTqLovHf3LdvxqWAf
QGur6W3vO/XLXI9AKIxYJCH3DwR+zQmw5X0tXYjm9xlG/h2b3s3oTvaOOLQAjfidaed2cpPa8FA0
/B1vRaVW6oDjS3emWlWT7ngYPti6Fw1s5biQ7VI4FGNQNu/ac+j1ibX0Y4fWzf3SHO6fIL5Qcjyh
UiUUjuAfOvz9Kf9d5zHt0xwxQ/94lptQ8wr8nYucaOn8pMUoZo8XsYtD4MYHwPCzE890hVMKl6/b
cbSMzK1hhRk1Me671qOTRDwFBGKxrf9yqf4YLF563u8r61m3E2wf9PRPUk/NGG2cKsid8lbXeDzE
HfVv08l928A4cFjHTilITdO2qCwuRVMwkTwJqVgIppo+mfRUuN2jLwD4YAjjqGuqb3ibCXcaM7C5
b01rwwxSnd9dw3Kj079ZcOM8yxRdCgE1CmjftFYSPAeepnDjqPxsf6WtoIzv5t+LjRM/5c9IC9Aw
VuCK4/LEWHVdtuXHDF7RcK1Qcl35FzkfU2O7DopTPY1OeGmouTlfMItBWUW87twzpSidirxdHqZx
r0BFjWpCYhVjq1HiwoOEEHHMZTJGmNbaXdGsNKz9qxgUe/QzQh+TJ13rg1UN/WKgxKOdNEG0jTMY
lvEC04w+mMEL/pKzGwfG59uGe+iF5kzszBDI7uRKu5u1Bf11NgtY5UDDng//oiHL8Oetw4DhCr1z
ooACJ5vRWTQP5NgnesesNUtORbj+bq71E83V6AulWfRYlrXXSp9NEAdaEKnPqn6ueH8qysDKta+L
igtjPP4EzsAX+H43+gWpJhVwSiy7IOTN/VhoyMhIY+7r/KBiqUxtUuOglS1jZD/9bgFQ178b8BtD
6HyB9AYEHs7uZ+N+2n943CdOMhoD1vGSp6wMfoCwqsfdcjkePuA1qnTyhtQXTDigz0Vii1HQdZeY
IWzbm6rl4MpU4Zv7/dvxKU8y7XkBdd5uZKk7LmWVCDSUxBB1lhMZ7l9pvqwzFdlF6QOiU0sxW+HN
Rg7H3Oek5BUHRfIYGjIPdj9gtHcY33pp5IeutbmlkMdGOpi2TB45oH6kTlyRpnMTY18EbK1LxeG/
Cub6ZW0iUGTEae1C0QcVEUd6erkxMiouIW0rkZtN6vLSX7rP9+2dx+Nf1CUP/8JSoLzIeoGDmI9J
lOaGYLjlwdWP78zTf9w4vW9s2usLgZo0CR0sXdjzxVEEM9s6nrkgQIhvmNWZIGTG4ubqH/Oy4fHs
6hS7cqHiHoslVnwJLLEbu045nTgkP13cff/ZPrahBA+GJmQx1yUtaexZNfQVE4Cs9Z2mbHOt1mXZ
2aBnZ5XqeiQ1DKlJkVb77bcJmsaddRHMMeM4gbZ+LMpknsC7LOl98mzMfo36o0C79JjLgZuJk00K
xSAqlE7GvjrdPQu9LYZX6DK81Dw1yIkp9RX81hm0x98nzpE7Hf3Lf86nO0izFeHNZAP68DJaqGrO
p395FHv9BhEuezTr7dlVQ9Rs1Cb11lupsIrYZ4hsXoX+LvNbk/epUe7FC+8vF+geoDNB83knAORk
bV4yqnGcmKzWHcBxsRZSfZOiFYKvFFnhT4JD9DtdbQoBYqoTA8cYlVOhsMuERoEa94woUG1gUc0P
1iQAT07Hjac5ui5y9YhioIVmH8Ak40au9k/KIj+jNNoACLLicKc79fTqNeQ0DxrBsaQlWopb0s2s
Ody6Ac3sXPW8Kxm96qyjytNPc0rmcuhZLL4Y8KkPJ7ciaVDyLoEnUdjv5d9+ch1XpTqc6p6v0Ai9
Dcw6Ylcxi5otZXZB5vbEOKF3HUubbbrdSD9oDRrnJGRWFo77KnhRPZQsGePB7pqC+WHwTot/GWL7
+ifMrtfo5fw+lMczWkcUsOxuCahfUfRaJxgZ1U/Fx0BT756tdeif2LRJ4sOJaxTUKuwIc1FlJVSx
zsZhmySZh3aRGP/ovwvQTyf0/Uy0YAytfyTx1ErCU3YjShPMEdRGvjkPOX+p9Jg2bxLxGsKE3Rma
1EbFhgxJerzP80SIN+JmjQ5vOAUw94YHYhHhrYf39dSZdFc/xuTmpGMVhtW0RsGKjWZwcQN8+G+q
4Q+5SiUwVy0pavtO6WO2saTMlZb5AZ3KEMAgSnFuCpzD+5pDlBnW6SgdX+oHWvuFSjYlpaF99Wuj
NLm7Tay6iYQfeakg8aO5nRqDke79kpuDNwsWCzdqVTwCNFRDCjm1q2pml7o4jYrUywA2y5D3XUp5
dUOz8iC1/+pn7bawRpotc2El2yEnzPnlPPeHb+MOJY8BxXe0O+DIdbCR4zi2WOi6BYmpaRp7ZRVx
heBcFE7vKA3eNsVdIGVnO400IV7kOoUDUquoXYZq7RCgGov8WcGaCvUtKKFuSgygryNXClGz276J
Jkp/HPNdJTgnS9bMDHx9UWnxeVg+ZV1a7yJLlCiskMzqZgATGVOQ2HghZ4kDmyNjlLXGd5oUUVf9
wDEWQAqayBIt/tLDAmkWsNEVTSbwyBwORhZlhGH0Exb3Oq2zOyEyl2qI5sTbpXI2/7myvb75Z2Uo
xyb+iWbdKYwfxQynoO7xumkiFbH355ihXQMmj+LH374+Sb5pnyqW9S5AIAsT1NzrxYt8sghkAb7T
rjtExAYmKdBjB01ASQNB/v7UEJXq6vHrg2aRbp/QWtmWikOrkwarIBEHw1Grmg+GIrg41/pHkV43
SjZB+55GWhTlSvXvV6SJMjM5YaprgV05lSbQs/GUL77jRt2wiKbdTory7igcpaDkOoXUD/0IgycW
dnz/OoXxN3YrMwlwG1nRiLXUURmwM4LdScFcgirMVBL+pm9uDCnXQX18cK3GFSiKUls0kQYIQsD5
63bwWOt5esruJ38TAHT05h8nEggFHyM/3KExsr5qDpN3mgq2Lwl/VrZZz7r5qEYi+5U/0zU+wqy8
jANGprfMU4hgu4hgQO6uGbkXtAiYS6JqGSgB86di1B8/l7YqHpHfQJAUKUPpcW61jQbNO6rlLEv2
PuBIEnPJrJaf48nHCy5otfiYSOot1xitJ3xeBl65/LbHJmpWaVhxBC8iPEAgZBmJmpdnxYzlNjAO
Vx1ltVzTexbIai7NBAXD3DjPkCcv6shBt7TvYWA89nJrzSEI9eoORIhKE7P/2PamgBaaZ8aDqgY5
wOkxz+hpQzhQ2JwzBq7vlKelbo5TuXiR4ndtQpB7dX1Eo7auFko44IB2BxMrVjk2fIDLqkaytcFS
4HgNqz7rGZDpywvkCv0qDTibt0uws9biMXuqx4ApkWOHHHOpfcd2yyPs2zZiWC+LTbFhJcS1JobR
uf41oEfEmMbw45TxeqrJPLj6A5B1mx3xNGNNz2fW6Ok5MZyi+PmNwO5vGamO/s/+EYAtiZdmoWV2
eosUMJIUXEFQtasDDq+OHp2vKUwOPidtF9OVG+wu+jl71jtiWstdZNaggXW0wdGlPe5CVCcsUQWb
rpAfiR27J9WM4BR74CmwSd4S60IFVBhfoY6gtIQ3qRmNqikBfqvylMGQaYM9IVztsTZJQ89XHPUr
V8UzTFJIpTPvuTUQH9MZ58GnCQ1Hh9tiROrPCsd4T67FBInltmLXZzAuqgMInUmXwAynKXYX5Yl/
lL94ffy/uaiD7+yvZ9Jr0qBmw+BoYWCCrFRaXrYeVNCk27HFCpdGma0PCXhht0QZsjaqunf6A/YZ
MQ2aQBiCFang4pmnHtJcp7Yb1eRMOzYyJAslrX+yIDGRGTstNJIw7tmbm7oc80T4HzU2hwoXDAMW
K5UGFk1vb1eTfHBtwvPCYN1veic/HeR68k+aI1/Re9F2fu60udWX49ZxTVI3psZILmesSxAVeFcd
XfMB0QL6kGWGtMegmghEF+QtX0sRLWQxBWywDZjVwJAZUjJqAQYBsl+/JMVLeynzjHhgWv4Pej1S
kq6+BnTulqaDnP/TLBIGqPWnDG9MzdroV5DEWc2Gikii2oZ2J5R87bw6EnGF3zHlxXuJsI+NZFrX
3XKhD7jnIi4KwXi2EFZMNidgmPRolEPh56iQPYLFfdy8bhBgjf1/Pz9pQq9VIcveTYegnC/n817A
XMzboOvkwenREbcpGdrpIYhPAXPybuU4KcA16RmtGy08Rr26Yi7sFiOtObBCSVXqXwWfSOW822PS
uOWGYvbFkUArC6noxM1iF/w4FgOPraRtNSTdgl+tHB11P5eYobJUmgJtyO/wFvAcGVe+miXpJkEW
7W+hWiPBItUocYbU9RqgK4QP6yQYkV2NBibELUbAXdCsdkL9KHm4SbFHLhJlUEwyEEcc5mq0pmfG
br1J10dzcypJkV5GwhzUYn6S9iazn6TE8q3vON59G1zbhJyc+j7yHRSYZn1WiIsnleCbOlk35Ugl
VV00RRfwswWwGhpw5hEiMoj1nOun6FNIMNEMMf2qCkkPA1X2ifRTVm1G2DBp2e7vkPRT5ciVqkEx
VD0WyH1dTqVPrHUUiYMhvzGnd1dRsZ8YvQst5gVhiqSyfTN0L6L89XeyQtUMlhtLJG+qUB3zU+2O
Moshy6LM5vWNA8qZbDDD4MEWVPfEHq/NzI7+NVhz05cMTw4O7adi7L1AcUvXXX9ruD+hlJx3F9iA
v0/CX0DLzIspvNy5AwjDmB9HezxnfcRMBVOA/HNq1ep/LNLwZwvWr/7JN2Bmh8QhFvJA71W1ns+g
vkST5pbgdx4xAWxfcNnYXE1M8bLve12rnEoGHuYNmGgW1FN6KOlFJoapYU+imZKqQHcgURvgGyor
uPUWfld/+FGMKMTLsG05DkrClZCUcTO+88jLs1+sx752nqNukUb7624F/Pan322nyCRcOACfs9rt
7Ugg3cRd8U3qeDGb7Rrp54MKCy1zHsn4Cfh5ERtVTdY8NW5HVn5oZI+Eafif8wtcbQibYuYurO/g
T0+uBvNrUNK1/ulLtnaYk4j3E56l97kx8g5M3UQUCkrkKzcabUEsDr7XCFxlT6b0PytTNRCNlkKo
FLPG7THuQRFiX9hUXCKu2tdN9fCUqxdjCSXhW98GmngvBuSn+Nn437veMaQb1tYkBIKpKk9/Pe7p
J4DbrgKo0WHf3QZzxERIbU+LHBg/5BLvpJpBV9HFsaHJ1WJvwr2OaJ7PNCz4gNt1pXf7WGqN9paZ
KMR2t/fwtyPMiyStHSRM1NQs4KhEFeNd116cgU00KhNI+3qaOOBZb162zdbf5qETsXk0SefVqvef
KQdhSzl29GfllvnhNCVV9Zwav1zXKA/p7FE1TzOptyX3YpjNvLBDxxc0FzFuXNmYPBaLYYXj28Uv
zUA1apKZX+f+nzcKBMF4cMjQgXcyRGyP+iJAkWWVhWzu2pcMUDhzU38QcR168N4FULLCiqlQQHl/
Is/gODni72BQMiSfF3cFDSbCLN0sCnyihUhwj4U9LTjGx3vc1WTxYslhIxkF6TFHGOjeolt6FZsd
KDBn8ZfE6ZegXZYkSepgdIiuvrQ4ifBnF174QvtRUMbpwbXc+rj4mWg69kM56bNgcR07FfJBooII
WR0h9goUJ93rtYvydnhj8xPBRLQkGBdotmPk3bF5rRF+CCbsU9Br+5qmzJFBGETutkwGfg1bz2E1
hhsYSAGUP/5QuoupRwUs8Icbu6xXq3kaijWOmlyETTSXWY5kt+ZdF6QeejL61OTuz92vMbdlZfbH
GRM+jK8IIRxsnglgKl6B0cmkzTN0fbMRbyWMzOXvAgSaygRydrmO+HBET/UEm//QjsEpVR6c2xw/
THCH7LACNSb5EKCcSkMN09MbzM9jrUq+tQ3O5rY1QQIkJImQTrnl103Bx/aemrYI7JrHEkHMG/Ln
mgn5Hi6O0JmRsL0UZ4QrN15PnY5oXMJILYjV5tTGUC7AqvPX0WHO6olBbQfmgzJqhm+aN/3+7R9U
Nouxfv6RzEnsvOpl2Yk6IxkwGHapLyItCa/stZmvhnNHt631MSUB4n3hOFpw7Q5HV877hO9R+f14
vUQbwIU6jA0vGI+upCbgp7bFqsTj3fqUdhMYzVXWzSvB4IixgDSXJzjqtFYARA6OiKGFdRUvS3Rj
ehwo85UHB8qpQJPKNDZZZoPYDRJ/Mlzjp6KxrU383j6LowTKlE7hrp7mfcutlwl12iMZks1FqOni
STvWNiyoKQqk6KZi7bVDtcBLsbo4x3s+7GTBziqDX/dD44AMD/9E4TQ/gq7vrbG+gL+Cj8Zc7Yes
D6V16rjDIBl/azmkyCrK5KcKrQ7hCd+kbEwNw2pKuaL3YuuzIN1aCpzHwiMT05QxEl4KsEt+YObN
chZKjJoWVDwunKhrJNq6EiWmaS8d+GDOqgm1cmUuetZIHBQ2wY1OKGzVvJiyTEc2HVIBEeP99A94
NEhpx+F8OfEj/+ra/6r+92/rm/g4bxG7nus9j8RjjpeYqWlrUtVVVv/qlHStM/CJKIJIBVjX4a/w
U9bxBi/ueknG8Q6mKEEGs1X0cPaosUXlUVWNu88rSJiM1gN+DZqFl1KjTwQlQugEMAFhKl1zwvwg
ZLG0gngYl6L0NmXS28oJZYO5nmEClKd+O8fF1pasRlFoIL8hNCfq7hzMx+E2bDPVnQ1lgQb7bHit
UBlW0cU/r+xA/0jl51A1epZxeLH5cbMwEDO3d+dS8B7b7EDT3ghtGmG+cBlsIimWPFaI3hhp/xmd
3xIxKLCBZVXzfNc9jXPO9X4DC7a4U96YM5QHGQDEY8e+JpLwV/NSHWNwFGYASZLLtWZSLh9bdqUa
TjrEoSfNGYdOFKcsRPXYRxVj9CDUJlJxJhaypiA7FZB8q0Ter0bfiTPDFhbbuUyQL3rbEXlqe2IF
Fx5HwoEvguY3M/u/1G7Q1EEg4+HmO/mL+LYxXiBWurD7gvsgmGWGy1gu32J86v5Mf3OlJUazTXNp
qWbYWk0jY3BEPHG2Du0drx/T30pratK/zvb5VM18sv7dQTdU9IjJ/W20Gm3nK4/quVxJPqLsRIOP
jQIRyIbPTNr8FkL69ITyAAsg/s5ysbcXevOSdM7yaZFxwvdmb96MkKsTuTF5GlgKXQiAbSH2GjVb
Ge6k6Io+yNgOPHX29usJ/kAdhaZVBmPeSqPPiAK5c63gji51gyrpNDQAbiiysZe4vnXSEPpGvnFd
2pviEdue24RCZeZmaR2sz7IJdjCKnbDVTR7sahLViQbpaGis7v+e1b2Jkknftw30amPBC44HRtB/
4Ofyr1EBREKUXZ1uZ4X94vLnl48eekEb4zmVj+ui7MTUsFJ56anhbLJMp7KCiKEOjLzk2ivYXFaJ
v+4cbw0y7swcafuUtLFlFKNe6FhzmjlDUOTkD5JoJ1HSa+auBB6GTe5N3F/qfP1TUYvnIdWrwK4S
lq/1xJjdIXQXYiPasVmj6vnxNDPTfU9cMKrM2oFXf/raIm0CsgWDwVal+CstdxZEMztv4CL/3+po
p5NXsVFrZ9nvAD4l45ssPv6dzHPSaTIYssSA8p9LqmXkyQCKEnJ0gzGZMjmeg88T3hBqF/GSm6K6
CrLnRWaPd4qkWnSgnt3fWuKmHrK+gmOvDuJdFZ/GdNACy1UcZ2SpX7y/g8VpVQVROaBy0Y+BcE5J
yG2r0ZO2uPTUoITtjSU+HuZrNKARbcEdt4raDq0p4QZfB0Cb378I4ZQnLQA2KoDgaOviBDEZqEoR
I9Ma4hdKl7/Q6ynmRVqcXjzdIn056n8es4CrxlRr+2I5dI9uMNP76zkguOCS+KfeiO8FIHTRdfGH
PYesuZ4sTuLwCxd/gB0hRaJt7uAiAvE75VTylxo9haNvOrodbVNseshmJgZd5HsaTK4uKy0ZCfwE
0sY5fRYOllQTYMf4a1cXdDCXMBBp8Ag6xlczDBy3wzPkzfbOy8oohd2rIVYo2v7RV1nu9XfwbR+x
4d2VV6Qv5kW8Z5JpHZUFCygdEuthsTU8H5fMfK9M2F197I4ThulS8LWhXjBvIK1p21JA8Jjz4qFx
yCc/y02uSbKgjlZAZJOv7EyGZFwszg3E4wBPghtJerUPGhpBxE1EacW2ntnU+ES+HWdyFNcvDR5X
Hs7xyZglgi+UsjDrJjYNAFzJ5kH8YdsWBdCwOOGWbuALC5/4Jvq5yEZaekpVZxxCNOwVHi5c/R9E
yE4VX19wNQ3zulrPTmpFuhyWJY+Famnj1aBpad7qitQ3CSdeRyXLodDhXInu/gwdqd3v5rBp3yUZ
OtqyPo2t5KThpSW6yTXOtkFym66+85UvOi1hx8pOeh+cMlVwWxbwDoaYY39ypNU6GEUS4D7Zg+lP
37BXTzdtOArutCVT4D4n5rbFcSq+CE9oR4nx+1dSNGAcbLVv+Ydo/7bW8doFqAio1olpokNN0On2
I8wTphdPIxrinNfbO+AAJPzQJ/nYqKaOdCoTQwWhjPpFxGqUEc2iGatMEPMygQQKZ7L89maPImai
KFvifZT3176gFgBGFfJiP2DIAZLFVUlHM/NqUlvNbwJnlglHxjA01Q4gGLDjf9iKHFN9T6ylVMZI
Uk0QjCtfL/R1aGVxZs1eGudiJeqlITb7Kgc4AfZv4vy8QMxd+e7hd+Foj4n+Rs2bZdnChOndxRjy
XmkQOqIH8G1pXSSJ/RdM0YWkPGPEcai4Kg7p7APmUxhVZ2X4zWrVeJdo5Li9NnBoYtH9mrPI605J
Bga9KVKIpp/0uuWCE108i/glIdHKnDd2gja5FNK3fuQ2zrC0AcSNaOUp14zPjBuS7/j1h50Cn5g+
sYZLw1W9AZ6nD/6s4VxLeIOxXytoDx78bDVtaDQjZLZgEpStZCyau750KyNh9RQRZbloLLqKJb95
phY8xtcFLpRzQOKq8swVB4FyrJIWtk4AK554eb23/lry7Hs2n4Eqf8V5xJxAOopHoBValRBG5v/I
iKIAM63/gfG2uiH32hdaaEU76HGBiwg1bhaHnDRN//LwgjL3KeZkDxSdPYHf0QgVASwD4fgT/Flo
4RqwBRxBDDmzbl83rQVta/WhJAlNfcx9UELn7uot0OUD1Vdqn8Fg8lv3OetJ8vzzDn/Cp23oHOLJ
XPkoZLZ0AYWnJUTw4vUfzRhNUCzjc6apMTYYES9+cHfxmZrnJIutxxVB1Dmjo6DxyWto9A8YPVhO
QohjrzAyrbOftFJFtJAWKksLDdWqayfYGNz5Qj/GHlESg73iN5cjWkBKgzGFIlLD/lwMLvTckWNq
a0YI5HiVQhD66nCTs4A9qqdpxzYwAmDQAftJkBCzcXWNufw961+bUH7FYly3J57aQ9329bsiV2Dt
nybe1ljZJpHsZ9oWUlstHarzwSWkDx3kpUHgvoWCVKjxipW0pZT7xqbVtmZ8juoEuwn5IAayebkX
7nDMqxo8dO3d5mB6ggjeKoU9V3bA9Xb9BADw0YH0hPZciP0IyTDWAawtOE8UlRjopDFle+iVhlrA
cjXJI4fYuvqBf+UIBNNQXTzCrAhAEqOh8MUGpfcyYdhhI7NVNAKQXzyh7AGdXg8w0ObI47STbuj7
4WzMkt+dYkHAincafCCqEOC04f7eby8/3RRBlfoxEMrJV+DhcNrzR8wDCYzKnAQjUfG8VBdRJ83w
JQgqZJDLabky1J8eDjQ9L/ynfgejcnQDw2E5G0v/h4tSRlFXj+aExuV4B4SOz4cs6trvdhNSEtjA
/Y8KReHXn+w0kZJV7F9wdPO0XuVTk5OxfqEjUl4fnq3s7Nqm09yzGusnOTNcvnLrJX4VktgWo+cm
1RSwESOcfg2CL5GGwESyCuz2sEFe46ir2guoX4ZwmRbd93968RHRBs99qEh1Qnr8Q9wwL0I6HaT/
BIkSo64qmH4vxT6eCGNVIliu8zsAqzvgJTYMSr43Pba1/fSsY3On7bH16ztxatgNDMdNjb2S2Bci
7we/J9bkeXCB+CL4mVPVs/41Osg4lu6ffYw2GO/XPhhpxUEYQvfJyBMX6F5BquRYzRtkQ2z99qvJ
jPw6mrdk+MRJzDbJzFpPGBH02OaTj32gQ3W/NqRLtLziVIzMO1smTFKeKtQpfJ7MKYrYO+hB8PMT
+ucl+UFpKSyI68yxasHMIbjGd3t1F2YaRTBafEu7ULjTSPZreSPFfS7qYv6rznJOQXma5iUSQnUh
sf4n1WRKOJon5G5bSJhOyde9V2qyuqFBFMESbyMt9M16VbjJ80J7YXxrjhbdR54OG7gfrV1+j7Tv
QCanwZ40uz90Qln26nMZWsRULY8tXzLdP7nu8hGuw/8vUXz2z2v4RBNwTiDw9U8q1/v2u3GFo49X
bHMiyxbCaKS7yYP3xABUwbkBOVtVoUg18RJb8+NG2yIruMfy4Q7Mk9hn7lbYewqN+++qs/a2I+Is
K2I0AaqB2ApRTzWG3ohV9McGWkvXG0FcooCfJCVQTmx48bon5MvWtHpI6ul64zYwVpAbU61C4nEq
Z+J6r+mi/ZbsH9yS2p/I5KTL4SdTiZC8KBajDkjZNtwgJDv44U/Kkj+4hCTfNBegRsnVR77c3d7/
11vAU3Fn+1aVp6iIiDnYQdhDX57a2a2/f3WJNOlX8S7LrQa0oIgRt4LUq1ZGchYzf5x8OGANe1t4
ySbqRyDqAw0XbcveQXNP4xP6dOleph4ydMevt9Gi8otZP8Af88w9hodF2put73Vpupb7y2o0qy0Y
vs3rCE5TXdee3buOWbJw5y9YrgKotTO2M9AmnrYBC+CrfHVrj/dsFE403aMFoUINuiDq7TF7fKk6
5LIbficfM30sQXkZIRgQ18y+GZoLmTBOpQw4xUcRmWRbYcmkiJ5MpmuhEHaaLrouz1cQc63tbMyy
kq1Tpj7nXMBcTQSBDFWCUmoGmsa1p8sjVkjjmmWqSxwRhzPgwPONIW9H1BgUU0SSLLRJm1FyuCK8
m3tf4+1Ap3SST90Z9FULg9We2vetgwkNGaCYfqKQSvpCEyJAkPjB3HAu7X4CyUsxFc44UYCL3fXA
xgxhREQfE8MFL3IDlHWXaV0w+zCGVynUzKAS3pyOOYRRhk3Pvw7PQ+xPXiXffOSeivwNbB8E39p2
J1FudRlC+v5tcqz5gM+QQX+mEHHmp+AorjvTpjwLsDADW+/PQqDW+FdnmmFgOy3Ui5Vcbc1EJerV
WiJ1AnY1BBtXMYzVNIOj9DBgoADOZ8szd/bSHrX+hSOSmY/groHm7dJsCZFmZSAY1Sg3uRLsRvtq
8IyqOAxe1G4m3Db1bxMcYQHKDhghf4R1V+hOAnJ0mPiWDBWg6kpnxxw8D2qMYvOR9/q0k5+RMrBk
jbL0xlJ+SMrf35ri+bdCFyBx+ixOd3CJTQkG+FwfODaYO/lkLRQk0W48ut3kZkkPxi4X0tWhfnlY
hvAd+HTihXLTvPmkRTvDgDkVvm1n4qor3rIC69F9Z1CaSm2m/dwi8wI18KWT884wQZ+ULKd8AY39
5TGKConvShK43zYCPSAGrSeRpWkIPJ3RYX/ZS2dMAYRF6y2JmMjira956yCl/E4OW5otopd59qoy
oFoAB2/yVzZ1H+qrYKmblpBDGB9FtfNdAWBMQn3ojGcqWaneYtFoIkLaowAQBgbpkSXESlxIRJBC
FwbSoPo+aNog6zcmKMlUhLCXAmnPBzPiykJ/gRyPgaCLuN/F3f3CPs5Yz073cfVusTNewAwBGnPH
lqJsab/F+jT22SEzdZ+nka7LV0H33pedwprbSG77dUrL6SYosytfKamOA+r/luLp+UTd6/pjbpOc
OL9Bc9dYmSI8ZAuNxlc27TDclQffTv29vo43YV86kHAR3dHBBToBIEaIvuBPJz4hm37bcCL2S8DM
BVhR0OB05zSeM1z4ZENciBtXm5P11zXKMkxSMKOUmianjoI1mavW9woxdu19VxNbqlDwg/UbvYxM
6vecO/1jBFUnIAw/l8jC8JNKPa+o5PzpaxOw4YdgewxfhEQ3BUXhoMVGZMrOzHyXK6/nVoNzct3C
yt3YTVngHgiNvTkTwiKvGvhkPC5vm/iQs+77//7V0WaNPGgAPHAd8Glc2N5uWSgD1nxIPtCBMzU5
ErvSfQNfhImt0KffopLPW1v8D7syuC1PTaW99uWiPpbedf96OPgnWdoyx87r8xVEn2hr1pHlwqhD
ouiCO6yrqMlcIS8hGrVC4LQoJdDRm4J/mYT1AQCv7kgIb0vrkqYSBSAC+NRIKP3mviWGLtzSGrs4
GRG11IsLKRsPlcRfaYFIF0cv0XwpfRM08MKazCgittRFxWUEafVEK8ZSkAvbP4StiHnR69OySC4I
yXf8MSvzSPM4MuIjDT+H/c6IFuUrgEE9AnwkIfTD956LT0mrFgIZ9/9LVDy7hPU7tmfiBfb3oVzy
dT2QUlD220d7rARXog4DhUACCuPdscMjlRmVHYejZ6HoThaJM15K1EC8l86OCP8UMaUbk4IisIc8
sTwpPx+0I4iQo0ewRnRb1D8vEc7g93cLtTdBYhR6PJdsLnNnUz4ENNsCdOGj5twfNg17BwiQOQms
0HuyvoVFQ8aixxGfhtVizxfCPZWGMEfBICIvGDxdyf7uOIy50m9Ii0UTn0srY1dwIAk3+NDz2Kww
qXmMROZhUv2qSAOZsW8ytEOfB8anGv3PpPJgv4b5L5xeiAQEsa6scLV1dYBUzt9dvPw849jwhEnq
ilREcZ6Zh3iVU3tkiah2fKc5lusBx0uu8T0MXCeUR0Sn9kJBaAAXyQnycxm4bbYTUfaiOJlkYjIn
Z070jgjKISm+g1m2PbebysX+sGz3WGDMy/qUXL2X/quC9RMHqzE3gWjcGM3sN+hdQBtAqZYYhBkA
h77HV9yOZTvxCwPlWjiE5VxzcsqQGJ1kRl5rNHJJEyTT28ej0SSiZkc1wpZxz/ep8rBht6580u8h
zYWfS9C/6qPeogl/1LOgPj2Tro1YLUeN2amZbEOGJElZyI0wyeOb6gAI6hkbifcOFsIbbpEQqICm
zqgu4e7QV2YrIXxXCPumCfCCKt9Pr9wneXBGtKq7KIr7rn8f6Vi4tev7H9i0MAJj6z3Qwcwhvii5
siuObnNLMUtOKnqpJ12gfbYAdjEgnxSCpLlXf+x1eL/eCB4MazNg7+evvVYSm0Hh4dNpyMF0f9jM
9En57ouR4DRKnNDyjmEaZh3rhTewNt/ECeH0Xd8KEPeHnndjIrPDX92vmN9rwT8nftwQ1qEm9uNR
GtLdJ3KimZ7eMCve7QBIUUfIqaQENtUmkPUQcT5A5Atjb9LsCIlDsVKh3w31SRJgmy9v8qVIhnIQ
kJ1Gx81542WQ22mEV1E3D5vvudOjkznoe7q3B3QN9LFBCcyjJGRoBojtaz3MQBeM9Eet9lMu0RUp
BDl4macKtscCjeYyf2uLeRWvBLZqMIt0lbcp729WeSkFSYaR0hiB5mJrimc/6shylh0bNuiGL8Wd
zS+qlJX8Av6Cn68wxGXLGHs5uJ/Biy9V2USCCfb3gKk5B9lfLCzSJiQ2FbIEk1UEpe6I1DewBgLe
7lWwp5yXKY4h/OuZNwLiSz1Vklw8FOqZaCd0UVhSovWCJcsBGPRvSQaqYB7Kz8wbUrFfagwMoXpc
wRk5sqhVpX+u7Y8TQKNRaTXI94Uqkio0t3BNKbSAS0/MYB/f7QL/aTZChXsMEM5eT3D4Gv+9PfLg
3ghsWc7epF0Nnc3D+0frajJaHRUHF0tkJ0PH8LK9qtsIEvlxJ9KB30CpMLT/AQUb8ODSmxfoj2ou
KiAoOVnrP4JrvFyZpTs4HmrqUzQHaXSF8miwKrPAPu3cpM/MDuqusakEiw8a5JkCkucfGkMHeVbw
bLaK4DVujc7S9B8NsQdeY9fwfOfiju+ggLvK3L8m8/Uu45ZoxfqwC+XDbwLYVZS3ASWQLoejs6wL
99VGVGwNFt75sW68vfEkWYDytWx3qmen6qytX47Nk2YGsByfvki8m7nw90uQwz4rVIbyH7getdvW
tmPQlJKcBdpRijw1Op5vn7dHN9/yOrOE+6UzJSxH0uT8uJo4mgrMaBEApGWZI309DpZJ5ewGfWC4
tftLf+NNA+znmOsZUdD9zYdP00JPYoOy7XSzcldtRGuP9AJa5flW465usmkYKc+JO1eeRMhu+SBU
KimBfzjjLY/CqUIIQAQyGH/AkdbzIPG+Z5BWPFl2ZpvEYz6v6y5qJh7GqvYdrnTlQcYGwyihL/+n
eXg718hcNPpgPL5F6sVZEiOxswTG82l20z6LCsknorGsI8lVlQhMfDqq/GlWz48+fvYmMFcqfyFo
Xp9YokUYKv7nDCWjLICUW6VlOTLd02/4zEHRkjTzUSp0C7j+Q43qucS89JKKFQH9C70KXd6hNkjd
ddxYMaFZ8RYV5AZKaHaGnjzV6tH0TUXguPymLwRfxQzH3jV51aeDIEgbemJYxgRPtOo6PiwXVAf3
bHS+qXVioAC/kWQmLA7On3AJFh5kOYmDCBsj2DR5EPUvFiAdOOQyUvjzE6Vt0VcVfjBEpDHYMxc/
2ubzZ+Adn5oMoIZhqFLTAyvEWpcz1tnwLOie+9pYgAyEah8guo6BpGx2u3IWeFRDzmW67ID7/Lok
aAwGWkYtKLMMpM3PD8OHuPhGc1VqnRd50gjrqR1/RMvmZhrh6w0qvMdcSh9RyJMTMxxn1sOBKoHD
v7ukrrcS4xSTEKikcO86tVYT0gnaYnQJxvsZsLLW6zOaNF6agVmEGO9HoDtRJm3y0462OBYM6hIv
fL8cJOKuiM2DC593v4odHS4QIqNo3O0v6r0iQMpTWFSvieRtYBhttAPieS+g2ixcD/AlxYquNBZA
j3nio7o6dLkVOkRGOjhGglPB+p0IMd77jtkggZRfdnWB/IVnPSs/ClcF1U9UZN8EuCE3hPkRxpao
eD1Y66d9ozcOy3c6BNqF7m6yH4ijnnIVbTNsG/sMVmliiSjbuLPKRjXd7grFTDdZOwX6iK7FgUT/
tYF6Oc/J4tYOx8nLEx9N+5degy7jntQIqR/5rlCj+b7iEgizYiC02PF8QP0Vii+sJStD+zFv9pe5
/PucPXDg06YQTNWnQVb9F/1ZpmAATTmIwSf1XSifwxL7zuTWvdqxOaGVtWMbeoue9Yt99xKNOWUN
aUwWqO9MV+3EaNkm7h9rX7vecJcH2k7EdHiHtMzwNqQAapOaIOQGaKAs6C+mRhVesOXH5NqgMW7Y
F30sJX7m2tghRb5Z40PR6JWiU1L1y+ILIKNRcLs4bRBnUjS9XD5KhVoljYGKNfWiBDG+KZzZDcw9
IOSwPMmpKjoTytVoyNMxCx2aNUDUEC2h6LycPvHMafuU9AssFvoQ67tcl1+pr/rdM/esKwgsD6fd
ccJP4MIQd1zbGPDB+nJC7aCQysh6Y0Pvs/KhcJ64cjIWaGuvXPFWOuVGqr0wD4RVG6F9eUtLhNGh
nIj9fGyYpEbr+le+m8SiDBbCynvgYZObvwTqprbn1a0oBEHZadZb7AQkW7Uwc9Aq1AZ9zSSvA1fI
4U8VIs1khlYcD9/0Hb6wjygBxfqg6RJ31KMHi5pOvwk+qukZ9RSi9J4MjW/qYod5xOmkPUm1ZG2P
Vf9XNKaan9OIccM5OJB+9Xk/sl2zCLrTlAxES9CS8hUM3s5WI4l0JnsgY/yvp2zDLAJUFNo5W297
QB3H1O8QUeUw6CQZ5n2C+EkQdXXFI+OIByFVahdUsxxfhgl3W40fEwmxKbfdQW68uusG8rIF9D7U
ymej6DnOlqHHtoI4MbTv3T8IXNMI+gwA/xE/Q8O1q0uowfXd3iOWjovmPleLqPPm04qOUtldXko2
3KoVRZ4ipPnN7PdMNwAryTtmENJTvMOebzEGmGXqT+nvqo/ZIk8NPtJt9lFhnOARCns8cu0j9h4X
yrbAewP3zRUqEYcvmDUxP7ABwoZKkJ0nx3rqONG7Scx3iysd3/sDlTS/+Aa7P60VoUAF95idrz87
sErSfs0uZ24dbCAhz34/NHEa4gbirwPGsjvM3wHLsp9iGEJZBh6LYTxBm2KmFujgOS9cAByvkUss
T8dkmnEJgiF6jBzACnUd8JRkLwKda09tFiIHJlEQ0SilUJdUIchkBfVEtxdc9aJv2v+ku3TE5Eh+
4yqEoxqjCb+/iAxL3slteOaAjkkgjOVyhnk+UeyJKw2IjjIrwVjTxatW3rDXk89G3WC2IqytoEAL
8dm2CgXJl+pnP2g+yj5vkL2v1oP2NPakvJ+UylnXjfHWhBz2aocTWRhBNCIqefEzyPHwD13O999f
ZWS55BUzs7HbJK5PIO//n/X3mdLJHdl3vNI92/cDK6xyFdv5j3/M6gouFdFN9jLBp6gaH2QloBCL
86HLywiVOTOEN0gIQ+O8DRAtcL6urRey2bqLxVk+bZS8Q5avpHoIgpi3J5BIdGQL8puH+0H6PqaW
g3qBnyuDEoiYQpS1rQS05C34UiJpKyU1j+N9foGuYybdhBHKNEklbjsW49vUZYfAGbkGt3lsNJDy
ZIjn8sbzFt5YGD1fVvLMeOShVp6AiDoG6wB8+C4uwZGyEeJWLLQFWwx+HxlFBC7qpUKq2CvTHeqR
BgotNhLbVf8zOlWuiDT2xsIp1hG7LX1bN/E/pR3z/WxmXIVS2sqz8/Sp6a/OtggiNWfj3ziOO0xb
YDoQRGg8ePG6c1w+FGJuqeAN1Ty+PSmtfns8eeVZ8trygvzjwAFpkhvaRUHX/VZfavP08BKV3tHM
jW55jVMSnPGBoFxfiEFr0sglTUdv79pjJGSL5NAWA1nPYNxZJQJ6jkqO9hYs++Q28cs9QQxsIC+Q
agtXbPWtljGKE2RappjDa4qQjXBI5BMS2km6gks0K+ehsGkxxSOtN+Wl0hwiDVPTAhxXypuDXrNN
c5iuGIp6hnJsWnOyHqPfyzt9nJBtKvnO8RIDT8t9cuq2Wn8TsvTu8VFZ1vFzANoaJqHJMOK0GBSg
onElPNUcPPOAqjPwxkQLFlQw8T/o8inu9+s9AVdJNEp6/2HvRs3rEosiK8TYNtUuSAqROXqaqDeE
idozBGtERBn9K+xx+BHYMHd4/7kPFln0e01xBYMA0/RTxNjziUtG+UUtlG/RvpSs38l19gsRFEk7
1l0+bhRYvPp/VdZ/U/SNJu0ZAn8E88fWr2mdBd2eo0/qup23joMEAbzYK5q3ndCYiEva8p/ioVhb
lF+2EEGMT8ek9f7LW4NI9dPC6HCx3/lWgP7IAP0XqYcBJb9egFMS3BaeFM6308+kpwU+/mGe7Roq
z8cIG6wZv5z6eKxIoKKT7Pu2+H9PSweTjk0hg7ySYz7ODx+pHm5H7qLSWPuxvt/rJyCOPnsG5lYV
3n33LQKcWQWJa6wwHM+Dpbg9+I3CT62BbaOfIVPr+1UGkeGVDAeyoW96jnyPdCsvtYVtkfK08Hnx
iPlzT7Olvc+MEovgEaqXZYdSfy58dFgIkMUn2fDFFwje2XptfBSrDujN79u1FrKi3wxICIu//ZmN
l3LJGTR5B7mf6dHAncex80lPECSmWIuAieo94WYWEq0uuMGtiFkrG3RoZ1VrjlqQqwgiPcw/QUmV
5z3Mh5MTMGXHHVAAy4OpqOvquGnjgbA1QhB7DMcXgfg5PFPmkTSl0l1XReElmvstg2c3NouYR07s
XzLak+e9ikYrR/MNtqzbCCrjbzNL8UU5JpM2fOHC/mWBoZyy+l2yPiHkwwClpY74b714ViT89Haq
ih7wV4wn0z8AjPztrpwJw7EHPclatMNENrXW0PmjIZoyqzRFpwJQPh6TnlX55+hi8bvzEMe2MJCa
in+JfKNCKygA2OJ3p8zGNGWUQpeVph5eys8hmmaxZwDFTPIltDTBxltX/m3ObLR7tg5jaS8yDZWA
G6D+0wm/6xRMa4y1rcVYwqHuEgXCYxpwcx3JiSpvUwO5jygAtKyNtwkUZ+JoSJqhh8lHWflwtwi/
au+ow2hej7+TmbUiBta0d95FFZkxcsUvtAscV4G5a8Jj+MZSInKhjKgOI3t5J468UkQCqDddiqby
xjtWb/gX+H5WrCVJv7GcX15d7Uks/mph+L2mQwxjMtCl9odsuv8cbUZidzZBvVlNg5N5AvJDdgFi
Lzf9PLLoya5R3lOHAC6Rlc12zLqbtyIOpLK/pQFA64pq0HfWxmc0Yjtla5usHoqqLC1B/h4FAb4J
xSeEgVqDI+PlZjCmbuEcFCLsIS0I/am0wEWNRO81frQnE/hg6BD3tFapXuJ9sGCY1/R1Pgu/RDiV
Iy8r4CMxZILSLCs5GVMpX9Y8vctX0EXElBW7gjln5Drj/Q23nnB0np2O57WsjHy9lrkUjIUg0CNC
PgaCFvhJMlYw5jnl5mgkkQiEvkg9nj1F87Cgql/5ScL2Ii00zTYz7rP6Ef9XZAwERLyXEJ7k/sa+
8cTUim9dPrTeMHSYkTmkr2FMufYL1qisPCC/oVTy38zsjB0laeU9TFjGmdwYWA4ffE4Shl37qH13
qO6vx4I/uUe/iJOtUR1mkLCKv9u74T4cv3nwV+tPlntjYJDCISP1qvOs2mh2RVKSWNGpkVg19nFX
FdqlgYvl9FTjveXMKVFSW8HsM1Jdu5Rl4EgdcAZcwq47VY0io5lcr5XzsOCvEg8u8Yj3HOtsCoDr
iPoVOWbX+0T7HijMp4qnRysz0rZV9o/DTtJZ7UnpUk/3ZlKSoS92RaJhu/+JeXYdHOG6EWbTJOqX
DWF7YzbKQhZWJcwHnJHB5eNuGg/9BxGJ5c0p5TZb6Cm68eMzuvOMbBD5whVnY+Vn8hGK5pu4EIwn
odcHGLyD8EIl360WpjBo/N4c8NhsO+0a+3JXVHk/XBqRatIt1du1lAu7wLdyVNh0ctGnUai1hcfx
6DbE/JRiHgn/rCv1C82zxjtOOVsLq5ZFjdeF4O4k2pmnQW+QWXyoqbHT4SAMnbL4eySQvPiyHc14
AziNGB7/Z+SYTcHw8sl7Z6uNSuJx5gLf+ld/H1PUd9e7S2fNNdOf1GbYb0e0L58++xnzZJ4J/Y2N
FtnTdqJqNjgI+aR3u+0UPrTgRfW45yaNBQ2hPx8m7j6NBchSK/wiKd9FdXn8jLMNnL4KERED3aEP
0oBVUZge2RoXNbocz0rdJ/wGzSUdEw4/gEpCaXgJIhh0u4MFo79aj5OJ2Ew5NL08cMUJ80DC3ypy
eb8Z57zaUQQ1iTfFyNvic+lVAzIYpsgk79iNGP8pt8ymMgwJMrrWB6kMPzg2zrBbgit7CLgK2c0m
+/7aKm5S9scX6rxPaQlEY5LIewzSSnh+mvlGKpjnEGdmeW+NeJQCS2UquVcrq/jzp5UoFzBMMmo+
UbQtuRtv2Jviv8YcKk4LtLhVltZ3zcgFpUfbUQOU8BJYMrrzl6xcaIfKzdMUZ3/GJVsuzvcc4CaS
21qOHO3t8+pn44WQHRq75nn5Q3l7n0qjzi6znxZAgeCp1r6gVD02K3K+MXjWlFR5Uu7oDOsSPGg4
gvJ2pI+ELwpUC3crcG8hxgW+BP+JM2nSHn2OLsV12tZfWnVBrusVcY9KynzgctIYOp/aNRCQWgl2
fyjojZNlAbWWZFGLYFNkBgkYfKWT6XHeaYFLQwUoBGuKyoeSoTyn4PX0cqO1/+lYVIB/0AWeV9Gw
OceX1pNNAhTUofJ4CYp35kiVBdbcbtiXwkWorNUZ+ZJVdYXQ51LPLJC+5hobf9xNNprlhypLVjTQ
dUmM2tDOuxuVauso0ymPd9aELdSNqG6psSSRk4obbatBwq/H2thWTJUBpHRsdSe2IkRirWrqZGpd
wdPtm22cskbvsi0XD69yt5esrFfvrinVLAyH3jAeoIHdTzvzT+88a/J0P27iEzrOE011hRoLwfqA
wMCLIxoiD9iWrPIE/SCb56I5lCpjaZIl7IxD8jS9G6AXwnZEyDAl1KYGH0ily7N5V0t60oe0oCZD
NM+3+orRuWclWdlf3WZzaDEgWFuCHW5Xe+BgXPmk3TtS1Ciq6fJF3/K6+MZWL78vGF50gCVC8Iqo
naeXkKUllGgSiTxmZz2wz1jSLrKyBy0V9BISdofyaaftFMzDVETJ6GvgOjhv/8/k6KL30ohGIZuZ
o6M86XvgZmWsGBE9BLc5UgqLd4v4+hQgeVQ/9suGb2f3yfglqDmsCfHhBmegPrrC3iVCYqBxpJfG
taoloxtz2L+cTKmFEUC76aP2jFG6pWau2oXY45snz0V+7AuJs1uUacr8fw8cui0zwXmvFlolGAOr
IufKx/s/gETckbgors02QS2L4koQxJq0G762RabAE+29x6LIOy1RIlG/xYZ93X+QgML/15YVW50T
jjpWhZE6bdq/dnqpKSHpaWmWoyML1/nvbZlBqm930JaPmG3Kx6HiLZ1al+Dhv1IKroeVKAmGmO2Q
tpBxiJ0IwU26LkPLICJIxhtTN9EwMNtO8dPG/EIFWB8McxHQV5o5paL+MOlILwm5rJjHwcC3ESNV
A9rmGsMa2w3ukIJN66Gb5qPQYgrw+nI9uzG0iIwWfeG7eBV/ErYgNPgHN/jaY//83bfuoYZrIrvW
S976Q/6b9QsOY/uSlez+6HAnKt1EurOJzqfbJb1O3JRBJi4ke2LGvq9qDhKzXsO9dsYZHVuppVzV
CZShvP5qoUu32OiHGckjDpvzVSxU1gR5vboWcEc6o6N/E96ogxH8XixoHOE6zTQvP1AMYuaG8zQU
m388JnmrxBn8ss3khTB5Sqh7GrZC33iFSrZADTeKg7ytn5XdVQrbslxPC7M32vNwwkf+c7oHS7/0
kddJq6NNSWddsdIQYBfji2iqgzQFPYSdSfQvj6CAc9f9QN+sscw0cJ4YZ857id80ZqmLLPb2yynE
Yt2zOqnhJcZSNfr+CRdo/tAWiWDuMEHHhY5VkmW3SfaCDoKojXDwj0eL+G5VnorK5x6Ssrf4t6mU
1BuOJtXNmvkJXSul21cJlxbcA2eu71/RorN79JD/SnfTG8hGjTVWAZOuOyiBOXpmkdjAwgR9Y03e
xOphP04IsdqosCapHHkMKby/HAQL6cHytF9nyywanHa6ptiUkJq553GW4pu4G1G2yRWmKGJbBvs4
WWjUVlrYTpeWHA051v0uBevllJgL5tpTCs1YIfHy9fJs76bIRjERyLNpTgwW/IDlcbymX31nwqnK
eXOZg55xqcGfF6A0pMM9bjCzl4GTn+axMvrdEF9RusjOdQkKofKDtxXmY8FrgcE/HQ1uwYhp58hx
fa2hscShakSISz9CqMlqKdLpKGh76J2uRPzQL8DwQaW/aGkzH0rxZ1nU4vfxYggQSr7KTcvYo3LY
kpi0B6Ou4qGvEszRyjPbzDCEg27rPRP4HQts1jawhQgj5g9JoYzqhMM9S/SFg95BMvb9ncqzLXXj
r5RuvYSv/Bm+CW6ZNGgSFnV9L2y/Sv4a9srM0ETD1tNUCZtFP+TQrE+z4gKSVE6/vNZ1VPlq4MON
m79BvBAMMYkKvMFDe/nI/eKU2/MCUpnVGXaq/UfWraoCJ540ASx3x+O2GUrhSXGbwVLLpmiHN0ER
74xbSg6hbEf7K6NURDJ8hpBkIEMsLryfvoowd1eda2MfXNdvGFTDeL8jx3YvVURYF5y9yrKbLrzu
GqW0GCWLYWeb8Ua8fFi+6fX6Mehq/cEjENrUL0kjmGvCVK9wlhahSMgn8flQiYWu0kLubiHOYbEL
9mBxrmEssH0/AAyuw12coZr0xuBqyqM10NiNMz+v5DVa+4uOrhW6fk5fRnLkaWKbfPTUuf17zJ5Z
z8ySbpGjx6fB2Hs61pKqIOpP9WCCGYL2DVJJwmhCpH88qYLkEIiprnnjTQcBOYjOPV90viSgir36
SXKfZ9syYXKzaFTra1IzsR7xneKgk4gVeSL9XZmSTvWhUsLu9uuGTDBzWDFI06eYIUkdJv9PCMDr
rfO3XQeLGd/Gq0VQOPqjgdo9Hk4TAbTNKHvb/N3pFItRnZejRFq1ia/oRGOx9+eQ7kfoBflDKkCd
HJtQ48HkYD+xp6ZLtA3nKzfuq7jHQ97DT1G7/eEI1fSD1D10qeJnoe9s8HpEw9EaGw9+RcXqgPGU
BwuhoT3bnhE7kwwhLJuHlxS3cPdbeu3TkAAO/LJyM95nQj6GWJKWdpr5k+SwJRYOSfwrvAYZ2Q17
8IgCriul2ugvT4Q4Z6gxauoZ49ZNQHSESHbuNPuOz3K2XJ+2v2tu6SvARrN40pwpwHs6JU2VDuK4
XsZg9TB1O9U3d9BQQttWMEprAKN0pspiA0ajfShY/BZW3TNdMSLKA7vUABV+Js5PKVdSIHP704Sg
5J8CN0Cu1kZVe5UCyGF/zkUiwoqnzSdY3XjPNGtjIho5Db2+KeUG74GjXPCf1LZ/sd3DsDdbnRSe
/2s8bacRSaZPNrOKtq2k4UzRlIO1Gtb/zuuZcQyiwhfQVBzP1MjHSwr0/ahsgApdHGwG3SqaSY5g
QRySUiaFWuU3Whj9SwHQQBGJaqWFckPxRnrV+gzZikKF9+g1XhIr3fscNdENcHUUDpytT7Z9rKCN
JqxDVFl9+klFicq9daZcmYo9jZEZVfZLMJQFw4EiUs+Nve1oWJ97LUby+TbBkNN4ZwZV1SNftJXi
lf63QQAmRX6g6VFf/kutDX6wNJ7G5Cjkw2fNtvx+v9Fd6JuEZLQs9qy+ZdFVyCbDbvfl3BexWKrb
PLl39DJZX3iv4rCJNEbyzJZbl6VHNMO/MsthgxKgMPJ6saPUFqxVrT5HvXPzCviivwJnoMc5+RUQ
BXmqZELT2z8iMffx8xNUwVj33KMMgq6ROgSTFoCgp8L94zaDCg3HgdsmVUipMMaa1rRzPjBRH7ki
wF9YOItZotcK3FY3mIWcOeyr6AF8ABF+Il29wztB7uaFIuDPXcSIK+7D//AjMOxGH0p2nxREfp8Z
lBUZHCGddKvZkhCVI3MJ9MTZOrzhYZ2TPyx+EqUZzGlfK9ZSyr9xpfPWe16+ybHXWQQQvOnpNecp
daDix3+MzDgMXSbQYUTX8lSchPWXkTq9gFoKYarIlCO+lsfffW8KOoQGo7z9Spx6lwURuiYnQoIG
t2GSKcCiVrGWNAM+yYA/dPvSNvzX3oe2Z8SeKJA6kKwI0iSMVZLTdcA1Yu53Lyv1eytqKvNMYasD
fdCFetJt766eFpKzLMfL0PAeqSa2MG9C+mukXJbV24GjgZQJ0XsdLKSCJWTqUgkZ12q5zjqOxIba
DvkpJi+jItbucwVbJHdKILGqNfMHN3XXe5R9dwCTdaC0fnie3IUGosFK7LiOl+9iHCAUYEsm64V5
XhDt1AcxJWFbh1TgdMygMwoyDl5KKYO8mUYKzzvh/axj6PSQj+RcVj5uSJfAVq1NYNklhRV+Hm0j
WUMkSeMzmi7t8o/EcqgjyUVcT2mrOF2Z6LfxXIsfNAJM0hjYXYl3hI0XzO/Bzx51Rk/TisSPEK4o
uVo9o95B8rr8L0QObmmcgXg+ikThS6CdADstb0tRunlkyYUzuc3HhXhorUkMqA/exGd0bY1cqlhG
g6wmiTrm5HxqOUTZ73hdMlo7Qg7hUELDmdm+flSeG1nxXBkLbT3Cn2MQnXFVz1fHa0yAoRjF3/PO
qiYhlbasMZVGP+hYGe9rd5FYJONKyM0Owh8CUlcdrKzFy8o24y1isUugN7cvltuzjB2T16R5zurZ
79IaOzjDgVi7HD00blklJ4sGUekN26gQy8A0owsdg0mLm/enCPET4uB5booqumVg560eohTiETib
9At8hX9mA8BgC6d8K7taalN/dyGlRz3m9opNOt/aElrEgtKnRuN6x3ZMMZnOn2gk4vQFIZeinea5
1VJByGBU3rho7P0Bo/EES9ddAkvI00k25bH/sO/o9RE3xMZJNZYuJYAiMd2Cn4Uxu6Dd8EzK6Dk4
PCXcm2CchQcGYopyIoXJmFEEOY0Ohnz8ikLVlDbvueKQzU2fYrYB+reG1cwQRAs12s2L+JqwfWbP
VW5eXW4oYg0Zq6SVECcz/o4ee0oervS/0eYx3COOqYzSSLuMrF7SjS1yIqfo2NRlwFqLysRAzjhO
nGRf/KRB1AZsQZQL9rAaU0+k2WDEcaNvuEkqiHihZKeqPmM3L2N9wpI4u/qsTmCWYsOR8l4epbp/
uzQpKHYRY6IBr2guRCKDYhVMWwO9cK2S6c6S/DAggR5F1JOZxK4+0omRZaQQdlhWiccLphqtqOnW
U9HGPeX7x9aqdK6RWgTSGPTyHkaCveD1+7ByEhh3C+xG3hVHhILjR2VkbW4RyyelxvbmtInxQtHj
NObsVQObiPqz97Yfz/aFh4wDgw/fJTt5ZHXk8SC/u9P8vgRAWX+IcUV5pfaSk4rGB+E80t1aJLdG
UgcLpnFMV/aVK5SOgeRehSyM9iL2gjp/uILxlFqda7UBcugQpSwiKHIzoOwPtJ5AP4Pv0r356/yu
/nIrMDnqQpqno77Kn65OmsiuhJW+JruQzbdjuMHOnC/RnIA9SoxBlCdchi23jFGdvUcPTZJvJsqL
XGBG4SdRz1Br7hrDawxFRj17FcnUyF+CnDJCc5pAP9mthCNjgCl2WWbxSU86eo71MHLxsoBwPjM8
JCLNflGadJtIupKVj1DvoQaG9hVZCUfoZBCRes6Mu0MwvfEKaNBDGjimDHfVdQQeydLs3h7aQJRY
mLK3J8xmyBI8EeWLuqUJOC2owJ3iF3iAvKhdEai1RS5Wyzfx0wImUwWCLQUy6QSjYYko8y0c6Ibi
9KIMfKONWKLJNbJLlYmPnjGTZkyly4XY4UeISL3l6KlqAW9MSgd38vZGa4qz0zyhbQkDRRZBHeJ/
MvYbYh7wtqgKegV30lS64nnuGzdktCQLEDl5X43rm5SG3k65Iv/TTXkbF6L7p0QPwFRKhXdnjNur
DvtoNCnQv6ObZJoLYEeb69H15zLro6h0P5I7cag2zA0cXVoQXgAEukwqIQVyacyoV0r8DNOlzNci
3O4iyGNPyluDTRhsUeTY4ENMzubVATtj2I6mhkl2bvwyBHUvEI6s4E6XcH+KivtwjRLeXJ37emLB
u4T/0KEO62ReMClHzYJmP2Ml7pfmnyOyys1NWCblp1RZq73eCAsIB3nGY8NUzIRJ6NjJjbce7HmC
Z9IpMQqPwRhaz2K5FrR/5skH9b4N2YQFaD0j3V7jBTiJFRiU9lh4IE8FP7ru2+J5e9J+U58i5N04
LoIh1HsDBWFM1O5KSdyJWu270FpsFpZne6mlcWJdPphxbPZmUFEzlC7dmpPWEk7G/a8yvWOqYOAx
k9FP2r3M3RjVPB7Od09JkJrIRUX6VhbThU9Nhpnryjnj4ZSmLFBUyvi4JdXnFgP28v36HHg6J1mG
CTbe6DZUzBosxL7cumKJQ+t4CfxpAsDZ+z5+9deNzjXiyBoQDdXZp5zmREK6IJDsQvcwssrLCint
jM3vFpc/+0bYBiRcsk88rJABfMYsMGuP28ZfIm+Sok3gBhGVf/r/gNgy1OQZ+WzgIhrgKWizfqEa
YNAzJtt8qICCirTVOXtE2Ef48iFYH9GW0GZbtHBs0NEMlMW2ANGOcvEgOOr+xaZWXPtnebLaVCY0
EoaFaTG+yheDx6Tdepr7MkrAR6i5AIBgtArMeX8Yx1AFc7VUeUB1M+Qg1TTTuppSxWOfcsu+X4xk
S4FmB4zL+mi5oCKTIJh/TlyRS0FiKgqTuEdT0TvPSpgsK3Ct2egb3BvTeWxOrPEreJ2/vI72Od+J
+BwBXfJNTQKSblb0a1HkLihQC98A/q+HsdLlqHov17OVAGvje8/F7D80P9e3XwXTJq+JuCPChqUI
hKBhJE2qENzkc6coPYHh3z2tyEVHWrhgLLTO4l8f80lDwxdoRWCqUYQdFNw1r6c+3JVxmaVrvVJR
ClPlbgPQqv6nLjK/5VgS1V166QNKqXil9Ga9Dp/3t2uFPCxW0zZPqolwEdFUES1lUm9ksMM3Jv7p
P90sKJxqxoY6jtKPtVYXPXDawYUD+yvw2nRi6aMy/31pdWi0A/+qJhQDCVI2XT+OTvO67ByVZN4Z
zBrmZftz60kOsUlEzV0p+D1Ay8okHBg2Go6xCP7gIkJmzV1N2WJUQNONEmRJs6TgE4Utepd6KOlB
65+HavUmTt2FoU5nTDxDjQf4GOhXA/UkioUnCmzjUZ4ay/JilvJgqIDG5Y/2jce7S4pT0vgL252J
Zo3C7wfwzfj+1P5Bvt/n+hg9ZHwQuiInezboirqVcrh46XvkOCR34pRyk14wsZOyP0Z30dTyKbHc
SCBcX2T0r1WXYqvVXncTaKQcZazpJhxhgWujjBwspvkQuXJiiCBe6+Wr9BrxEeM0eaNQsuyAZrU0
+64jLtWHtv5W+ym61sJvvZx8n1se7u4pa/Nt6Uw/6EljzJ31gW410GxQ9qo9tQkm7kWsPu75zosz
+wSSdItDPe/jOCRmqQXlSN68YS6SSpcIEQEP/tQvAjt7V2X8Y6DLOvcl1CQPMJrqjda12zJfILoZ
+LUHx2BeMp60fWIFoJInZlJDt3h4s/Cz6SqGL6VPokoVZhw4ZYZcoYurglW/wmg+pP2CJAyo+659
kTFljSLFuBWOHNcFH4AGcyHkC6Q3OzqzS2T8/H32DgGuviEkGJfQAsezN+nKkgGcyiZcQjWBCIL4
114/y5S/iUZRlnJMYPUx2/I1Ml4dTJO7ftUBHfle71OCI7H+FNe0z7FEbbBVIFhPfhZ52xnhgbdB
b2dJPGlCeaMHV24Nj1sWO/uMSMPM9I18zhr7PPbdEfi0p4ipE8RRahatx+8MxiTWerHRTOFygxke
a+HAeMEOjhuntI09CR2M08lS+ze8Oxs74M+KIUCYtYGAolbyJQJM7crZoYZKgdQ/rPu3nYqDL/xs
pfVTh9VfVQDtaLvCVUEmgJhWtQ4BBEMf+pcLmn9dblUGiFF3z3HeobV6Df4QgscN6J28nxlpWy/Y
ZP/1P1UJJHLVPiOU0CSJgG9kMBuVCnSx+DL6kllvmdt4gZQ/Xd5Pa2weub54UFbVj/Hu0mkphOQ4
Hm0KLBNKsSSAH3uQwUND9XnXlUaO2fv3xNhGN/LE6QBC36LLPAyCxj3dLYkm/hZcGKbxQz3A668G
16HdZpO0RsHs57AovVvm0gssAwScswHaHshGo6S7FD4fH4qzKTs+s0qmUpP6yPHut38hiUhOHTQD
YB/dT9zIP2RFzQbCnXlFf2xbbAkUPtyF5ikfdYDnMSiKigUml8xZVhtRzSsE1/HCQwuiNkofIJUv
H5Yk1vD1OJOUPNA4Q86st43NXUqy3uMBK498HZrz3rdXEwLh7/N6XGGbUIMDlmTjJyQA2UpvSEQq
FGYeilJ7tX8irxbewVXj2jB5szHmd5AlpA0HLyWOKqg8lS4qmTaxOkD1HfDxk6oVz71myJ0ct2VS
lUKDCqyx6YF6iq4mJPcCSLVGaw+KoA7pGR+kLqnOz86aCvGJtPo7sDJtrEHpw7k+1BLg8MnV+Ecr
7QJdTssPTeQkWiY+3fimASGbrJbXpEjmf+WxxollV3OugLN47/hBzdpuUhuJX5AHx0sSCgVxVkSQ
ZUq1y+ukg1W9dZRWe4L+j1daAUD0znGJacgf+VHXg3gCiQatRQ70hjaMkS4aa8GhSS3ZRa+CXnI8
D2k5N+xSPRDjbNcR0YUH3WeaLOWYIWlx+/tsQJBwqJRCgEks1KEYXzjwQzNhpAX5WRZTI1/XoB9g
byFxkDbnrwnoaAfNcjYQpsUce5XX3yCjy2VAgmLpdWsudl8owS0/kaPbK1gYfFHSHnO2/EOcl8ue
Esf5nJCaLT2Sbqd7zhnbh0jHkPyx9A5cvDNxwvlcUB04t2RbzfZuzq5UnzhbByVujSnHBIq0Wa+d
cnBGcaDAEER/+Tlfbyv3fkof89NTbPGuIxnWtqT6gVWfB8cEPjBvHWgOhW72kn0BY86mxII9XnIu
/ek/m/uuGDw2bZ3Qpwfcp/H5K4gkBf8xkNA6jiIhAc3IdO92CYM5BUt8/UizhdmUBVOOLLQ7Qgbf
Y9Qff61SCwZ2viOGs0PVk+ANUE6+TjmZRgE0CbT5Eo7CcbZn/ItMgQbN/xgHR597AMXX8ze5dZ9r
GamHe4tXMNVhnsD9LZ07CTPIDwsNy+65lCfGgJ1/nccj/3/dGDpz/+uE8Pk39NyyIbnmzOSW5ezk
kSjs2G+wHP7RcHhhTjECWgpYonaLLnJRayDCPeSqqbqmD2g0GV9cJF79TVVKWJS3Z4SuKaEhYsLD
jRO5XbW1vmrvNSqGPYnXwvgb5VxIYzEzjrTwzDIHsdEg5Cg506iy+dI8jFgJ6srTBTVyhMxtRrAs
F5e0zLKSCPUEjGNsAPppo1WClWMslo18glfW+K5go8GAqEbW8A1eTOACBvorldyXD5cFOKKbsUDS
wTEGp9omAS1LihnKABMxg0AKAu70ZGXv4EOfSmZGeZVKQGhOMZHAHB8Ve0ooMzxyvlE/+fGUnyOk
Bsvb4GamFXEi6bZFAPoIT86EfLxMZyJDSk8lH1BStMqtzQc/+8KiQyV7A7ShipobtiPEqwb/qeem
mFtvmB2/LvoVwR8G6ihP98YyzLjDkgt5GkP8UpCv4yb4IpEmR2pH3GnZbCtkljNww1fzewNHBygN
SHl5Vd6ZGOlG64HdZBAGKjaxeYAsNDXRuYHdxi0YKhISJpDs0QsJRe1nFd4Wn+JKbsaPFPT8PC6B
5DOjXAnaBCQyXQWBuKkQz03aC6dKhvWOFwJL6lmR1sEJ6UpkPsdMbn9cddYmor5TNTPylH8UWLaJ
Mq8J1++4krpMsbeeggjbdNiePX0XRaxJ1CAW91KrNa24iHCKheX2VbEstkJHISYfzPzmbtOuAkSB
nlBUfUJHOlqWtv41jmygRAstX/Jz+6jAbSVP/lG7L0GawsJUYftJHtjIZ5frNZC3urv6KYwU7OXE
zfSYUNSPMpFZcjHcNK0jMERET1PD02TosaQRunZHM8Ux54p+qa0LRTWm9zlpi18J/mshGkCqmHhd
S8hRS69/kerAwrunXeMvdeUkffhVh4rkGpmgEQQNe82ovQFaXVfm1MLUdgM4RGs6zfwnU+Vg6fSt
GIsChW6xotKodBSNLnFiWgOG0vqeN/uOMBVa4CbNwmbSka6P7u8vGIp7naWvbjTCCUxavIkIw5MT
hE582Hx/bjNBLtB0LiAF3DibTn5QJDiXssf2a1JiW1/i0iThpeiYR8kBidOIw2CrKjaQB2tPd4aZ
+UDzGLjbDDDXFfCZcsPBRn/vGPFhecKdQtO1FPdkchI/TuyFW/Fxt0AoAUxAtItWOWhJ7gkzfZ2I
TsxarrjmAZqEYS6IZGfMuD0vLoboDkIKkx43AdW+beaonupobDSy9Fz/R4YjafPe6J9loi4+26Og
pZ5BjJOlaXqmVq6MUl18gy3H7lGJe0KlkGWdg360sxM/F6hCk+8Bs6i4fc41JwAzL0+aVCgUrJf0
J8nKtrEAhVhdH5yW5UclY2mqre2bAK+WOFUHJluxd6LrLkzRMuMO6S0C1CHK8xRp8C4PZCbPO0He
9woEVd9L1e8RaQq1KMvw/0529Qq4BA7Igqa+gUtH7hDQU0KqPwSzADlATg+OKncnKnZA9D7He2QC
xmjZWHMoI+i6thqUcMGs/vDWPUnM1WDyx3SNruGSDwBq0zAtmyx6UtwAJ4RzZVsItbK5a9tJUck9
GMfmI8y9uJlRKESBSpE32c7oTwJkTFa69ynvnIfLODhkgVmgqpMNnBlsV2NLbFYIwqtSpf/M3S4T
hIE2vhpQh4ke5xDMb3VBSzBZny8+VQKBcTrLfFiQjXdRxUtwd2EvB0EqXp6HfpGB2icF7x6wq4Is
u5dBWtBMsfQMNFkoDCLEudRYSBzBW4F4rwjGU9J4B/5SQuS+HMnq+LMm7x14rFf1PKQLqdoLRYjP
lX5ubS54rN3jflhYGyD+YoPC1mL6ilZdxe1dgEb4qYHJIwkzgsw9b5/sHka61aNxUbFAB9p4cOjP
7VFDtEYEvmT1BXVtx9wxy9CXl41RiRP6Co1yO5WaAgGnz+piOhDZH9l8o4vgpGyEse3VUqSNHffb
kyEk9RcYB5KHJ4BmRe2gdifBsO8kS68d7uVP7ORR0eSLNGl3QZK6fKVtV5BE3RU/u/EKnqjz7Bca
Gbm9hbd5Yabw/QlBxF2XU4IPxVjXpj2QzcHdm8PWSmy1r2H/ene1MCwHj/AQPL3uVvUma51mKpDQ
d70qho0cF4jI9TRfhiN6w3nSEGaQtpaaV5bXqcsUK523i1RuTQYPSYfVtaUJYE7kKoz5yMzCIFMP
3nKDkc7D1sqL/XmUVuzYLOFSnHIajtRv0BMEr5+pihM0A2X6AuqFrTmEIQUG5IdmL0bM5wNJA08x
WAwL4PAlV4XXmePsa9koDJ3uSs0A7WkROtTbOgbn3hHN/IRALpjRGwZOyYvqVl6b2HKGQyHFs6Wh
/P8+8nNfJlaj22M06wOhs6FRybhRRBQEibc33z4oqZ55I+LQlbvFZQ/W/xSBiep6HLHHFgd+zRx+
zh1wp4uk/uJWzKD4WFCrg9J/HVsO+DzeEbJ1k2g1iHFdXZBbbZ/Kbh4KBr5rcw9kCGZMuUkItnCA
wxRHChjZ1guUugnSuOD9nEmloJm4VzXmbsj54rQ9z+JAVFLp6tc13tWaJ0M6OhRojvXkmKkT/k6I
igVI+JoA4CRMTPStXgrP+Ca1ttUAzEkxIx8+mZCfhkYAY5aUqO+tfejEAq39CRoeeLp1g9gEKI0x
ssYcGtsItask/dV8uZjIU/pWyqFMQCqT+vLapzbYBD+OVD9ggTxH3GMV+btBvc//96pwtvjCWS7S
hik2tf3rtfv3NF7UyrMNrIlLPf+9EMwsWgy1xwsjS41seyyFlBVjkYTL9htQjWwLB38lMD5kUAvl
bTTYOdUbaBTdSCS7HDQGPuuHAWynE3am62Ye5+yU4xteIh/4aK8vBVmByXlVSab8XUfDDBuby2tc
uqsJUCcGIvd+mB3xpVheQ3Oncsn2Fz/NRC92E7sQI3prLPOS+hflE9mpXR77Ki6OzPscXy1oldOJ
cKwQdJwqwVc0BxGbCJGo0OGUIDrjebbcR9s5FMuuLIGOMxNuCz1G02uLXiuzlRkHN2Gn1lTh2x/p
+ekRvrcCSwhFcih0kaBWQRobC3cVXwzN22z91yJNvRs7proy/RzQzlPOKPwli44Z+jWpHH2QtdND
TYp9VfXccMJ3RSJYKzMw+q3A5ZqYF6LL/wEXG8rzuR8Bw5evhml5oxeO4wNebtlOqmLHt0K3LfTJ
s4Bw2RIka6Akww6NIszNNcOkG/CGUEuMqxaGAmyRbnEXJYR3+5DhxNRPOZyMMF2zA9qf738q9X20
DMqHufiR2KOSQ98GLNdFJ1JjVpgywTya34TbKLiDNOow/jYqiazTiy+aQk4SSOT7P2lxZo0zh29/
C0e/8PppkPeQyhhq+3v5nsDxkXCQl5V4vxyZ6K++2CfsBV9nhF+mUpCGLDS7vBx5EkrXh/haxoDN
rMOPRbzddT0+sJQ6/VfrUVhnAR8+VbEAgC6tjwKPaSqlLtZitNqqSnqTV35jG++wtl8zoOCEB9tJ
uM7qOvxqGh7qtICS36aTFju5pinp+O7/oaPd4H8XeKplf+5no4uL56ppM8b3SRz1XjW8vQviOuoT
0IIeC0hNqM9bq0BXnp1aQe+2z3ZdX+JaCCOai2ypPiVwmauJUfa8IKAWO9IBU9njEEUoojr5EZby
mFGYBow4ScAqlvGL6QmuqJJl6DTJuUGoLlgrp5nfOkwngfZTVGnxVPWjq3KzxCu0UXUTYBLVgD/m
5cFJdGspYqsWGUWhBXy5vcxFQRVD+KDYBZKQTJZ5yTxDM/gvYv1nf0yYe7VwmrYlRsD23sKi3Nzm
f441gqYTZfQCF6rYQsDsaUEufjLmZx1rNO5Vq1WV0lREmM8SnaG/3o+sZrsZ+jTvnD2Rpu4O5OKI
O0F/NUDqkJTikmOS4/+ZIqNfnCmuTgsxMPnSj5iT6eWrH0ii0Ba+gkxJmsgnWGc7ZOgO815h1B9G
6uBC63zGfiBR0pbdfOOlc9FGA30ZKrmwxPrFm1onjNXWmIm6JHd3BqwZ1AwI92b1/PhZEqnoknyj
IXmMMANS1GDkhnSCJ94RspQAefLR27jp5AEydx1/fyfoTDrdXtJkzfoAi9p7cAnPXrUqiVGLDVTy
86F2sibx1PrNW1zj2K1IoGeBiB6F2oLmu1HFhUckoK7h1ngEabrt2aydKN8qwI5laz4Qaq+uYD1b
vX6AB6kjDYrTcEzjMYzOvoGgzJSMHcrlztxH5FpyQnicr21lHaZFiIVOFTA6P35ufWJDmcs4iWB9
EgqK2je5VIyLid2xISvmShM0OlWU4oXLURY20bKUXhKO8wFWQRtn2hihy151Apo/zAVLwwVQY+FK
KjcazZpzGIQ/Apfevedw7YU8Kp2gh/qNxIGwQzLDyfi4lTRsDiJkMOHiO71gQyCG/ltubypG0De2
jRgwQUmQ6Sgd5C2WvjUvnyXTAaFkLriDq0/VDVMj4Ngc5qMCbArZbJ0NdiJHeGk0o62EQcx36u70
D07IgkfNnVr2cTgBOqnioogE1OS3GMuNM5lZMzRRFPTP7EX9kQVKjR+LTUXdTPZYgEJiBPslszuT
DwXeAC1NWT5pb8fg+w831RUjYurM1/Xry+F5770BQ1Y+tsf/gms744cGEdRhuafqwYvpzL4y46Np
ZeHaxN9AOYi+bYuwOFsfSIdvmnbK7wzDKe9ByyOhqUhIi6kr7cDkSCwUv7VrjWd7GZzqPh5HBlxc
tWpIOcOCnmgQAVqPkJbxhJfbxEW/HW07FeRIGn9LbmpmqhZE0pDjOJXjwQROv4aZJp85W8jkPmBI
PlyuCqqW12vfzClLcRwQyFI72Pa9jhNzyWuOj6GSB+/0x5mdXxZI4nNPK4bdl1Xz6La8fNWm7751
7ABx2k+Oav4u/26pV43vLPTwnGLEN83aSzgPNN1nNqvalPeEwwa3ceCrp5uptkO8xSSWE3J9wtCM
zl+9sI41P4YeFc5fnp+2UILgJON8YDaKmKw2KB0paLrBsmBRRwujFS1mKXiQoDGR7Vtn2U6tQ9lA
FxAH2i2aQX77hEG32THVjNpVsvhNiznDJYKg3JUHpXQYLpzbQUec5YJexKr/RneSnwkqJUSQFgvs
EChGNtgWvrMWQlRAUOg0bOoQmXFpiuCkR+DHcMw64YhpdVTLLrOQsuY4bEb0ck+Ck6oL1lSClGGO
0vPAU3eNjpABKXs/mzStpW5EzuQ+6ROWE9sUiBXn6x5r7K/Psf4gN52gkCx4cevBQHLEApoP5yb9
4yDSrqF5se05e+zCmJlC8QmdJNTKJoRKERAIY0qkt9sXbULsq9zEHyEYBaSeq+LMotKfNlXnYAMt
J5hZEUTBZCHK3qci724Dy1pRSfnLyJQJBgI0YBJY8Wd5h4DTWVIJLneNor21zU/31yMjofqkw/WV
Rx1rVAeTCDAU+eW1Zi7PCE0MXLi6RkqJDSb9BT4iKrWnyN5FASxNxirrQlzcU0w6NKjLVnwm4JTq
PqJn37VUR6T5M8G68MOt+wdoU2REgvXgVI5VWYh5C+DWB4EFTUBKJqr4+ePthSjI8gMUd6+75MwN
aZnPOL0O2eQxLvFkL7TKdwGzPt8Pq8SgUpnkDvbZXf5MuWgEk2O5aK4SA8o9kwWyRycQImAyvs/S
UkeH7hPCo3ZrJr5Gq6gEh93ME4iZQuiI78yxkI2cKimnb0HmKbyH8PTW13QKgr1DjcCFf5c8LGA0
F4VkIXqw7wQLJXril9DYSM269stc5wshAamf6yk72OCwBnVaZAFzFzFB9nmAD/R4ncf7Gyp2rjpF
5zlTYq+IvWcSJ9Um5dnn78uMBw9HxAc6ChmajtBkFcAEvmJSjNzVIWC6TbSYG7ydRN2tYRBQSIHL
ZQAe5BgdbLNrorpuhqSlpekFnxmjjWtvFQsojCee+VkFLH4/4C7Th7txuGryrSczDoowOQAuvK2N
J9o5y3F0O/PHE/DGaYwEvcogktNE696bKpUFPL1rIo0nVnU9PtJRsW2qVp6G9rjHVo4EgpoTndRf
vyG4otRBiGjhh9wdkCbF2aVjAHdLBfSx/RRLt0SDNWpC1Gf4jFwBgdb/BUHEy7qCVClC/WFyKVQU
iE17jfAYzVPU3+5ZKr8idIonDl8Z5ZHkM5EDrXH25EB6DTc4/huICQq+g7IUpBnyffZYpwMecvGN
H9D1WugolOJy85NnndvqzAgVsyJpV2adCnjipr4vHHCF7M7M0bmLWRTDrmVmP2X+dfvsyu+47wS3
2m2mcirukJ3/9OxJK2VXiaED5VVHO5n39EHA3i0sOzc++XaqmOOLX8E25Xrfi0O9J1gh0JvG55vj
ms3DC557+WfHDNEXGBmfRIDXEGQFIPw9MdJuQFEpoBjAeWS85qH1gpJuWiY9VG0NfiPfc+f6MLwq
DCzNihmHJgWJ9DHF4fNTgtUIA6GbElpicyYnYf3mTxeXRrwXco6QAD++F93W7adJxMJOZ4QZo2jc
IMDArQhu2KyiOzEcQEdcjkXe/wijWh5RwgmzFRHk1VTlR0rty+MlbaOwz3P9/5mFdo5YQSCT4Vjx
LYwxpht2hy+g4ggydkdH0D3x2qwwf8Q7k4li45TqLkLtshLv6vQ7cei+f2TWWjPNUBormDXrO4ig
T0sOPSruUE+L9VghHcLMUdE8X2IBQo+SAT6MviyhVkwMRtPwS4lMRcCGmu3tq2lI9nNuni+rzuTb
Fi7yaZngiXishrGPjHgswpjt/56Ik+te6nLA2YPWwmwnxa0nV1AwJVZaLEtv2TT6VrfUDmdnQVon
6FoaayBilD0VL/JskWENMoCp7kbZZ7nu/t9izW6SITP/lOO4XQI3P7MdxfNuZrIfEY42gZNO4+Qi
pILBgJFvI2U9/JjuaR/+qKOUZ4ZqHjh30fAJ2PX76LNEdQjNZNd8C6iiVGIHs4AeaX7qtQoL/E6q
ninDGiPKrCyZn8AVRz7UWUgF+gi5v89V/EhJQxykgH755y0cPpSLfgiqWGSjJ/2PmP6RA+7Gdkdm
2i9FoG7ncBNuc8YZCucH0oFF5CM0X0Ek4MzN66ZjmSfbXfTk98CXkKzf1bRKqmGBxsAgQanqWr1F
x9rYVZk88hTpn8sel5aFw1UkVVt3NQawdnociJSelmQPkvJJoLV7dSV/AcjYPJcoQyjNZDRDcudz
Rpd/oK8XLgkhmHOuzKFNZIB8K4z1bwzkhIebfF9IT3QlkH0KEI6LThYYBErl/eXIj9rH+CYAda5w
9GDL4mIvKYPxXEbYtaQLnIKm+cpQ8K6lQzG8otWxLw1PXvwk/ZcEbgggglF1pjU1h9sxclnaQlPx
c+dvHjvttqjXjd9dNRm87Gppsl0MyfkJMx7dmEbfOEpoqb1D8mZWh3dpqiLExEkw60tfKOagKiO/
C1GEZvjq9650PlsF4loxfTJaMf1FTejUj/lIP38N2uL8UGOFa60FAE8OJs3+5H1oVJkN82/RMXT9
c3X9pHyiyy2WNeMsZwWaoNTAKQZ+DI71OO7k3fhI4uWpMX5eQKgS6QAAEJ5B0iorBQo+W8NXCya1
qx03k68YRzM/N7Tj+R3K9qsB3jv6ODdrIhHVCMI6lw43G7wLsN1ygeE0vUftp6KZs0qC+Sw7OiCS
bEvT3ky5esfHHfU6R519avBP4oBIkQU15RNudvST4IDixoLk3+1M5MEi932v+BR5qJBKyeT4Qtzp
zVJDueHqswNk76PMe8prA+wvBeeG5Lc88U5nQJf5Of4Xl5biKnmXGn7KyLlovzvRmUj0AWtb6bdo
FpMuE7ZJnHNX+btfgbqsf+s4G/S4RFQD5yfBH6YbndIvOPhhqfvedMsoh9rSUheMSAryRd6lcDFU
QENImUyES4LgopB/8ulxw7vQSgDryLe+jvAoLNFAsKBRnB+CiI8roPt4EF2myD/Wjds4o9ZJ/e7G
edFUbLU1RoMesL6p+5Vl9YMk/n51N6as15nxnxbGKEICPgFZuXpuDAHmnqgZfLVy1mBIWg15MoMP
psO4+BRNf/8vyaBFCOhg7JmgV2IOrsJO9lPCnBe/Bx2Rc7H7/+bTAa0diBPzJM7WfK+9xiahmNnG
jsu8tRzV40IGqRSytCW+45exboSOiyIZBInUwhZJbW1HTD7yCrEMgmlfnCWMXrLFQ7NExZDpTdml
FKa1JgbFnv3173cGh4w5CATtTN4mepnLZiYfbGaiWu4+aoNrd8GQkhx62JLeJ6voHb1+vKbS25PH
+gmMLu7ONkxz98tt2liYiXBzNP6J4AdHG52dVU7+kmMUfsiYyoJPw6Qbvsrio7LQ6AOLL2dOnPzz
mRZIBHXylJKAYqU5peyLZSbfg/5r5Jxdw/VsSqrvre0itjz+cPVREGnuasL+UGETUag1vXvw7tqo
7sndO4Mh5RDVG9aUrfx6WplNJjaNFA/oNdJgrb6ZtEqHtyE7QXlNFfo9BtdNohKZBEH61PWaLC3e
ZeY2PHbl31XsXr4+YpAiOKWJBNCh1E8PndemGPqOPVsXuVDbeizWsiJ106gHB0Qh4gHrMTJCICUa
DhDffZn7jqpW/JC7dr1XskKFdy65KCuxHbgr+tZGlLZV3dVKqaEBMjZ+M+pt+qkc8uTzSVBVqQNf
MyxjrIQULq8kbTqn7uLAKR2bCHU87K95xH5hV6hheCYOZ6SiIfL0U8EFl8WcXK7/6whToHZXmxyp
7JODoojBlUo0FavlvJQcaR166XLVCSyyjmuTPLMeDZawqqaT+u6s0Nt0wHvK0pRKvMk7iW8a8dF0
xLQEg0W23zkMNcFFkFxKjXJrbhgI1oDeoTiAT2NPPbwLLWSKx1gnJWUFdAq+5ylYtvxE7gc7a/63
l4IjXPPSiXb014WU5btKkAYEByrKnfRqUdP/U90vbQvAnXTFhCFawrWYlmNq0LTLIWwfGP/Kw+ii
hVkiWtb8M31ZWST/Q8NZ5mIG92Hc0jfJjufqChhE8SZ9z44iK8GrsH5I1kNqt05NppwjLhJJ9Pi9
yJ0q5WECbE2252RSHoSU2Q67IyaRzmLaDk0vwVF2cZP7anCavm9s5vPaAgP8djV1xG/Gw+pR0LZb
oRgocBe0+h/qRQiJpO9h0jfAWSeMLy4+lwH3kCymf5Nnb31dBc1YHR+LK3E1StG+Iq9CA1pzMktY
d7fxihvhy9WL6swdhMXcb2KlZ/pOlGn7ymjSCPgt79X/uQ714Qmw6XNhNf+BSZniumVuQyymdKpM
qWYBIK4yw1Wh5TqP2t0b/pU0AwlZ6vLrKA6uOHwDmUFotW9UjFMejvgvJVQNkrpjTk6lzTzoJOTL
taAzOG7qSiCFTQl7b5OJwQvwFAZQUWYqQl88PcxPboi/K9Ek8E6FiAnn52XK6nixgXPh5zOR/NPK
yHOBP63sInpvcBAGHCoiCgcAC0J6To+dgbeE3Zccow4iUi6rgSBxu0C4X8aruOLK7p/PCC2a7n2v
sgGY9y6wjD50QJUbxK53C9rYgn6JvuYzeTLfF+2KdAK/iMRRbzU2+ACBkZzQNfoyuqSbgVTaQro5
PQWyHw1xY+BG3spRhSPRlA1LlW5pu52WoUqaJzrQ6D5a5vu3ARr+buH/9ixTHmL5un9UIAhFonGm
Tvdtdc1znY2mE+xgHKHe2TCY0cOQ+dJCJtTR2kNQIYDt22uI7vAFw7UegFo1FtsZLIM2ifcQJsVc
sqhfO9PgINKIN/1CwRbD0cDh2XgdOhY/QQlNz5d5dlFMybInfDo5ycHgEZDJZa3eCe6gAibyfM1E
hXkDy12nW78qcf0LpxXbFJ6DD4tujIEY2OIMA9jO+k/uPYeS+8Qsycykob4rrciwRmnFbaRLgxj9
JOKTNrMhgvqhbprhmI4sKasKoLjyOBHAcnskBwlblz3Ob5Yf+EnhDO5L+265SAWVw6C5Cgto4XUv
v7yFbxcWR0crXVxz9dX3lg0pn/9oa/a4SmExA6640QeNplPe6n7pa/CxuzXWNeTu2V31jwx/K4g5
uoyu4f1CtjXGLCzlemIcBSqALHxKs6sKvotsUL4GSspoXtZcYNY1qDAaiBDJlG51DLQl+1Jmm2I3
kYbHtn23/T2OavLW3Le+M2ccJGBqVQn0oV3RukuRNvvSRJoCuNr5dCywoEyqYYuLzOMqfCZvG7l9
sVwcsTGILZSjV3/+RfDRBdgy95H9bl4OiDXUW/hHroRth37LA0MzS0TQiS2KXD7KKf7vaX4uGQ3O
cMxR5HbOMtU9tluHZ7DjGpkZSoBsfXZsZnzGx/K/5mZlq+5W9lovFQe12yLCTqrlNnt8cXZibFhP
yNK6TI/Eyff1aRJohoaX8o0G4sludYUpmv9nUQzXdwsi7bWupQqouiw7cTOmxdjBm4VLqs70X3BS
jtfwZE1giSmx+BfD7S1YvNJqrc9/iEldcGxFQ1xXrS1egKjoNDWhTahydGOffwAJTpZXSJFuoxcA
yNMCeb5pn2d/fQH46rFETyvtre80FweXbk3y0+nFizSf4sVUsE1pZTIzOTo3PyIEZGvtgFYkvPrb
CwfkPWJtEybaZBxi429tV1jw0LSuTrd8uDRlQyhD/Oj+VkQ/Sr9XKiFYHaxlLMcFiFkCWsLVYb5U
Qk0wC3BuyXmjWAxJ38Dszy3HiZs6vE9waC889C+842BavVEFEPn5uiuwXRhO5TtcX2m4qJ+MFlj5
08Z3HnIs+e6VoUUOg05ERkINwW9d+jU/9vmr338IPwyPa8Old6YzUAUuPX1eo+J8TDisK3CopQLy
oH94X5OJ68J2RnIsYBL8eqCgfDgOUim2tI+8hATm7JVLXo+oySUXcToAW97rbSutI7Ub5vc92O0c
PjHa0hgQnh7INIYZUKD454QR1J9OWl/S3k/Vm4GwebxcgsWq+B1W36r1CpTD5eRUVSfTtmjg5u0n
EFw3IhN4VblyrCSEHxJZQSjDThnNExpl3F+fFNV/YNc24d3KbE7+TTXQ3jOsWsYYJnXMi5ySsZ5j
aQ9ogtsvotIL+S508EtSw95h46oe+YLHfA22oYj/NL0LuFTyOU1tRpyzit9hhf3fYFaN1d/sJy8P
rCTVLC97USocNquF2Q+x2xdFxWsfOHxgWhmVLlUlDUs/VH/iQwGtIeF495JsA9G7pTKxKTtdTF+E
9XrTCHBfeK6T+Odg75j3KY2AAX4LZjQX/tu3jWnvNnEPw8XYlM9W1AKIEMVnfZOmeRqyJh+W07eV
tP0AdwdsD1fiDjwc3gjHgQVHz+k0ERlKWL+Lcbv/OwVciX5IfMgaHEipzNmcJ5oVNCP7lCkkiqjH
n/4TUtw5gh2Vk5lXAJrKE2gfpaJfg9zXjfIHJZ5Rn7SRUljUgDvbDL/jbP3W2X53y9spEPGb03xD
k0yaVI3DmuiwJ232i2Ce5iTAl3YyYIWZgUYz1CSQzS7+7+u7WpmoQXayywYfbR+XSYAR1UGd1ZBG
75cBeTF8LPjOzhhcUgGkoPy3+caOW8TnWzUzfwUv9F6fl1qPvUeOrVg4e7Mw9P+EC+qG7sxIZRVu
eBgqRDyGH7sL/LB9y9lITiVIXp/ZQ9dajKQ4L/4grHTjDH8viAlrm8ubIZYgY0OoZ37FNlUt/7q5
u1J9jlE28i2whrnbDDBWT4UvAud/WM0CiEYiN1gmFLmw12qeko/Zqs4m6Dqna1WHxP0bhBTnzZo8
KYZTD0TrfW2ni2E8uLAfFHZ/NDPy1o3i5dvhcxmHqGm5+JqoVvtl6rn5UH6YnrxfaCLS5YvVKN16
gTQTU4Xu6ZrkRK8tgndB8WCTzz1a7yFmyTLyZmJuMRl7IothgrhEq+FRgPkhMRVXK75l0YvTL+1H
ycGcmXIU69NPAJLw24/Uz1yr2dikxrPmNb/F1cRU81cVkiC4rOMdpuSv+kqnOBheqKb0f0XKIdz5
4DJfdsLGgbqn19A+qwpGgJiVhlEl/TExHu2o9wGnqqRYsHxbTrxSBWU9YangFiV1qQGIim4iYoGD
PY4y4SJ/gHByF/cVRIfTK3zmn4xIQgWEkvigbk5KTN9WMJM8D1iiohNd1oD0UuwiJmMRHUZHTvg+
tiV8J7cREd53SoLn9+n8Nz00g+jz0LouKMR7942Z0/90dv5GDbEPVilpYYEPT6Qyz27V8P07PgUW
j0CfVnZOv9MC1Vb4P7mrrlidRVoUwsdeVqGzPbl3Q0aaahUsHTY6TCkuml/r25GaOBOHP2YF2RgB
dBXE51rCF6l+l1lyYrTuKb/XXvcKwOK85BxwSteKY4AwpTj/NW5muq6b7HlfDZlIYJpLONqVLI1s
Ll3tZIEqAE9XRJ254WloXxetS9HaHbeyRCFeqKZEkPPMbevKnwtnXuDtOwu4S1K3UJvMO8F8cvtg
u1Is4P3AdV4RtDGJ4U3sgjvWAWb+MJP2/vhsycvylFqkqaV73lQ7cXq9cd1dwUYyJDagq38hiC8U
EZDp24KvfqQLHgE9VQ0PqITRCq5QMddzWLptWckz0SL89PnfiYfkqJ+/uyzDx3p1Jsoh4NeOXfqR
mrUxClRdc8C+tKhEuJ1J4U7JLEv0o7oJ8F+Pu/MH+oMBkuIPV8r702DdPVbWlknv9aoH27WNDFOw
qjFGClwaImO83toQjTxxTX9+l9U9/ZyKUu+9RnFv4USFtrwMPshMKgx59hSElkdtHA8MZAJCkfmg
7AlWf6hMy2pjdwcZdP2YGrFOIyJ6gpFXvPSxbW/JmFmqBPAL03AvdMIZhI/juoUX17Ph3a0DS+bV
28OTxnn++ZbkLD2O4S74Atn9gtH3+t/QR+RyVDhZAiMiWEVS/eyiQGIfx22gYjz00ttXoZbbQVxj
foK9wmgG/OKtYoiC3niq9cWrFysrWwsbXKTGtzwFGHnRSymDnucD/Hy2/ixTrH/d/Tf29XV3sM2a
yQ1fO77Aqd4jEsrDTCWBcjhY94NJlevjc8yPdMo5q+NQVzcfSfyTVyVS6FBqemKQbp4+MZl+i1J3
SUXJ3W62FSDctKRML/eqitB7gvaHz42cvBqku4H4BxD1yaNh7GwKbJTJNn74vIGLKlaLWkSQFN1B
ypWNP3EPawtecv0UQ1DWU3fDc7j2apyK7BmIFjB3KlAvaeLTxiWrv6G4xVHtfYqKnXTYADhF5XlB
vu2j0JctctW5mr4UPamEK7tGPBVtDjaQ8Aq/+OPOFZogEuuWrOSLWax7WFLQo3CyttWRXC+64GVl
OhXfDx8BQylg510OVzR62tT5QY/ult9TgVv3U/hSrlp/LcAZWS9l0Ve/Tm44nk+PvtNo/6/aUAEt
trC+fdHVl/p0N6gofEXunt7P/acRznjvnbBhWq0X7Y5rIVn2fM8Pbz4tb0mT11B+Qdjx/YtXeLV2
2JTCCJ5nqpKDO+rfP7DC0cEVjrS6lwXS7Qv8wqTLmFE00Wb3pB8LYiUGTK0oZwnJ/ssjcX9y/dUR
diMyhj07G8Y81f0BCyNYXJRxT/CQBFudjBfW/oBr/UIiAD9WSTo2bqnbcm4neRUXi9XtYYROU9te
NjacFLfJefrO0PIZwkZhOBgyIaXiACKnAtwxyi5lbjtWeNli3/d/aVaFBeaifVj0ZNANLbmlK2rW
hDOsXH9a811ajIU2hl14w4/QfadkTCnUM+wy0WDQPt0clh3QKo1Ma3sXxOiBr9d1b/beTqXZobMR
TwetnkZvVJpGUdv3ratEJjauE8tyopQJS1RHL3AZdM6QQE+TfQ7gvhIaFJhbEdlEoy8RJNMkWZN4
V2gshIdyEs2lwfGrfSpS+jX10Eh/usAANLyKFaIRpIZ4xYAMjAyR9BZ4jsRp8YG98zPPE6WCcPPF
Sa7BoBdosyIP/HuEYVwXQqBXGNTDEmUPeXw2fc4GN7cyfIpb0MxSnXHLhQTudEdubzVdT2scDPsA
CwshBx7J1RO9j0UjICvkQ/qQVwriFpkOC1Ez5UcLoTYeEzhzMMD+y6lUt827lAVKPf5LeGeaYqft
CyVQzA8s7IQKw3EFsPLWK9rI0g9eEny5TP/NnhyIzvAPE0sNkfSVie7z4JuHLeu94hywKMid9HeT
HbpW+bvUt5XEwwVwJtLx5unSc6Zp/2TAjC8asyk/qfi6P76wkzxfjtJwUdKVaHZ557bAZ00Ng4fh
mDasBgmmc2BH7aFuqhHRizyHxOwOc2UgP1mSgy+K1XVJCFOxL4VUDN5LDZ9/qYfTDTRGUOZF0dK/
lFzPrD/pyUBkBEXrdl7XBtOi+/0VHqfciG29wYHlRiBHHzTokm/9qvF8Nk136Cw2TemQmkt0ldwH
sZbuytaQOiQrPBnYOCqHlWUxpaIyord2tvcsxx9aXcmwogYuUxxrHWGyVZMpmi64eiM0/TteATIs
1aPjvQCjOldkWkkl9cAWP7S/lvAnBCN+YxLO2l+r3UFiabMcRK35nZsHLW3nzBt0qQlMt7GMCpJJ
DMGOLhqvfU5Kp5jgSwDZF8vAwg0hQetRbmadEmHokWbgVyUDLLO0dB+QjxWitCLKsXAKS25u/RRQ
M4fcBewPhqVv3xYUI+ZwLFbyO9pvOEdYZZK+J69Y3Ke/YVO9DV7iCcLb6XkWoXGZ5nix+WpqsdBR
en3pCVmKvX7CWub+o7kCN+fUDJ09+vmyBZpD19mdhxuQ7q1xPdjEndY4eKUs/OEsSyZqcUD4oug2
8HVFINQWFI61KjqQB10srsXuNJl7MiWTNrZAG8EkG+dnpecTkiHEdNydHW3J9TvF/TS2MHnx22bV
tSBmSdQ2LyeGg7OCPQptc6Gm7WfAn2Jj5i+5En9KQ4wwVGsKm82j8OWnfSnuWNxFz7GfXhjdzSlR
eeDgDUO2JcbVHjxjwaCL9+vaFB0Sw4ndPhBouOuMTRka/a4RrmcXUhr7EL7RvYk8unTXKra8JB4f
FrvyTZMBnCcTOFt25gbwIC+g84HOzujpXCUbSZzERCEV84649tX7F0xydyPkRMWJwxa1b2tgU07y
Vs7N30nmNMOsm2evxhIN4EwyoCaCQttiv7NeqwL8SLYDc4TTtAoRqtB8m0+KMtcDNgZYcooePY/z
oGQlhG1qs8qeXyOQGr82cbd5GaL679ty6fXkzjYG5hH58hf532NWpw+9aPntGacKUdmlAwRaZKfx
LZ8h0yA91dYj98X2H8NXsmjrkkKaHmnyTJW5/3tXIC62rXXKXxX12e6+TI9QDMDr69WIHluO/NHo
RpyugkM8kdKLkVn6ACkFWTWgFa3ycGFVy385WpNQm5fJ2OWpOlGfHcH297gqV8TYr/S+a3B/lqGb
O6jwnBKcFAMosyW/pZouA6OOtHKigaxPKOAhi/VAMvtb+Tk86eVmcguHC/qcli5cFfyIsKorwBvF
YABX6uTi6PtMSX3VHwva2/3lzvv+yIgVOVhjnY0llVI6GQ/2nOvEBZhHD1AwWVI+kRZSwexKp95e
iBRIQQvFw94AQQXm47ZH6Jbw0t6taxlCktS7IaVzPjqQxcZTm8LH4zYE2+y+sL1rFJaPw8GeZlRT
Tgf9rI9AXEPPWEjPmAzhMo5AMZFU+EUqfHKatKDVAiI9shWZt4UcRNl2/jbwQ13xR9KzMoQbCMR8
mZy6g3W8STaE/i95Bg4JfsubIJocRhUbrFsAiyaGlspnafCfpVIqW9y3ZjhXRtGEDH1t20/uoX9u
1xGUJmsfUMSQM2EUJvENhywZp7UpBlG21ZpvXL3UTpmFsc1lqGB2R+19Aw8VuHLUSurahek4mI4B
akwFykP9rAKnDuy1Adz4s+9yAFcxSIds4ktBq75XSHSV6ezxZmI8IBN5o2t7se7vJZq9NFt/2VD/
k8iHuBPfT30IviAfKINXmB351F9jCBBNVwfyTIOv7S4NwWd3nGpBL84Tjg29KnpAO31/54EuMbNq
9YB5nEoLF10vyQB3PDxPUr/v4jvbG0FG0zXTNfp3tgWtiFqUdpZ+WERlJYPTewRfqyOQcydqZdOa
gPECSMdPlN0qHr/+Ze80nET7iAvJrFgU/ndFHoYPsOIv+MUq5hC/+WnU+tbDcJ4jakzP/xZWY3Tl
1C1CR9/I45qU08/gJrzPzi/pEAVL1GWdIdrpySY893PRKpai46jOTOiGPcc/JI4ff/XjdTKRhBTT
z4N3xeS8LUzlETuEaxLs9ZxoPn3IMMUfbvAQWUsQ+EdgQEdh+47K5W/PkJ6bZ3s659WmRxaPtjqw
Vzzi/Iq5IH9Epun1EkMQU4IANJoJvCWlaZ+qzgld2LrO7Tzg11cWtP++QrHhBIwQ5ZkbA7IeLCCX
5NHa8SZJA6MW80q/tUL6L9ZO0jk0kYICPb1aNDjVvc91DgQaIEPGquS0y4fPT3QvI6WvGMj3cCan
u7itimXQV0Gm6rCtXm+8O+yfA7sGWSZFCG1M+zCyTfS+8VtF88C4BhvvqylZurs60Vig5Kty9qxY
bfEOmJvV6Gz9kVftLO4XLNQGffI3Rs4fo+PpCS1pUZ2BvWD4KXIvrudAFglhpHCKzVf+T9qW2g4U
bRUW8fOIKHYrnulA+qyGqUSwla1etfOb3oWL1EDtscA9BxOLwt66u5kxmLUP6rE9Y4plJQicNZid
vbZp2geCwWjagxIuFndzTtf4mpNkTpb7xbHFzBDf5GoxzVMjpkD7kRwGFNjKg40iUczsyz9WxgAh
YzgyE5WQBANG5E01ka9HLUSpFtYpB3KkJ67d5lI5hf9FWz4QaaUXmloDdY5te4BFq0BlD/6m4Z+h
pcYzWIWSC84xpiSD4xyhDZCkEp8vtqwIGPGnWpxDij6hJlQJiGGH6ZryrU/XVyVLN2hJ9cDu8zr5
Chwm26ucL1rL1t8Ky+OiIIsF/DgTCK37DQCMnbL2kOAqJKfYqLIKZlY3Hcs4M57+mR7erQSqPAfh
/Z7owydSK7kNUcZSb8cjniEmmvCfp6oqjrk7HnK/WiO21FgoMlijutjkbFPypKHlACJqdTm2hHsR
LE/UbzN6lUTKaCgg2HwPoLoCAyGLw2VBYQCWv000W4j+4JhUC2oqWy6DrsIpgIKP3GhObh9Qiddv
2kYyj37+W5QTvZmYjp2+RDrM8VhELj/Mha6RIhO/DQVsMz7POCx00Kn7wZvGEbF7fJ3DCkD4iJAO
VpHOHrpNk6t6G3V30U57luJ78pN+twq/LamnULqwRSfG0xxiC4/P7mwdC5AlZqa3s1s7pHlBWAl0
YcDyHdotHZN4EkaV8DRMuTmWHiI/CZGGYgRAEGW1iHtxC7JA+LVpnDx07WBhG47VEkoxnmMs/rI4
NkQsoL3KT2zfNNye4TenR4dDjyl87cNrXWyX+UbDAGRWsqDf+6gX3/ZMgyPo3JF3iy40Fpo/PH8m
kwTXgkQtsBOIPm3TTdLx+lg6xI//qJOcd3GV1U1yXXaJEGNCK97p1OgS5GPY50f+d/fN++1UR99L
iFtoHWcgfol8ntH277WTVt0c35Glel+0VdjHPFBAVJdzB/Hk24FTwFdXgiUBr/abS0ADgE1dGKn/
llZDOr7iMDdQNOOcoo9EIT0E2Wq7kbVusKfEikV85N45yNLOJHnq5GMWzWOWUDZKzO5VR9FGe1G7
OwgW2t8TthCE+goSjkiQ0OnNmEEFLFJlZOF9/s+/h+oD1Pvk5wQ0uWPjXH7R0xAv0mKm1lQso00h
kZIdWeRXyS92wevmpbYmqW9TkhcqEKnRab78BrNzwdOjJteGUo3BHpF0gRn9VuKTqJvyMNBfyACc
nbLxSY0ZtvRr+NOEr5eHuQQXRDHA7wIIMBBFgxzPN0bZBHvXCqudDEoyVBzud7LJwuqt6fUVXvd3
paPuIvgvShJhVoSlEAkPCfr/rCARXAYzpa6Xmf9i24d7nGAJYiM8ekNxwmFWVBMkWmioYt6i9c44
sP9JmlAmZodNTHStUiBOUPWLBZa0CPNn2buxBhphs3U45VEdm0hat9CoWY1b553dRVh5t9U3G8Z0
Z0dRzyvk2kOiwfzrU8hXbYAkkiNREnROe5fLP2tVrj+03/+bT12IJ9J/iaNFIbLnpW3tjL9BZITD
T7ZkRLTPOP4jfzpPxmR04HuV/xxRvGczuIQfwdzOeYgmAGGRoXRkH2SkT0HhhNxKzo6yQjp0DTYD
Vu8S+YE8+i4ykyIHkjbj/ULt2rfd/FCpDmOaGk7c4zaS9yl9xW1pZ6FjJ1T/I1RcbLMGFdA/L1Me
itN2zJCppTau/f//w535ykK2bapo4NI+a0OjV7y0li1s9HTB4HoK1en8GPyBectF8ugA1EguWLmv
nS975qsQjSy18T/7rPdmcqP1K22yNSHmIDKqHjmDIhfTrzlEHEY5FwYRbnTjfxf+Z0uLKw2doAVa
jGRN5VISPyDDaIKYNGlxZE/XgM+ToCzkH7e5YcSTQLveICBhLbn3RqehxT/UGREF0HKBr8W4oFH1
1Vw7ITOq8kPuhyQDxEMUlln2YpXtVjIIFhzcDnrC2XTJF/ULBwL3qFw1kAp2jrH3vpL1YjxBsmlY
93xVRowR39TY71ZrxvSZi8VdWVQzEQ0ebLhTdJderk3bNd3ACbQiST9tMObOX/HZNYDSvht/4NY0
JrfJUFxqRc6D3A5ftYQ+YK6JOf6Mh6cmK2MuI6Id8XOULgenIkRp4aV3ldOocLm4+hTPp5grQ0Se
MCEfYb0xXfCvrECmVNU86JctQyB6oou+BuPOSXNC3tcjboLh+Js7ZceF8D3WYHoEvhidfJXGfXAO
nz5thKNZmazbT27WQqmLQciDM9ahzBcX1xG6NyP0AAYPnarNeSNTzqBYdETFRYBeoMY0vwXX5r7B
glBDfrUStUIDrUbPz8+5vRJY7c7eexW7Y1T/z+bBQat9W+Wghaj/7PRgPCEGrl6ICe6VDZ9EUNUl
jv3a8mMIstctwtSZ/6xUbbwDcT0GXXTToS2C0YJLJcOMb7PwVn2ulalifa7QugXzAwdr0PvL99lg
PgIiYwAsZZv1VN6BAhL3dklYmyfKgN10YzUHRaf5E72NI/Gucio+0tr6J+TiY9DKriy81mwowHZr
Kw800aLea9a/dD45GthNwRWbKHJfVeJVr5xeVl5KFJItcl4+vkyRALjuaJpssqVarkNKAWb+/CMq
SibwETqFtFz0yBJxu8qkSZ3YdA1uTEejmsYkWAfCToHg9YSlfoYjDKhy1z6oVfQPqUs1rMe4Xzn2
92FiRFIso+yTb06IaFm4WJUlTJX9ANrcRvn0qGvW0XllIx38tkrfFq6ALjFq6dUnY9EyUFpAuDQ3
bb0rT/xoOfDCmXpwyUTaYVRW715s9jkSQuv2spIZ0XcFNZ+eaKYs+sdDKfOXGflrMVC0hqWqKLZP
bkAr+HW0NsC1Fso0NHU+0jKeHx9tyM7f8Wltc83/xtZ9ageqlfDS1MIBRZovtJz/JXg8vGgqIkDi
Fq9wxY5IvqXIstxnCLddTt5Fo45RrmqTJNOxTVP6O1jScfN5OE7fr9Cjs9j4hvydx1bS+VKgsHzV
S+Du4AHQ89ZKJjkjUAduuptYvQsYXU1MgcBtb0eKNaFO6bUGwRgexZk+KVwNARizzzep/jgVstOR
OHVk8Te+rhlJYFSybr+HmgOkA2WAtAyaFshfnOlNrz/tX0j/8yFhpgJkzhOYAPc4Gy7kGZ8Zdixa
I3S1Yd21dBxS0w/PnO1qWBjfykVXTFLFqoJYbm+aEi76lux+vCfHBkmENgoeUOQjSyPp1OcEQfwK
vSqqjqJSkCD/zYbcqt3RO42fXDgvfLxd7FKkAgq/x/CNUZtuCl48astUkfeQ0iOFEYpIt/teemtY
fZxkTvySXHQwSaRAZ/zWdu/r8NIsvpz50uUkJn3xiQpT1JABcZH8bQ3NbX63S0AWK6PFjhVJ7YlB
nDvm2MpNRKeCFM16amzViuwKT4B/tOyXEV4odX6GPv/2pQMlcZ7Hw+RlMnGlNRKB3LuhLszsY2nq
pmMrZjmwtUnCp9pZrDYf4kNfmJvACYkCvqcdULKPQpI+SdYu4WDiBhvAbP/StfuU7k0kWBP10vMb
UjeEYld1g8/RALo5Lz0By+iI0q70G1ZjdE+9fAvz6sW385qFhEo0DUiY4Zo+HLcoxxwDDnISZvNp
p6abNko2Orx0E8vUHUhfAnhDFxhWb8zo/KEPiq6G59J6G0hPgiFWyV/vXVqY4x32TuCUQB7alUxN
gTNftLUJBesY1xkeFT8dVgX8wc3ts9wcy8Ynnd87zMN2fRPmT+uZGFw8J4VJ+ZOFeHsWzHuqcMI7
EyGGJaGn5KzmjV58AsocGGWNJemyxS2wlp7/kOW2ekC3JgHTTR8MJB98LbCWCdIbO9qT6lksobvi
kyS/Mugac2i1sqWIB8rKWS2rtobvsnpdMpknjbFnPL+MMT+D7jeVsHL2s+/pIEm/CAkVnHAvsL1X
AJkuLbo+iWkD4s0WGYt9CMNPJawos2KsLMZ24CUjxESh5YzvYHXp1cVLME40aZ9C8i+yS0eoXqFL
UChvUiylGw8SwFPGN052WWfxzvv4jFvOnr4OS0Fk2Lg8Ic4PW9DSGChvrq6V5zJ/RaKz5XL0iubh
eAUvyH7vqXAFUOJ4fKLPu04XQqW2O8IuvlaB0eFpwiluEeElh5WEOnak2nJaaEC+9kbTiVPVYbIG
CNqSZRY5KJspnXIiOXBDG2pvoJoqeXxrEwzjcAUDLPVHTPdXBNaMT+oQHHrKG4pLv7c9lr+zdq5S
WGFmttxhA1QrhLjR5pHiVJIUrS6zRqO/GLLPJjka9sm8EAYhkMwuLMeK+A+CrAKrTp0t0/SwB93H
rr/vPDq34RiCJRqD0/QY3WdBySdcph2rdQdCfJCIZVHVA7GIAYBgKjUe9ZjamVqvdDskgFYBIPjM
mjFtkmhaVzJNQoyk8q3hoIIhdv5l29RuW5bDmocTjaf/6KKXm95wcR/BNplEwhTelQzfo5kwe9LK
6gfEo04eTW0RR8FMuFj5Dy4pSfw27DIYY7yd3NakS/ZbBJIJwn7PhvoKSpBfz6lIpPfnsXaekWqT
RHAU3LOi7ULsda4el/WUYd1uxUOfiIYAiqTEdZa5wQzEHXw8LV5D/EUNOosy25boYlRJ5VtagbGU
r10gHxe4sq4VGhkEvAzkwOZdXOJmezue/oehvyj47dTfmAQZwLQKJQD7NWGZ4mIoGqXXaG1kaL3B
DJ8yoFnWB+5l0m/r9JCck2hukmI6GED3rHTUl/806IE3bqRtt1xPyedWlNdF/bGz4hzZ/8EsYfiS
KJ9Z3oK+lZ1A1cf7eOTblt9xk8zWIQJdq61g+scFFEBapr2dEK8GzYdq2hM3rnMPeVmfWpBCy9Im
fn4RyPeaFc1wXnUAjUDCICNDvgy39FmCHmP8Yy7qq+KFA0Rr/c+6remBf5F2boZTm3wtarLQFgZX
/xiDEHGB9E3rGk4+cd2CjQBHN0YczQGKBaruloxY+086xrTuL6KoKXNFxDOSKW3Y/iZVSBaxa1kR
QV5c/nyUCZ8B8wAFUnQwdTPm0L4yObtMvJyIAt8Si5oCS6UHT658YzY1VX93qqCuAfxsArr6UG52
2sjDMA3GdiLksJGQ9B2Hob9yk7qlPH8GBwSrWKf8oSbrTH5AU5XdCp/NtK+vEkEyLo9esXxaneiZ
yoQLTHvrSBp52pg3ij/BedpWXHyeEeSaidx9UsxgvdfuOJ5Sh1SwpogLpoRrQFv1BvTVWRSxxJoF
DCTjm8p0+phJ1X/bQ6YZPFcDjECw0i39UDCycQuxDJivzKq+HW13Sdoq0IhM2+zUO1Ij6aj9tL2A
96Lw/ARq+EGJmXGg43dg39HJ/kh3hiA8s2vEtU0D+QP383bMnndN/3pQGyucPl2HlUU+l7FttXOX
H1nckmWgxz+ga77QThtN0ahRKlUalZdvXnkIsppjbqwxqEmTZEkH2jKRN0fTHgh+jIIZahon3qjx
tWQ3lX90dfYSRTRSSzL+CTxeDIK8CIsmL3GZKWKMGLjeTxGKVLONHjqT1EKfV8+pd/7xdgkPYweY
peYoOtW48BTQEeMzc0OlSDWFmKrk1m4R+KjtEQAVz/UTs10DMMET22ea0MPA2nDLplyJVzPTC4cu
XrxBy5Bn0b6nueYC9WDWn0IiAsLVMGChR3LBW3r1+Y+Gnb9mh/nAJJVKFdYShyL3AqMoP6QVMg4E
Gfs4t35oxLf0VAdzXuT4l8dR9uLg864h83KkstS/TjpSv5GCQlqY5i537ZEdBaL0oetSH8OpQwtP
xPW7EA/alV4nNrdiZg6zuShwLwvTzEZV+ocEALmSGFF2hEeqxnHusgBmVU90ZX82eFujvfDBI+jT
17UhK3VWar4zX1LVAZaR6+jlKuIaAYD+0TnaK5zam1HfGwt2lyZl62nSa0Rmx0OIkC27UDKdUOMn
w7zCDkD65EGj68iVdgJFf/vaL+XbBPiD2OReOToPbjeI6F7v8WBjicaWC/sBkADrgRSO8fNmT5Pd
DPz1J1rzTL2EB1WHoNBofE9H2QZ0MN7yp6X77vW/be/vBcTxz5zlK9KtWaYjqj4301qLC9dxh4a1
PpLM/c140IltNiQR4eUkZyeofIP6z3GRotvDD1yuii29VIpftCmvYYNTjW1Wk1SCL4AiPmK2k4mn
w8ymvX8D6WLRPOKsqqmc01ROoYKfhoLxdX/jCA1py2Xm9sxsE7rCsvQ0LWDIKYMhyzDgi+9XtyEO
qQutYG5xVonjjp2/W3tIRMfpT5IwRBmBpns3aDtDbv/f2+UNTdL9E3VQdfwCvZCATVG1vCeYzvhR
QxqB8lkBJ3U9cDrf+cKgzjNT5G6hn+5uOnyFrW4rDPHwV2NtRyV138guc14iRWtD11rpOVoM/rn6
cho32E9Mk7mwgTWj+NhuU/eisUKkW+/CdpRSpxuX5us+hKntmJMsPpN8EtBC01RtyeYGO8r52Fl+
zmIfecxpiR+mh3xlhGdj4dnqWWyMk6LgwxxzY5SfNlucaCgdvKKtKnSQnkR5/JgO62CXP2xeUCAd
a1RijRYluiW+UbxbTEmw4dsqL6BC4FCIkbcbNtF0AA43rFup7/eJYe9RtxLET9ZCt6Huv6gxQHnx
v4aLPA/G1SGmHRqMy5CoGPInVjlNHGia8XzaLTOUROzeaM14O+6lwNaLUDw6Pci/Aj8SQ6ycu1KA
bJxnO4fH5wof4KlAQhKgZROveacLBNg34dubp1ANrF5BRhx9z+lLTRfadYmZVc9Cxrzu8EN3Gcti
DVc22e8kDRxBJTd4eJYFVd9rwpCI92FqiHykDDDbBaHW5ESEetOEytahYD2IilaNeisg8QGJbFKa
JERxAqC8IN3kF9rFSWRCIlradJhEIeP6Awrny+nWVEdfvckIzR3ucTbquwVZ0cgu3W+az5BPUF9p
mvOMSBi1Zw78YHdHy9Er/izfdioRR17hFGQZyR+JvuPJhjBHAGEjt3wnJkQdXnExpcGpm9xYQIyW
gBjK9uJsnp+TiluCS60IY2uzb1sUUHcYCx4KEyMW/nfwOOeVdgNdfWfdnPoRzOvlNw/19s9tHIF6
DWbVxKk+m5Bte9kFgLKwXzX//753I9lmdpqMu3U8VtJMylXdtK0N5RDDNMgOg6mnHWieJdXsFrNb
AC8z0rPblNu0P41l4poAreoWHCbajfYmHZSkXyKBA6z2o6xQHcZX40ZdkGl+/pbaTlABHNmcZfvZ
VaQSSyJOsrKelm3rwR3B0Z7jt8SvaHdJdnhLG/LUJI3PXZ2pgFeGM8ro2xetQWQJy23BX2bN/rst
uqoQ+7p8SOGqQZU/p9/4QIya2axNebZESgU4x3VMkWcZj7X+YJHRmHa0xvpsjC5roAsQbJNq83IP
+G1rMciwvLvI3kGaE1lzhtCyJCO/LbqKm/0AFIxcpRTLnArEeswaARMuobEjruu1aCbjaofQavZB
U7pQytQi/WMqnlUzRdd+8DABg6E7tW49iFRZCnB9zFIcO2i22OhuF0GK/tkI8L5nr57YD4Oxae+P
gDuReLfssQGUU4pZFyNPN5D8qa7dYT68s9Wy/6HU2yx60bNXaEPm9nZXM8Q6j2eREfzTqAMS0d9R
BTk6zjE1rAM2u3otP3SXj1i4R4n1ApbpwgDREP+5kKHV10oBnOrOeLUc46Eo0P8fU6ZC4fyLZ4MF
PlxnquPGcZB1BDWTBjAfHZdcC01XvCzI5MUcGpRq1/xxCOufd0c6IqXVSohhyaSwYL2JvcgEkSHA
/DaYidXbaFgmud5YdrqXa7ycwmgZmQWj/wDxjOTshHyTqeo2djZ5h0qlxxgSGP86bOM0z9Q/MisX
Wq99oklRo0duA0/IGRg9a4dK45HY0nN+uY2kI8X2QHQs6jsAH1xojd58ahk81E1bLZm02qgxn4y8
f1Dpv5w9ulEKXMm5R2fgw76TjbEKmr09Bo8pu2GKjHmXVmcn8ITuQLp9APwXgryqjWF2ARuuvvJ+
3NwOYYhDN1aBGCz1woxXS5xwBFqw9LgflyFmn5TWV/hSy2kX5d9MpcYvXgyFkANtH776RyAKXruF
To4HLryL3jrsD/X+3gB0Wo2HKMiUeM7Mdybe0MkgoxKp6YBNKV4XABFZX8nKYNzGyWRIPxU5iwhI
ARQUZ9g/Fl1qRGGj1ulCZdWeeOJ9XNfg7A5Jor9Y86nhY32qMDEzKwPn5c2FaLz9O+foq83wLWpJ
HhFZCzX5v5BceeYSD6SuZ7UtWrYs2U4kNc77VcuebAu/FuDVNcVLKKQCmsJp28Z1JBiXmDadQa3H
zIBzkQoz4rFXJfaK5KHW9jm1vErEptXjnG4t8j7ak08KMQzgl+av7JV8/HW4kmE7RjZQHDe0foG4
qCAmiEaqBVeT3bzhByh84+k6/+AFoU7vANN+8icGP+TsiurNWKgZgn5rTDh0UwG7oWyv5N4B391d
9psdJpHTCI3FXKtW3jVs1JLxFEyLNV+Sl54SJw7O+Dxt84qdmrbI6FkvNmmq3aedI4apQtxmSmGY
Bef42H+KsEwLGSmzqEfcr3PHzA6wVa0x+cjhRp/3YKVsEuhNQiItEpWKQWwTfN7u8MwZV/AcjVJ2
NcngZcuFbiTgoUa9gHuhgERik+1exjh/jEi/Hr+7cJ6KmKsULAaZvDYaIR7hZoNRK4UFjzr8nIfE
b3mwL7TnTK32Vljr9vURbOyAW27qBlTtHmShjxFeTBdZNv4fYNeVyuaiRdCx2qKVqIyv9kQfk7At
rplTsb4Ns3pu/YUpanO7IlcNgflRJ9vHls0sDyg0tccTQrjs+XIr8PJxDkxR8LO3vg0NcWRQgBo2
7AoKAxaFRyehvpq/HoWbNEUDfH2fw/sz5KX0Wgxc6TckfrRIgkRrWlFG0ewJLCpXZ00NAGLF2wIh
xab4BFkqz2zhvdpKD10LxSV65kn4DZEHkNxJzKFzI0z0XX9jU7g7eEUf8Qgq0qG0jQcatpFOTqUu
tN9nxlv+qmBqbdJzYXm8BTJgp4XRVItaxNWT5LwIoQ4PU1W0GU+FyQ+CqP3yo2oj/spTpLWQkje8
S5ioHhomlYbPdTkv6EYPc38J3LF3VlKylSDH+1v8BCabP3UnDnti6eJxQwof6y9UyLlfFgiaGG0U
LwQgwjZNvYIl2f7B2k+x85Z8eHHcABYF5SAnxZqVdAJWlRIj6E48CYFItV3ePLOkVK3uFjDHiDpi
auTlJpSZ7sY4QJgQARw446FNUZrJjWntvnFHNryNr2o+IRuudTHytrzZ2X0vInw7SyXvWhO9CqHz
VJyZtMuZBf7Gq671OJdmhTYdNPnRY78a9ncv1iF1KArd5nCQa+fPNMTv1xCGp6WHhXZ4xHLhwXdB
gd0D7ZFsSWuXhzzbdzM5HCj+hCIJuOD0rNP5dsEvLUYCpeCusZ8l3uVTRYCxfGykMxAMbBmnPIVj
eB5IKB/9XPuOgCGg9LaYTaPlvj+vgEYPbUE2qMjUApRx2I7pFzGxOlpAi5xNUz9d0JkWI+ca7U7A
JOhYWkRYX4vdNmBtjGe6or259jxry2be/pEOvtOLJY/AWkGuHHSCcUb3M1CixBexsJeccVvUcuMz
BAn6zrW9PhY7FsrJ7b7vXKkDhULIuN8drPitIDoVkMwz96OVyvIfVRsm6kSdkbGvQyqhWhB7jSrD
EhH+KOJ6sv4BpjIkHnSnEMwohVGkrb0tgwbRyrlIAC3w1WnM8UBi/Zi6FDcVM5Zt0JZFXaOLf8DK
LFjNWVwsMG5hC7pKgiZvn7Jk+k0BpoKXy2zELMf4s19vVSZ7GOsRuHhY6Xjr/3WEN1L6B2JvXQU2
G3omMa5FH7hBMVY6tG8o7Fbh2j1/lLFQDHezIFD3uucyjmtFi8vq2SSQwMeyA09f1ZKGJ8NPI5Pr
QamYSSx0XgmvK1KSMugJUbtWYzyVRbOHAXOWi4fBlZffCR0smRsovO0pgoNG8EKTJnaJLIDjioZk
9oUqVm0r45dMpmrPXiicip+78A+CVbFuwGPUiDahBQZKgiC5qyRckA06rgZOWo9+FXbaxWpdYwBM
NNzyHoSagqoVSZo+AlA8XtjGnlV7dAHhr9laJHsiuki6HOTG/pF0+PMNOI4cozqOdhgpGIGqJdts
zK8ZTxNuhGjV3kHywBOJpmFp6INk97UD4eoGqcgtFWWMSlltwIM19rNJ+fwR5qfVfKBwb5+F941G
xaU/rIOnW5/o+afDs4Taotxm0989MvZOTV/GOBjVEP1dPy65Ovi+wf+lC99EvfoI1wTSJgdzfN9t
MZdK9txmUZ1/AbV9UgV3O4GWhty3UKC2YLZ0dwH1mJDnQS7mcjugygY1D0vEuRrrekbbDMrVgJQI
eLWNQnu+d5qP6rxhs1BoPq65rWnUehwn650hp6U3831Z58OLFlNIzlCkNzSiSog1xqHlV7O3nrPu
Fk09VhJc8LNZoWa10ZXeL4a24xCy2RLtVjvuyvSE/JoWjYMXB433nPMHzIPLnnjzn4EWh2/YfihL
hNOPtot4poXFSerVW/V2z6ySiPH5aRQNNxD0KlKvswK+QJ92XWHeCpMBpf1lBkGnh6buqpMcDHVe
9bYlqfWnpuqFnSaYgGKkwQyO7TFcVrYS6JQMyFFAKg4LnLRDsvrXrjvnxncza7T2NoxGu9uabl63
0o0HxXfP6c3xqgNsJ7xZgAZOWX7/hbfi+wvizfxa1aElSM/O+BmoI+DYekowJ5DIotv0dGuF6yB2
+XPE2O7qrV2pCzMizEpsRK92O4pPMc59D3m7RFqWxlghXw2yZ96/6wApOX/hMyYq27k6xJUM6cyE
203EUtys3Kq/RHLKRqJ8LRHGURzIy6EKpUkHenjvaWs2BM9hd0nYqq8RUKFozQZ6H4rUa9A9Vaxp
A9UoVZDc7mX9sYSV16utD83z2k/+xjoRSM8ik98nhGoeN7eoNCe+UbTCaFipb3/2FajsXX6UP5gM
UoUmqBGO3O1ZnNjHEAvpZXmZt2FNIxbS6u7JL6boCTiAMAvl8SrrjGhjRkogpauTVam798ywbb4F
ZH32uzzlTwplayHJIymMyDZCyAfbWWijCjeGz3krsCmMSeuZTaKPMJNY8BJcknmPVTL/oFbkH4qv
t/zn3pI4uUc1ipIdA0HJaAa5swFAznIdiTl1H899qZ4mlJ2HW/qyMYSv8WEPs+FPizlB4P8aoiRE
sLhmRMK4YvbQLAdJn+Q4X16FO4VL6vhLmAsKS+4T6/66820lE9lcbes8FZeyBnuWBOd5jkaz3CYX
GRD3NBg0rU/dqlLPMfhaeSgeYF8GUzjjv6zU96xJwj0LBslVvgPTU0OGsFzN3QONDU+1wbdY4Ewn
DPCO90sxcR02Tr/p1MyJlC/w+fS9+WwLE6vNGfoR2af5RLuhJEjRH5JzDpJWt4JJh2G38zZCZArK
/BlhnKeCsZhmU1hQVnUPgI52dFCZs/WLGZjEjmlbkXNYeGhFKQM4AyowQsL6Ts2fzWaF38qeEtwN
MIS2KZfHtujBdTZuuMiw/7ocQA0ZIKlLFzN8YPuEw51BOaDlvJXwotzwtXkkVpNERciWoSVK6QQI
aRVvYeEouJyioUsqjLSLg9hfcZGkhukps6WH/bhu+csNbJ84HKGMWtW0cJ3lS55RCirTJlSAlqov
bXhXreFp4ypj7FoCrUeXUNPCowyrmyXA4P0GMqafJCOZyvYQAVm7z/NNKzvSVQtN6JZUeaJNWT5x
3xHhl/ttSEyel8pdUQjEzllGs9fEbypr8Be+PGYXladAhJ7/s1w4X/hQgy8cw9lUARKP0vo1GstJ
3TBmDoKPW6eznx4BFVqSeva7yKsx1oVs9NnlMj3Un1TUnVVhOL1RjtNr2il31LSL7ZXbJu98Gufh
eB0s0Xv2mkAAga86K8wxx5kATLTi9IkA8lxSqq9rRo1cIhhVz1R1ZEmG5jHw5mO5uN+fYpr6ZVpr
+nAjmsg69zKfiyfLt8wm5PS0wbZvBD/ACeTOf+bG/5YpEzMxD4obfW+l64O/pzP8Y2R1dylWSOAR
ZLBd3peabNBS5ojZipQ8L0J5QFGt650QNJuvBVEcM3dYLWaETDqXltel3aUYLciEwNzxqsu50W4Q
4AYgBQF4j8Efv0nwmgEwP69mmNq1H2UJ/vCEuJTPdqUzml7EyW8z4jpqDqqnuC9kzU3D+XrZUaDT
U++OUHr/ePqey+J76bZBNVYysHu/FRsdHXUVSwvYUXJ7K9rdP467CskGkJ6PNsm06ba0OEixLOxt
TctS/mXtXOnEJXgSbep52BnQl03wA7LNxM43+ftt/a8iB+0p1wqhVGtstX6fHnWSaUpuEcfnOpLe
Aoft+HITbn48mFpHqiMr2fH+u2vWzB1BcnEvFcAU0MIcI6lydNXZ0i4gl4jGP7GTihAYELRCMCQQ
+BNb1b3JBPlgoC5BNJiDYUlVGGnLi7G2X2tjyzgzI6UAVdKDs66d9JQg+fVLDgWfixOiTB1d4M/8
XIH2QkkAgFf/+PcOnHYCWKdI61feRGsg+oJnJl0UfoTuiifqVQE8YoIaOiS4PoYM5Uy3M61D1DDU
wguHoXAGvWIJAThhtTM7fElORqq3J8hPP/wdKZf/d8GprINEkrFNpAGMHhkvgA8RiGT35OzvqZHh
/k8ILLCMe7PMakJ9xEmjl4xY4eeYZwD4GY8STRALunt6hvF5G5w7csZ+E5Bn67sV6xv6jEghFp89
RMwE6qSNQjNqe0krWcRXWv6zB9GfjRYtv1Z5ydCeoXv4/bXaD3hqUP8DAaOGufDvHLBQgHYNWa1y
tyYNnNg0TyI4NQ2GO3AhifyfIyM0bEY3QaBrovvINCHPlNKuk7UPjW/7ps7Aaw18blVF+PGOcmU+
b8mGRix+H9fg0e9gVTfXOgIGzL+mbiRhuojxtvA+1VlG4ZwyfdGQxr2nETOIJGbC9CS4gd0jL4BH
PPpb6lwC20IHwxypCoowt+rt0CELNYCS6wMtCE7ri+2drHCy7Hf8JaPvZ3vIjkeOm2B6bgIM+/6P
iVrT+0TwUTllQ3zV2wpMs3dTJAvkpzfnzKXg1+yjjrip3seUXFIwS5M+Lr8kBDjNrUHgKdiQw1zK
P6d4YTemnUA8PlRCer2TYFlQ7Fk3ftY1wPSWO0+oqyOMcqDCIejP3+07owF+AfG4w3A1T4qhB6rb
l1GHM3iNA04X9yadC7H5Nba3P3OWag274PTf9P1b6eerYtJq+r4HD7rwdw6eiH/xpEXvmdjMgoQx
bXlfZxBaq/fn240lulUHs5vSDFQWWiDSQgI6wBkuv0qHn/aUPV1PiVkp+WTr4X6COXrgDQQvsNSD
A0P0EqQVe3RgJF7/Oth8HyDNcqp8QiDiAE1Kde7aOV8TCdd0gNYq43MJo8T8qJCNj5UMETfcgkW/
trvuHkR/NwnXMaTK94kKLJnJ8p4AZyX5st/IZavC83/OgpJicxuFdRXi86z3KXSrbhOJeF8pexOe
E4xmIS9i1kqAeQLVY2hnd9117laCuZa7i1Vaz+nnno+lU4PyR49SAWoHQSfDS0MEZBEGR3LUSKfR
aBP0rbbLFIo5fK77vhTz8b7mug76uTcIdwol6n5bzJceBPzxbVSXJFJHIsO4E2g+NyHeQngRqzFU
++E09KyhMGQdLOQdKKICp1JlFZkgoJ8meJLXqX4fJSYLbZiGeDo3DEa5iG17rbTRS9/K+pJTZVmf
R9fdyMu3UHtRt1Jt4H6RYo8vM6AK03nOup+q/znYPzxeRAvJAk7PDMdJ94TClFanLvgfE0ywhsVL
SbesT0pP2EWW3fSuFlGxKEPkwmG09Cp4jmKhuVS6GLiSDjUSp0jj7koDiW/D7XHubGhDwVY24d7Q
hi2XcWknHjkqjMnBC+Y1LvS41cbvI/OjRnuMHn7LbBsHEKsDKcMsHb23gvng8Xrf3E7uBvFZfJlj
u7BCD15RiaYE2kDgtFUN3C56+ZpPCIOf2pnSlkR4GKUEH9JjykLsDUaXYlt62J4wfClw6mm+4vc+
bnPd2VSFY7IF5Cybh3HCx4IgG/xf0iZQHZPT21qIJxHvpWk0092fyFp+0KAfGVHhWYuEUOJXpQkf
pj3dqvW/rNr+ol15b6kHtCHtPBlpIB6bdmSKw0d8SCs5g3BIWPpEn9pnEou+dNyEwSpZX2/5MBhR
nmettt/dqe69slkt8OLfH3u+J1NyIBMCk4T24r2lVPloVszyGD5C4wM4CJcv2s44Fs+QICnVyUiS
MOPYC3bLOZn0R/qgpLeIPT/CSWmjYSjoO90BE0w3XfCIl4Rl30HYbZ52VdYXruM8KRk0erinzJHd
+6Q8akOfRWRGvjXKZVSfUXnVnIUUpUVcZxn4qMxaDzuZaEacpM23TstaZkG+wJsASMtD8qbY8TvK
JsUDgUXzwDLREh9hj0UQ4oHoCQlfFZIAk4iepnhYZUMmZqsVgQyOf1JRHpunV+Fx/0sq2CvRYCmO
BWEe1SCXm+wrr+59DLkF0HvyvGaTFcE6Ixa7FX7aYEdP1QdURT4CeB76WgyWbf6XuKn/eTbFiM7j
QrDlZWYk/a/vZ4j9gDS97G0tmzTPZHONaeCoSFA7GiXPnVva7+AYCnB6+n797oM7741u4fMCBr/K
sLn0wM7EIFq5j6AaLfRR1YNBStlKRUrFijwk7JE51wLzxHlUC+7IZHirldSzUQ69hdNwbb1FRxZO
AKziHkXNmCf0Bt/FPNYmvVEBNGHKhPVw6Zjmrotfq8E+TgzWrq3GTlBWpHTQQwfIUWza2/fNITTd
VuOsI4wLyxDGLXAbwzuY2Vn7cG0RqWo1G9QkpWr7COd2iwZE90dRMXimYPh5fPiPFme2hColCvsu
YQTiOv207JdLCey9pN+Lxo5eYrjciyLiixtXMXzPa2h7jwBbIxjz7ot5GWNp8g35ePXIV3wbHeqg
1qCQOJhG1EdI0Ko5eK/DQcAzgOYbY0GQfaXVofCHpH5QXYgrrNLE/FewOW2llXfmKsJ0L+jy93yL
DFS8Cju9gtiVR/fiCmTGmMzTFdv5k1b9tiiouLn8UfB0//Jiy4HeeNyXZmZgY/LKkaZt4ifOSVVy
dfHNqFLz3HMmjfiYgLUM61ZfwQ75uSfjACqpyxmVlB8dBC1XmPWyZ/4Ni4IEp/mul9mb0Comb3GT
tjO6/meNARD6uyTOxPnicU0fuje9jPm5GC+hdBMK3IjP6lNbrtXz+QkU0PEU/NR1hb+Mokz43Nrm
dHDCZ6xnme8aGPmuBk9jvvDl4jwASrUqtXhHBbiFWH20uwufIWL14CN6kQ2Msr/5WdP4CAMBLHJP
s62pVOdLIR0v8TPn7uNh9kBVrfByJh1Q4YVYuH+ktEWAqlRAa2Y3B1MQfa61/FHPRThJbwLIcKRM
gbJ2/ztj/dntEK5u/oq0BEQww9Gam/DIIon827BmIbfvwhD7SuCGmml06OOWXb3LXc+Ce7xeXxJY
UoP/kWPD47ArQhXN6I6RMnANLB3mXB5on6F6sfcGig4AbvSWt0nF4SqqAQ3KrFNnz8+u5NlmjeXx
GlLUYWSzyk33taJoV4a3UDwre+OF4i5lqEG9tWrDd+7HajJvij4O1JFAcKJK259GqlRTRTbbQxB+
8u/W9ccZZ0NFUvU52eM/0kr1o39+WmbyTw0r16ZRsix+Flcaa0o4rw560ShsgnBqgu+s1MEdaTnq
/HxTv/A5atIAdQYrmmR4qHo448Wa3oCrble1sIQcysX9dTQoSVvSa17E2Ckx7NOt1BOSKgzYKsER
wBZ0eQYg6MXTZxhd5f0AQLl+Xa6DVKKF2XxGAfusYmNbiaIzU7HSOcbkLIESTSjWQvVGMMohfD2d
3EfSK0mfszJ2QsEJ/3+WI6bP5DT2xG/LPnGvvCMzhV4+KiOJQgba6NkDKpkXa0ANvVII+qtb5f4g
+hZlnGg3Yib+LkgEzJCQDte3LTQ0ZN9l5S6AbvOMFnNH5Z385Xnjze+rYEKxSUq/DXJxNrmhc98R
FngVoz7xzFphoqRuw+OgQPMwkWce2U+KGQhXEMB+wCS93xAV5rt5KDRjiOdugaxaEFHCfXkEwtpU
2ozId/PLxSiSGXY1AfTDvQRAkSXbT97qOCvm/gEKm1Uqh68H9dsiGnTuvIC9zoivvUdLh6WdkxPI
doP/akMgz7Aji3Du3yOCRComKxWcpWaWZr3dKnK9Zvl2wxRTJr5F49urwScu+LPqMmGFpPOFuWBx
BVClTRXllYWxUC4qt+WFUWMlsbUi7m5uhhJKsAXChAdtFvXyWGwBHI0v0XveJ2PIT5xomMJd4OZw
B+eBvC0IW8B3w+8kuNqe1zsLqQvJa5TlyX4y0t157pWviD8d3PngYTpNW6VkdhPmRRzHnNmiWw9u
6IZKm+At3H7V32CIjhowMs4bG0TbA4ia8hejPt8KMo9VVrksCu/g74Ln938BfHtxI0gEmbnH8EcY
HPqTIKvs7yZOdPjQWGbgVOgUKAseFkpsYCYWefvTfNyFZVL6iU/2n2quwfHtIaGBCKTTHl4ql71f
/+fb4q3D63iJOTVfmWVPGsJbKbKHdy4c/ph9mwvCM3bzBNhI14ApmnDfipZb+DVzZObv8OYMxJ/e
CJ4BqOeqoog8qaRCRWppKSJrwJr3p5hwZogjwi0e/rLWRWoMLrZ2PDRmcpyYMDgGMp53kpV0qgMa
UrLPSIW2xPCXYJ2hmUWLWIibOYSpFphER7Pu7Ml/sn9PD7BpTRm6gpTQjEUzHWyXDweH2NhVi2Fj
hr2ft6Eq3aLUqyYu46WDdp6EXjAKZqLWCcdk7Sqo9e/l0Ybz/H8cYUQr0kT1V+TrqLxYhxPZmuhi
kOE4DrCTPvA04ZhWeSyl12WAqb/V/1BA9xfiV4fHcb94Jc16GS5hJDj1KuU4iD+4qSSpVPx8mqVU
GfQyaoQgWfTyUpqnfOHmCE0QlQ9BQr+GKfDshTD49KLg/PhF3UQaphzKvfEliwXjRv9WwnRixW1M
bCtDkf3u9PGYqtusb49qAUEHnTgH1s/EMkFnw055N9/sJoZNH1HXfsyQPV03gnVgqfB1DQvUwuaD
nq9c/FDmoRZl/+jCjbp/CNB7U1sLM797P28kNfFnR+5ncz5y4TG9AZQvtlBSjBuZxaI+PYjs575o
stiy/HNbI6WDZLlBZPswOVxFL8aaQR9iX7gB948f3Du5CCpv6WD3AVosMjTcbXF/l8YhW8xhx0Dn
DAphhUfKD+4fo8kjtR8KeorPsTc4LY5ohNB/P3R/7fSZeMpO+6xFotu0AYNlhTQuMLgqAnHIkvHx
mMwPupUA1HlIqznWCj8bHGdkUSYNCW5BhVFQvbABkqv1AYCa3PYm6FsHbSKRmxRFwObIBBsEQiMP
pvDRhAxfVEHHQres1zl8plMEc1bNX1/V/7lGOyi0sFilK66YaKOHrgjTXmA4bjK0skRaZUgdV5LR
AXiJ+TAXww3tnPIp433hHkaN7ZZND/MedzfjWE6an1xnlIr4pOdPjuFmmZWxHkR4n5Ee/X6Blg1G
ZqVkqD+1nG0ClAZxPtYSnWCPIJ2+ePghRzzF3BzZFZuk52vf1y8ZVOrOVGEvfP5qNxxjJxeTngrp
tTuq4sZ+NOJU7b5KBaSuD30rH84DyR61h47vbWxwtY5idQ/qWmVsYfY02x9W1L2lPLomsaORVHgz
lojkVQLTVEs+3pHzag7DHQCGAYXAZU9ZFnNeNdHa1IKcAlMtMa2fXxtKYJaelVe+M4DX8gUCVXmz
nW6mdY7Y4wQyg9hBxtdSyM08avnXNhTbi8ggc50s/8i3Hmsg0V93tv6vxrW0/Ns8CF4oKBbPTZ04
j9CTTxQsgPKdtb4i9PmJAkAQE7NDMYm4d8w+Buy+IagxL/HWpAWVh5m7WhUuqfwlyl8X2BNUUbJM
PJSFMWUUeHX5evIKwoa9CKsotioPjMPxyyk/z3zv8uXUw/nR7FJH0g99moQzpPDB+fTFWs8KVPFb
lnPq3Mi0hXBz3h7owHam/BA6EkUIhXiCUIVNJJ/xN4ppnSHeQyvE21RJBNakV7hquolGi+N+2IIT
UhuOPEJuer1c2pQXjDskc7MVR/izguVmhW13Jq75joRWqL4iw/Dl4BB+e+cCotKvFKVOiflTJSE6
wgrMjLy7p8wtVIccCLPCDX+DG1mHe/3qByveiM3t26/CgloCg/x1gVaSi6Fhyu8Sx29ZL9v72RBd
BzsiddlrJwnV34rAQW0aKE9XX+C1RC5Ld3MzycOt2YBhq8zOyZJBsDrsLbBVjctBy4SgNZO99EeV
DssUA/VM734nrSJn3dgRB0NhRnkuB+8yH8Hhj31h12el2qvYNWeK8sjPt0qRZ7KH6PMhZEBkU9a+
UOuUd6aPXSkHBQ99a4rXTAq8JJdPlQL5Zh/o4mkL+SiGakb/rpQUdqOgzpOJzfkpbrjhq/iWmA9m
mp2MoDnEZrXbHGruWaru5ZRH9mpcpe3kzlG86d5RVB+zNbiRT7x7FTjoEkLrMf+CLZG0Fan1XoBj
raBDwV+Nh4hdCBTvTkoXL6j5PUWwunh3+rwjAjkHg9FjhKMQQSk2V38CuNaw8qZuWS10qjlXMTgi
rOcwBRfpeKsE7+eV2OKMgIxHVpfdE8wbs1bZ8O/SsLq5KCeVUdeW0IUR7pGpPMklTu51gcf0rkF+
wdtD1Hs7P6haOxiNUIvpNkA5donnUkkUG21qz2viAHN6cek0mOcqIlfVHshOrLVmzKxJZvW/Z7MJ
TLh47wJEeQegL9QtIgoSVHAOxPHOBGJecWTMd7smED8ObTM631+vBf6kqkh2FImBfiwNxGsoTUbp
A8AnkaFiwl45i/o+QXNSXihFbdgxIZPLHto6CzShGr4iQrioyeIRUkxaYh5FpZdXN8Vg4t36Hd3t
tLYDPNkMi9z62d6K2i0rPoTJpcCOeUjybk/I0dxs+++1Z669B86dfN2cxzkPmJaR/RLgnXNXA9VQ
YdE/uXnBwjudxJlWeFGGZJ8pOFxBv2YFMhdG1J7jeQg7wnXlYP02dPuwOhrLigvO84l1Ldi/JE7p
TDBXaMdl5zyI/ux7pzDSxXzUrsbGXeDqX+EseLwxEfXd8MXq3q7p1FEKLxV0vuRGjXL+w3snnxtf
XFe1l9Jh0oKCEfgLqseORSArYXq2jtoLdtRRl3dmTyw46vT7D94aQr9jkPk+UMklyr6Mu+ILD/yY
tVgY7DH+SJ1gxnyfE5AfoIdA9xFWHt3mQBxV8Ji8GGOz4Dk26fzRyjcM2dppxRFJ3/DF0wIDEr0+
Y1K+RSQ9+JezGGF9kBx5hoMViVsIOWVABJ972Mb8szYsEQyrbNcT9nQJEt5Q4wwueK281CddR/9s
1S/N2+E1EqxGn4fiOjbgb44U2YMkVc685HIOfSnloXF4IBgQ5zWJMMMyAtfX2jN/IW/VMyK21ddg
nVU/lIEcCYGpepSvqBsIxCLnO3owgWv9ksCX8j5SGQx/s/q7RuA7owD/St3geYOQOuvH0AwmjeXa
kbCby/F7PcocG9wd9aTvPm0IOT5rsN5dAcSizZfilbd2QuQOGxwab3RXjBseCbvHuAhnQOmBvtpy
FDunSWeCEsBem7RiEYRQsejQ65QboM1KC6D3J1H5etXhet70g3VsPqupdvjG37ObCUEjae5NFS8z
2+SPMGlOCtvZU/TXMKSnkzTWfE0LukZ2+sXMMPaDBjegWUm1dWH0W8ZLs4KeymUA0Bw78Ub1MwcW
l9KuERxa3Vj9cwrnuuCnkPMQqlDO4ey+oQBbh++Ms8x+q152GFRoy9GLUvDDKF0NlVuOJevg7WIX
Ei5S+vpB2piQlUlXkJbj/6dOeSg5nUCwsi67rArDpWPMgIxo48JdU/2ec175pdQUFvjhdG+o4X5T
gBC3X08hjhBNQkGYewJBpryn8a2HKvX9RpTBCU4D/AUrv1vjsD3y50Fba/W95WRHGwFdFpAVF0k1
ryzBf6e1AEjMZ1WBjvQAhH2DwMkEnb3x9g2hZt1Vst/3EiIyM/QCfimco9m1/ghoHAOhqRAhxuN4
UItJpTXDfdrD7fn3vu9EBwBMlXvXurFqYX/P9s8ahGzm6/YHfk7S2hhSssJSCTjnSLUiFVOBSOLm
eepiESNzhf0DrafmzsScurufXt9ndESPSJ1/1akLBI4cs36+uoA92ilgdycIjyuOInLLmVi+N1j3
WoWlTZ3fBYIvWR4Ys5Mw998SvAZTfh7rt/jeBwLUj9n9Y2EXvO63uadewE0SY7DGDMt2x1POx9N9
deskhVYf5S0Bixbepj4t5BxzhBTQXLdpjtfJ3+J0BsGm3JYL4o052MEpKsPtzuoXen0T2xqQ1ga9
t2v6a77BwgCnoXjZZHRwNRRCeoGVKq8/EU9IQdY7NpydgkE9aNWBqTT4RggoSyt8RpURDXCeuaY1
VHYPo9uJxxCUEI3aAuH2Cajqbf3rXy70cPq5WIrxm749d3WfnAoy43kIxlOuNHgyxsj1hAUmkMnE
4vkSNJfsAe5eM4/u2k8bYuPhDhUdsSvmnS9s0y60w3t4DykX3RN5yG60hHUOQq86giXNUvAcWk1I
6hDSvVoyYCKqnHP1qSEbSFmHkVrmQMF5WLitHfIX62rbkT7DzkGkd25giWOnmMT2j4IjE7JkdBEt
Q2ivJmGIaUr4Oxxr57zG75idkR3ag75ycV3+TeDnV0GVcRXsPvePZMzWKLQn996HC4x64X7L1RjT
QocGryx+TGGRTO400w2loLeIa8Ag2WmU908XVmy3I5D9c/IWprayt7NFcdwHx/mfXRUgfd8341jw
BNx52XEQUHxDTQ/+oBo7TEpHBQ9rFVAPbOJ0pcvDKrI6tnpzVTaXyJLxkA8zioRy+MO//9Sq0MEA
yBPocg8DzQRwG0d4i3JnDLiSb7J9a2JI2L+Un2iWY/LUGcPZYV8CUQ33J0/Qgc1N8h4ktysEvXvI
jSWVGUFRx2EoFITT1+l8KyjRMELheFGW4B+1ooCsGkbw4PDIHhF757IfSD+hlKjMIEYmcAy+lvyJ
e8EIxksHeqNwtt3Yc5Qtc7DODto8zIHqpHnT10q11LUWaIwwOPWs17b4zZsPp5KOLCWpR3Ygz4Zv
Z8Qi/hGcJ/mGEYa9yz1lRNNfuO9I5xrfEmmzoPwtpE9oEyBcysOOJfcAxIGWoYuARq1A9N/feAgb
czrHdMjMFhFUaDgZVENG+DkIFZCgMgeLiAJG72KoBQFmZDsnmWAPnvgcrS2JtXRl2jgqamB21e9+
OuW7kjqXxrfcHASU5CDy0Fyjl17GH+9BgUtVfwjToV2I3fEKzXLLOOjIbLkpQQpwEGPzpd+29x93
5WW2EphaZYwy4Renj0mfbxBEFz0wK19/+UTWZQoiMf6m/QoY1VlAFWy11fgJgqxe5Tucw3qwMW98
PF65IAW1QRQXjMPYz/3vKXPqPiwi5gUrfku7WNg5yjLh+6VGVmoTb8Y5wap9JbJAZFnofXQF31wN
rmPnwgqrYPyGTO9qj/JXT4kLSOM/mOCnQG7nLNnHp3YflggpfdJHISakaWr4YFc+gfDQHYcceJlS
/hKV1/PysNZds44t1zGeJ5TW4RF04zp5UlRNiQi8c4npwfNPPAQ7i50PezHFdr4z5wFYJ5UMU8Qf
Dy1raE0IT/Us4zw/nWnlyHllP90IIZbXhbRg4ayfh9XSg7pVDNrI4MPp5T9RnEJjkfzrDO932ruX
3EDLOSbA79+38/688HEKGRFkISWsDhpCnchCxL43Mcf2LNlM/xTQpZBSNU4av8ouvNDjKU8bwexB
y6dp/BNPdNAT6DRVyju8E0zEmenlNf4UJLIdsrZxnylxGr7jXr1uEO/lQCjMEmv1B8b8Rq3DgoY7
Szp5ma72RUByxad+YvXFjyd570ihF23Vq7buKRYcdYXj4C/3tAp7MUCkY33WL8N7TAvznAW+r2Ld
dRwNQTx2Iale8DD0thgts+e7XPlPYVPDWMLHsFB0VP4OMj8x2cQRECBGUURkJ4aSVj5BYf6QSaCz
hquXkFYD0s92qOnI87cxbfAc+r04joRG/Vw0z0o/8tQ30f0m/tPKtPwXOlCGmkVSJMjAD92PhtoV
tQ0l20pAAF26UG9mBMFLMgzVIvQi8an3GC/i2qJG/JvoVXSn0ln/rgB9v2YEJCLNdTKCiWhf2tMw
omU/B66h5DckXl47yLH3F6t2YetGJbhB7cZum4zeWI4Lv/wBlJBXOr7iP5nl/M3IEz5SxtU6OnOF
RTzDWHNg6StgezcjkVBWuf2lwqvBVmyzK4iFj8NpGx7A/bdolYcBlJoU6QRAgFc5VB+WxFUyB4hk
tgO6qYPSOMAFob4yaOSPaswLlxZKYYygMHmKcSiEePhC2cd/H3JgDxDfTsE1GFVjQL4YkBO1XmDD
+u3v+s05kMKSucJ2APxbqMrqU7xP+9t54Gk5mX+sfyGFqJXqBlKlxkPeSqiPxTCngTVY0yK2Xc0P
NP6hPyNtD7RD6de/TRacKWoKVLKlN7IUVmV6b/4B4PQsjX+COGsBj/bbTZWzwW9bQRMCedySUw2f
zR+jYRslhBD+4TkSvfjh1gzYja2dSlDLLxop6Xgn0Wia5mloPGHV4CSKp5vLX0XaIpCHfsTbK8EQ
XaoZvcUNbKBrPcQK+ElXxlfgR6EIFaOznpHUezSrKSNbsTyK8mt1iqRSBIdqtGuAiBP4V+mZDEqO
kmC4iDog5AIXwjZ2pCkL+6TLUGf6V3qfA2F6XEq0hOBLXzxgMqZvz2O4gc7N1MNTse6G7l/nGc2h
i8U7iZFbmZZo50PDfAIAHj4NILraEN4WnvZpb7kFyF8EiCDhcRX8ApT/X/ZzKw/5RB9/yF8N5FUc
V/qw7yXpmDs4YxojZkvXJTo20MZ1sJKNyFJH2I8ZpIEdkbAJu2GyTJ3GRkma9NYO/hgj7II0G0MH
byEpy7vxbHmrqpRkGDeXDFZ7UYL+GjgkFtq31+eZxEY3fB+ZXlyzZ+6QmF3zjaPGbQ7/MiYi9Txb
VffLnuMKcBgdqOU0NbVQ+3YlGgSrY4QuDl+WdEx63XHMvZQfsOPMmEKvpxVpyFRLmfys3+1w5WMG
g7BeZg2B1sx06q2F35w2x+DLcn8Vuv1u2ljR0WBjT6XBQcwUegdkY7nkcDr8ww5k1dGpgAVQLZoa
skDODdb0Qj0yr0L0cm74+3/GxbnS6LllAjo8+hbVbkEzU4XV1oVK+USlb3ooGnPMOfXrVZUuqGea
H5SJg81hLsK87WWA79oqVu1+U5I9PtyeWcju1yD8+PyEshwkcqX2pvtipn1aK3oAKUxNOaeszdCq
cOSvXNV4rmPlSHW2orx4bjdsz4hL8DVfsayPwVYX2G+Xk6ab6egJ6d/rv4adnmIUapGd9N5EwOyi
mnVgJ+vmw0PIkvYETSEGNUHkxg8atD9cFcGvXu770pv/CCWP510fMfKoQ3ATYwGrZdzdfkftq9ve
cFfK73ndNM+c92AtHwUAA4w6ZcJ6HtyTYD579/nKXoi0WQOOx8NjR13f1QmJcQA1XHvqZcQTTEyk
YCHRDlVM0uwB+0bRNgmLQdGiuw3rUcdghI4v+Uyk4nsNCX2sjmnvDGsot9yjYRC3L0272cLedHyP
RSz3FZvB31aLkr+cPDMgDtatYrH0mGCvmITZ35KRLp6Q5NXv3TggdwulhEabVWVcbqPQLI3RZUBY
y4o3ULBRwF7NVAWlac8UmEnX/0109aEFU+3OYzA089bwCb5m3n8PaxDlkkRW1Ha/DJaqv8qnYc9g
joEIU5DAfgc0/Mdwfp8Oj413ClFePIvjVxhqU6Y2RSEsj47YWuP356loJpDbqxSWowF3NWa1fPZN
BSRq44VMuXcSybBJfT8Fl+KYeu883ijICfiiqTEo086hg12aq4/lpC4nA/lBEyDyAxct+H5wQq61
4FP0aW6VnRgxycgjZ5gF9EYY5m06FBEMUY5NDSWBjnuyaY7fPTR0RDzrA4cnhwBgqSt04VF1aJzy
oOHImcIY89OWWAV6soTiF3/qOBwQRdeyQkrixWTFxzxjUQR0GLBroiGOIjAmPun/go4EQqZpW1X1
tklqxZS1AjeERhlvzpYCMKPzZSK6wAMZZyCQmObf0FTRnk2qAnLJrtrkj8CFvSjDH/esE9ZL8HXh
SZuRxYlr9PIsZqCzlUC0z56nTGieVflXKbLbj1h/cIFJVV3iI903P4fUO/fZl6PlTFxbaaA5q/Uh
TziMdcYNOlldkDdO3cJiVKYDXX9wg2g0IvVFaKeS238WGeHX4SN9xf+e4FUOqs0D/X3ZPjTbUPBd
lOJzAtjhLxSeTyfH3TUQBeuEPNlE6RmtAR702Veazx0p8vMfqIOIfejygdl3EigCCpYWbDGuIHxr
z9C7WvuuyDeuOQ+QOhPzUNXk7GrpX4FlxckRy+vGNUcCoKzEiEkriYvQEOdUNMx2toUL9iMFEYi5
3+8wxuJLqcsjNqPPcYTiIJKNC8BgXFCI6Trfd4D3Ee9xmr617Bjq1L52Yu4BSM1dD1ozBtqgAmYO
KAtcOWAm1aqe1hE00rZEhs7nEqCvHxixrQojQ4BwRUcii59vrgBni1DiEVXO/dcKFrmeG0ZcAvgl
vvYYAyPSNJ3uByPceCyekZfsAUvlDRtBxePo7/wXbHD8SQJKs+vqGxM/9vOPhcKWNOY+ghdQT+VQ
ID+Hbg0v+lqb7JL9Ouil8UQYYHZwikJ2G8q920OnxEw/fwTAhdKjXCOCK0g26uuZFgeM4z5rkdAF
nl0ogDTPJBj8DLYRZ1OBFvBO29bzu61ydT009mScpru7X8iM1d3ZnEekdTFiaDJ7PAV5SIkQXM1b
U/0gAHO+mETb8uxsiqPvCSmNO15XjExR7ymB3ES3D6cJGQ6+SP0eIrgZs1VyeVldQyoYd9sF8tzW
+xK0LaRzeAxOW6rq3A/y4tUQumxHvu1YQCiBcEfAgvzfTVjlgDSj/BOnBEKw3izyrEz5AWjwkf+1
F3VSxQvCCseRXY14NJWIYXbMxZRZFjctlIOMUC51HSChvGIbb0Wk2VFBDBhQgG7PIjBhPOJKrzXn
Phbr8rmCb2nOKXZdofLVAPpsqXYhKGsBQmU2s/1VWzcVZM82ubpnH31d3JJwKWKNqTO7sxNo0ilv
CmF5lwASw20NFDfhJYRy2P4WLssUzrWA+bgLvEuZavyjK2B38cIgkKuyYoFGSyZbqD675LwvCPPC
Pcc//52QEe8LfuDh3RCuSHPc5V5CWIeNvvHawqQbiYrWQ88h1r1NDnjmEdj7HjgXPAgVfiBtB56E
3uPSzM+rDkrLB1DtflRsXTURfoOH5swetwjRPyO/CKOY8xG8tx/HiIUMy3r8t425wm2byJc9doqv
nVj4hpymRb4/cUgKxUkj/7fnhX4ieOH+Ug3N4dmK7U8WlF0lGM8pjs37v8eUhNl34OeMObY+BBnM
+GqorCIViIM4RbFiurbuCn9EI1NjBvEqToWPsBl2tCMPr+n1TTQ6XNaqSkB21UFg6m6HMWsqZs9W
q5Pp8aJetb0MYZrh+RDv/CKhs7KEFN6zeN7s8DWUBoo9Ezxe3s2uyw/ghNFOCwJy/TekfsaeCf5B
57Y8dp6S/tmUxPHLLR32f+ex4uCPvofMhD5dWuyug7vUNgT2PHEC9SXphV+szypt9S2JWu8weXBd
PBw2OhSA6CUttlsi8gZfw5D2CduuwT9qyL4Dm1k2WBqcyQ/8C8Iex8ruzTDu3wzfeajEaVif6SM9
TGEqdjTgbUxuCu++WSZF5yh4aMomPEmyjuwXx830/TWzuj7Q2YfGq6BQcoeqWzl7RcO9o2BoczlJ
Fr3gy/vG0sWEbhDlJN9+fc5h55MSdNLfJcxbLmtT2eXlvuDrludy3L9T41dy0Ecfu/2MU+R2GziS
2rRGdq7JmGCPa5defRFNKMMix+UImsEYCUzRBGhZijjx4E3MFflw8a0HYSsXWoGwEFM/SSTE23O2
REHyUb0mLqXb15peyA6DGh9EdncDtKIcegb5i7AnMbpVne/cxfzzaGupUHgfqR++WOHdSYXnLISv
RoC/sx3hymeVIJinlQDYvy0/Fwj47IpNQ3MRCeLi43yNfiZu62816p+mENxmN5oRP4t6UXY++DHk
1DHE+htbkAH4zpVAi27AadPFMTIsU2oTCgSBn9lWzkNp1IpWZrX8+UH+tqOHp+YTBJH1sI/Tv2v1
5G9JwxkdXYA3ZbIf/wrAdj78UslvN2V3+1b52tDjwPbHaOv/HeRjV09XWGOnbTTU/HpfS4BDOS5u
y/m0FdZpKOl+PHgDuHG64FvVkUsWULmSkrAvm+5rFEHdqbgC35ohFCdXyxB60A6h4ggADFJRaqQr
MrUXLxn6NEC4MySAOhT9wEevXqZrkagk3chwoxYKWBk88Rof1kYiCdnhkyX2u2VYYym0lnxUBZiK
vc5ilw2WamcjU5cPUsETz/AMyrOZDfk7yNxhYXw625X8r0uyXJVzOrSnhpFFTUOh5xS5OZJ8LA/f
46DZCFnltearSCGms4gYafYPrPvzCGW9rrTPIhh8uEl3PizIbwXynaBJlJZCq0mpwXlx0CxLD2RI
HkMwAt2tT4Kxzu42kUB2fGSQpjQ9VjBx0TRcIZRQcE1KGdyes0iJJJnoRr7L1uZucHXaXE+DZf4+
HlKLn2BjFrUwVNfdYghLmxnkmI26YOKQ90DC2C95qUarV+rN9XLWC5QEE4eMb8DX+DrRDPVcaify
IRw/NkNOFe0m/jy4q6fEjn36SKwEGYtPEdPxUEH/MzE+4I88Wm38RkQYvWGZUi/ipc99gRZSy7wS
4T8jzZxq+9RvHEzSwP8TariPbiQll0SvYpfHWB+JdtUKbr7mKe9Jz1EQGhp8QK87LaDcos2Xz6By
Azpw1FDCwccZZK0lmUZ5DihGAltlcIk9C1lWv+QRONXI/CgXeteyRq/1k3MfTk5d7VRrQ5937nU3
spghfpNJepUQR6D7laFztTFlRhfx6NV4pwqJd9IPIUxqjpAyDU2PQ4mWqkSmBOvUClt9CWChIkQA
/EMkH/TAQ8TIRVElUT/At1Kqpr0r/veoFiL9YsJorBqROHG2JQ3EwF1N2udLpPovX48fxKEnHlQH
isVM+JIZiLC5zZkkMmFBhN4vyJYLcoIBP0JIChIQXcfmAboznMOisfBF6DeuQJg2zRHI5aERyEg2
jvzoGq0VumKAfFm24kFPvtCKBBydTvOQGonMmSSYp5R7BbsRJj0r6GaO1cCbrWnTQtQ/MreqHwKL
VGRR5LWZzBQwkEMZwEFaoMc2iJfYn95jtppkYrEQo0OgbMdYWVwEhhvy/+uhOsMjX2K1NTGjYnlP
vDvWzZQu1HY++fHKiDyCBFGWqm8vA0EqnmlrlhHP8iEJPyxsU/J1e6Mz8MHuSPevbY1f9A/wUF7N
7dWQ8oiU142oKrnkzO51FrWrgpOCHZMS1HEBuu/qIynIsNMACWjeECRoROHy2oL3zC1Vz4Xd98LZ
iemZNy6PwWXoYFe2w2ipqdrTvYDWutVYHl0TvpkWjaviCr5gZe/sghqdY6pfvM8zbeTpMrm5swaa
AAiKU9FEroGi3OPg4+LiLD2KMAWKtE6XPI05LuIEUVtcuG6WnH+nkv6lF8eGoQbrMBIUWgV+e/Ly
Zf2rM5peoACYxtY2LiOLQlnHm9qXJINqmPalTXukMSXTMq+hHX47ykUJGjCxHacv8ZOmdRnam6ez
bEPIpFSt9pHxigbr5U27ARo5Q8gWRFa5eli947Ga8ef6bZNHS1VSvmSe0c4JiZVJ4/UNc/vfeyO3
YaosVjdkRkZZaExB/V4MVbMIkkYTo5Q05qTscvOjHaYIOfhOJzeY4DnCiZ55oSdvxDn+zfJWokDU
5FeAKvgkXi6hsXYKO9YEpx7msPp589ZddsqlIzDckiKnkdJ9M2zv7qKDIstspVCIx8FEGZDGZY92
ctoQHNv6xQ7xhLP+5tgqpv0YVxMlzS9frQ2+qIpzEPFsXSIaQ5P2wkhP0g37GsfdLZL2U85iRHBN
D5tYSW7ND5sgh3ROj0iiGzA3wVNZ0aU2cQN8+DervEQ87lkFlfZZhlcgoJQeMlqbrFnxOjk3YMeA
+X6REyGqh63aXHV0MxLUgos11Mo6K0inYHAB267byNpI2iAcPBgfCw0MbvDjkxNDqO/eUSnynVHO
E/RxzLJbNKWokDys5dKT8krea9mFoOS3K+cIzbOeK6nMURYv0DFMBkQUGhAnEMOcgFOW1gQ6H4Ve
uOTctcrgIU22ZI3bDTELwhXlYuwabtzZcfl2tKrXL8yY0BjWT5oE91z8nHTj/7vjfvd5B/C4i6Ay
wIRg72Di2doG6+FAChlJCVmOEKMzisvxPQiadxjube+q6vy89YcLf18DQ/J1JlzFVQxbEFk0dHGs
3cqZy3C7mcX3exZCPpjSRWJPlvQlQqd9BJlQAT/iJqEw7aozy8rbRpRG8XJZLH1L55Fz8IdZS5ZW
eyG9d9DC0qPecOWMGF3CjE+bRtVbspYS7fqhX4XnO3/ef6iyaAr86nb76br4DTV3+RHmMk9ZiXdE
0pS6iumkwgWgd5l6tb0u5gGHsPU0dReza7VQpQX/QkRbuGeszQz1JsGE+pnUDuLcOOF9gHvTQ65M
vBOomoAMz650gxtrSGft5aA8e9hYmijBoeJ05TVI9eAw4QEbK6Go9ln6xI2XMF+LXyGdEAz6/pJt
HZoqVuRYRD5Y4YQ6y+Otjd469xjschgC86BfKfj9PVYQp5W/Gor2hTvLn9ECtcR2bFhkQ3RGJkTa
O0l6NcW7ZCbY4JjnpszCnSrMrcKxirYg2bPtn79H5YLVsJO00RlbLvRwHP3XhXEbdT+qxYxtXzFf
tYnOWEl7lRpfs6VWxw/VHbDTF6hsR68K2VFro4ReWjHI4kN6794auqKzp/W+6fUySiQQ/xZLPpFH
9lBwDvmy6LJsV51rQ6O3zsnvneXQ8kJUefkQswGrLdBuj+rnFP+MC7C2NvIizyZBZvS/ZtbwEgca
otRXUg1MCXRK3Ro21yRXjGdEURm9+VJP8zgtwoMCZEwg2h33mb2lA4KdAJgjMpfMT6hc2NPvrzC8
deQsN4Z0/M2mpLSf6ITS4IHgD6q2YRMiKeb1lEh7QBZUU8fz3u8hczvPcQiZBY77rpTMs3GmtSt4
ZUdjSDzJ+oIfYlZRgqwQEm/DjzBr5ak9UuRLNKqOtx+IB8MY82peFbIhZebxqq+zpO0IK6tpmJ22
Em3fdFnfjLQkxf092ekiPtGOordJVZB5QvEpkKdmnPdCJEwPM1jYT9mG2ZfIFKruI4KR0nT3LvSX
qxw34VtlKjaJbtx/HAPHrrrpnKHtna5+wqccGt/IBWfpKizrBisWLoqvi5rQlfHr3OXm8gJzOrIC
FLVhGCZZVGY7qfDH/tn4LyVblXarOkJXYb1wkOlywjM7oZ40r4q6lIq9mLWGfpQNbcFvlevdAppp
+kIF6q8NpWsoP3/TDacrM3SEUdwA0AFHWyLqEl8/1DvtXAAZuBg8KvX/eergfP6/maNQ3wJWhN8S
ZnodPJ3Rdi9+zAi0aRU2mroEjXUcdXkK/nuU8fW2/1jbXs1qGuKEvlYgu8LH8umxfR/mo73YXe+x
R2i1yxuu2mopYy2Q1v6/m+FeS5U3YUziF7kpDxxn0cDSB2uPEEc3K2COOcj7qyqwrv4o0vYtvcug
OE1XfqBau/sMcseaCem/HXOKqWTrxUK8uBWlGvOqBUYqjcMJs815hZiKH+7uM1rUWPZCEYQ7RKDB
M4D5JU4CONkkSeSOz6LeuTVjklrDs+GEyVAiURz9lK4v2lrZ4cDtBemGAB6vt8NaPEdaaXTck8SG
iKmBmRTOwN6/L/7Y1RtvarWWAjs2p0Wkxjn9JO+6oSTEnefQoc4pIjL6yxd57W2vsv635KRpxduh
6BclsRQgM1snASvdWZHS7EuAGyuCSNailjFiUi9Mkj+0+W0dwIvMBzbUAReNEZh4geB3l/VumKvA
S0cSkcHXoaK1pUMQZB4BMIGOnS558qpt+zLVG8HCnOExEKEnwiFADEPlYrWZ6mcqHQJSyfpD1oGH
pd2nP+zfeQGas/Rby1Z1WZRrbGw/GJ9d8gPbi44K711+c9qiL/E8Wf/qLwoJ/ThYw1xl7cceJpBc
5ULYZJQsLQHT0PpIstU+rNrNRhB7xBSwVlkS6xf4rh9+2XPXVSa4joPfOkuIHD37cznZ5CrCW4A3
Prf3BvweBkTy/dnPxazoE8fiZTuNO8amTWCsYDNaZnUDqGXb76wyflB25qWyT/H8zI+vQXLz61j8
w1gqIqq2iNHkXHuMmXx12AQ8s+SZHeS/PDQkheOLqUHf1QMuqdCCuIDpK/sdplV/O+uxyFfZST4P
oWGHHp9NOmU+qMNNDKSFGkBaE+hDa9FqSsup/dCMmkyPSyXSc0bSDyBaNxw5Ig4Qqi8a0FJJb9f8
6k8DQIQuwn02CxmftSebFqbYT+4lxwWWIM5abgAsEQRKd/XHrWesCqdhA5JDMsDWYbQjlhHg3vym
bBgI4kv9adY5ChPaZVeV8nlZ26QsF4nHIbs9TXTLKgDSR50UkR6pjLCYaHDHhxIvDouVNfWev8f6
RqKlz9TTe+ThdrEx1EjCTjB4LxpbkM/8v91hmH3/1yMMz6NzapZY65lY66Bg+TcYVwxflt2BGg7/
8AOTYjYyTD1koyUDDshP4Pqgty1CDxSsa2KnqRYeYO/cUEsWz8wNDNlDyNxN7IU+5qkfOnF1w5LE
NsAiuqw1cyQ9ue4h9FqPskPHiXIUQRceZEuEk1Q9Lp6OEYPMjAABjmlA1f0VuNnhUZQYhvAPGOgM
avmfvKVQMg9NPjW8NXBcMDyApgXEsJ2UUmallOJIun65ZMslJZ1Ke67zVaVB/l0n5z4N/9nBjywC
Ax2S/XTqAkpcqskrqkPJXUY4S7Sk76O/TmZWbiIsi+g94gxkOtavXwk4oKr+1BAzi/IlJM79wzc/
Sxadyzj6BieOKJ9qUt0wuFTAevBoL+RYHJCV3zhZBZ8A57EKFeYts0EJrGR4Hs/NdCzozvZX1vJv
lMT0YQBKcWcu8Q4vQwkaGbW47nd8c5QdPda+dl2EQVNjtmL28muq+rpTy0kisY4Bg0lZn23XJ+cX
bFYeuNBzXEoPh3zg4a/+R+dmo8dKN8o/XzD8pUTerqe9x5uXGggk6wHDqvLRsbyqs/RMtb2Vh0dk
QaYTOmbtfbgoouXbDYzJ3AwMHRViRtPnrQKVASdAPXIQfvRcINWzVrDfrEfPSOCsH01fHWMcyfI0
Jq536BMfORwIoWL6aZU1KvkVyj9ul7KDB2+gLdCft3w6Sf+FWrZPkN9kqF8wNO2vlWVoWpf2Lhua
kvSwcenkSg1chxF+N77jI9JXcgkDC/b9d3vY1jTt7rfTqZPlpoZOF0dEjsLFv/I+Rvib/sv8Udmt
SBMxFo7Zkw4TuSh3oibRrGWtahZiy01PGacd4bmgXIKvq6MF/PTsSQVXrRlzomMhd59C5Cj9nZBA
CXKaC6D9ybcW4vjPh+WcuJDn82luTJbnAaBCG5/KSuIV6doEXH7CTomoAoGA9ghEf5SwF82iiGDt
znSmD7KBpq7w+g89N+tmn2Nh11pWO+ejm2XwteF6RBekBFkoTEtg9KqcurAsBfJ4/798OP9xQyoM
cONiSo5YvO07TmnNdLxzvDFtx6oMNXgo+s15tDK5ulEPuCeVm94mAtDgLeA+BHP/Sb+DD+XRf+PN
9js1qqiFuIgP/RHtAReag+OYjCSTf6Nd4LTTe4ye/7JDX55rHeY552sKhRSpYUf4Ycsnf0yEKCRK
WJORaVLSLyjfGHXC8wBAVQB/kdy5Uj1ESFWdu3/2+8Ib/w/FWszdjCD5aQzMBbUQglDm3dQKfLcH
4EHeJSH8JM42uFyXTH/S48Gdm1a3zi4v+8SUAjKVm8qYcr92OSPwgtqEZkKkrfJbBsJbKlpLwGTr
0SIxhC9KEBoMEc21OSZClA4soQA9SgIrM8wWF8L9/Dpi8noGOUb0tbDgBu1Rv+30d2r4zANZJOui
XazRFzcHQeqEBNOXuByaICtJsClgWpM1bDB4jySTz2w769L005v+y9389rDV2lmeSUjPhqb+Ixew
sTg2ZqQQZGHdoaTf7iSnZgleNNnvVVlmpwNVJtlP5W3amZHboJGXpuCbtXeEU1J7stTdxZanlZlf
FMeNXXdplNEUtu/6QtpAgPIlOZf6+l14LXqTEvR1GzWR7soL0lFpSlL8ByKb9Xs1XUSdIrREogam
Sb7JKK08nuGYqgfUM/HVPGLJYvFqKk2R722sj+lXpNQeAaCRVR0cp2fTDnv7q/nMImFlVcI09XpE
Ru3Xw+QxgQiAX1RQ4nHmHAOsnhQyqWDYPU/j8GB90ZJvI37mJNoLLoUTwHEjNL6AEJHoDGQLDEoW
Xe09HmxXLxFUw5jlO/7IfLu6wxCEbBz7oi9LKxSaoDdZEBogDulM4OD0pYHr8lTXYqnma6c4cJ1u
pS+qaFpf0ohj5FxN3TBd6zW2W5rzdhalbfyn+8Ae1jKBKGC4zdXbpe74P+FCnfFouktJfwdbGu5J
bykDHkP+UWCC42MpKGkRjO0eo4G0UGqo6lbvUISZ4neq6KI+Hes6n9YxtK1fuBDlK0ohf4sN0OPc
lP99tCVDlx87u5rgmOGMmcQBXq+W9U93ogUuJKmMdtYu6t8ogQUE3YRXvskGD42BbhfUTtfDO/l4
znd20+IsP7vq9ukz6oma6PwPf3/5/dEznljYd8Pln/O74A/8y3FsOAxZnbL44CVzI2b6u7xKu3D2
l8b/J9ariAMlLqm7eK2PHGCTto371xw8UET0WAtSHgC8Zy5faHp0N5YllAt7V4pQsnO/MSH29gz/
uvQ/WAQ1x5qyX00FYi1X9YpfZjFl4e3gokILlf9aE23WhLdf7cr4dE5Q05P2ORuHZdS4LCb18TsY
0pEr8dPIhq41ytgaNBPumffwfqWsmQXJCOdqNl64qyfJpvLUhwtcc3xVum+NMBpACcQNDf3lp+Y5
jiK611buB5crna/gW6SC3JVa+JexDzymZYBA6/qmdhNmwUSGhwpkjdCngzLp3yn3oZiYxQfzXVBw
R4NC756Evn0b/vIlp0f08VGyck5gDj52Bx2KI/Ez8KeA36YVxOapyu+w5pvY9GycOKoVLIFntqdg
IG7hEQLBN6J3wvbeqKElpRMpZhrIYcurDH1DYAIRwNkzC4sfYkW/Qoiv7pRGm9GRwjBoNOrDCkUw
wxdvacbh2bYiT0EnOXS9BIgYqwD557hlC0LCLzVicUiCP5gnV/eUkM7/WiiDwdfU+5iit9I/GMp6
kmMdeUkZUloCbfFU4IO4MZ4Bz7QrVKfw19EaUmP98yQR73VSPnNK891HJAVneBz63OAnbY1ozVAB
TB2SzUndlzKGDis8J4U08xUrAZf40HLaeQ9+vClMzYtka2c3gjIVjJkmqrod/l3HmoYZcfoKlSg+
Ikc6bpdv0F2vKV7GaKdtCn9ObnjkeThblVRXujO9x4GaoXy5260Ro4N0z96UDK6Sp7tyQaFpV96c
4ejCyMB63Xt7YMuUVyf9JU+Zj3UPqw6IjRFaNHPuDaxzlfUsEokcaofPzaOYMthL2ZokxORGS37V
znseuc6zINkBZ+B25rDBAXyNQuCVcL5D/X41njpBOQHtL0SJctO6ouqXLRj3Qr6Z6+ylM5paiwfG
xEomhrHxfkVE53JYE4KkMBXTA+xgdMDB+z/gu9qi25dT6v/OwSm9lgXz9MX3K6I8nr9R2iyikYXM
QLsCvBq1p5bLz6QZ/GnLCxIROkIKTOZgCKW3iH4Pgz+fhmtRWuwPwUIk01Ribf9YG+Sw17aqetIG
NvI0swxx4L2a5BgsO8QWDwzvXdJRiqTZZbteQfUaHaB4TrE/LcMWq3mI3fiIQg14YrH6oC6K0hVG
rikysiJaqLGjCNtTnMOLSHwUDvl6QHkUV1RKFmWS7z5rYbAfOSc6Vpp3pdayoD9DNECj7dN8bvvQ
JTizWpPxXN4zrJt8J774TPzQPy8/s1ATR2hvpp5e0x821sAeAp/2ayns9rxLDWCKkAd4K2Vdk6Is
t3/OL1EF/RXojc91ERFW18XdVDTMjTt3BU7g0Cq05iASoOSx2djdVpzeMPVBEEdOvIF8kY+4Bdza
Gby2gb9HKQFQfzfrur2vnOlpj27hAa1X+mVylZULpcyBh+FBmdfHf0zuckQ7nIq0UodVmIvv78GS
QUZfPAig5/Ea4+ILY1/oKgJHzB99IGKX3ECOdbhIBSksrP9gpsNLR/HiBDYxpvdj8Cmz9Z9yE1ir
hViqfQ9lGHNoCuzjpxuTxUzJxzgGquUtwUIvpZvORXI4O/hTOIxQJHX0otiYhTDSMP/anoGbJsFV
QSlC1YM/+6JEOf4pUZo8dI4vuKwvHjetMQTOvtioUW9caNSSrdku3Dt5i5D5GgRBPTVTOeh5Q64t
CiVJSb2EZU8XK+c2vq6pTpTApn1l3wHPoj9NoNMMliQm15Yz8mn3abEFSmXad0U64vtctApTt8fW
CG5DtixfQUuuclWpvOKW26y6ADuY8MKDNpGfuZMyl6262YfjkNV0HwrKC6xgzI4WJsE7B+5ofAni
cGY4sX63gYau7bBNWMBC8+jPWdp0lo01v6Ygaza8xIrkLz0DqRfr+I8ZuyM+XpRiUwpmYxJuYfeL
8VtQ6jW+OeRIdBg/zc2j7xhxRr/llD6hRtHvMZu8RKGRlDXRG5kx8hlW/79oI0ssIaqDNVPwqsTr
FiCVucPthkAS9+2VkCFoZ2vFAeYx9ODR5gZ6FDhCb1MIwSLXww3G9KSPDNwOy8wCaGVbqITnGdT1
uiU68GEnnQRIKQYQ9HKD5cIioxsG3l79WE/tBc3RAjY7oVZ5EJwiHQViV6uEFA6GwjenOSgMGZaW
qsyS5rNIalxqDYGEWQSFZLIARjdOGdDAddTdxg+avDVyUMwd8SNZSB00SVK/lOqHbfBtwL7y3TMI
NIO2jHmxGtsLUdIkWud8BAIlnrmidxPuDcx/WykGYNfi/1XluuP1uWgrAHoJ+SmgTJ4ruWgBzjwh
UcVooMVTO2G5fhE21ZNZlwtM5Op5lgqRkbjZYp6zqdZ+9wNmk9GF6/X/F/pQOCAgqazReDNqCQHm
Q/PEy1wOY/u/vfRATjS5lutgaH/ixLRoKmD9Yuj+qvTFkkeDCzoROnlFrySIUbcTVd9PP0vV1fBL
JmpvKxoIOEtLXibFiMZ+gZ5pWwwG+rvgD+wxSidSNWyrisi3buK1YHmkTxFojJwWxjpi9TKxxgPR
+wnOm6zKbMrDvsOcueOHR3Puow0hsYFsRuTScHitnzMIhGLUyQqUUT70LAjZJKG3PtijihUSsn8V
unjnsoNn4uy6N0/qoKjZGKe1dAJKbHnGdBNRsVZNKqMzNYDHl5ebeY5y6udVEkAN0VyyhULW1lEk
2/Gp1JaxTka7aeXN2z1BkOzz7cwKNbsYpxtGl95Y8m7MPmo8k2QF4aew3EHuN/9UygCjUh6eRETK
tnbd47tvoEV8ghQ1sNe/DfttSmpOmjv1YmuTS44ICef4bz1GLCBFymtYl+GOFnqtXf7jqIEplGT0
8YmciCIp5RJL5zeixZld6Ynr95ZB7xXhkAISZ3NWtJD1Pd+kXHY6MEYJQxtLy2T/YdV2aVBod2hF
FRyqipBVawxPHeprdEfBlOBFYkJI3Zt2cwRWmj6rO5ry7C0HTPuTmU3h2rP+OzPRN6dwIRoGYDxN
oHSj53eOZJpSrQTp7ffr1519t/SQJReFAmYUCNFMFFycwapZrKXvOi0jdsN9HiubGB77aiUnIaAR
BYstK36I8WAW+liY2pl6zynJqF+Hudzc6R5wGEJrnf+cGEnGB3VyznTyZAKi+TWKALzqhydn41HC
vP2pCjB7pzEfPAQqqpIID8O+nYcgugbKQu9NquQGj3dNCZlc/YDGRTr0IkQyvrDzS/Zf2b2kt7Q+
UoyestHpMsEqsBrwYWBKTS/QpOqfla5MtQiJMf7gvHIGUWQ8J1GofhniKsKTezK5A+XgiKl33/Yk
VXfJpJnlWYcw/CwbnYwAqdIttA8Xa7vJfWonM0CBSfiB+oz6ynYTPpveApDHrSq03tElzQhHqkl+
TvZ0rHwjTQbDJ/gaCfp86RatfU3iF7PqEyMgOA5eT/5FxmC0Q5sjnZNAkD/4dFmPlXWQ8g0N9Q0P
dPtto1XUUdDFC112niR6EnXrDYHVdFejdazvlNhVtmxjZGK8Eus4DawdPL2o1cY0eprqwFp5TuN8
XfMAncGXi9M0wSOrJ49klYJNTP3UBDSDL42ZF7c1T3NbuRMfIM6Bl7N4pvaBdfPWDxt7V2OOexI+
A6yEloY+wLlnXtFs1ebSJrjZsLfAr2Vaii+i7SMGkI59hnYLFP0M1t3XgwtRlUQNzcqtKcbBfyyS
WUJ5dnwj6zw4lV5kg+LfZKKf0tGNpchMHJx8psI/9/LMkun39K+n/novXb8jWYhJLC+c00ZOrMoc
qKcnlYyNoOigEcfNp9yXrEl40lsj7aahCk2F4hmFqhB9kHovIsuuQgJ2Q9uwNqz1jroB4O5bsqCq
6RJFVfKOxYWxFc6278QFAX4WdvGYxsq1vVAJhb6Bf520MO8H2X9MbDbA8SQ1mExEJZs/70DIbD1D
9cKKIg2dvKh74BmaF64ZXIAypJXZKSA3em8cUquTVRPoLT0+4Nb1yLSAhRxYABWrndzZOgnpvSw3
tcDcDZtyPU7rccIU2JAQ47i51COucHyT1fu5cFvhtVQzmFZXg/Y4IS0I7xZxPiLoojfFoznN3wt9
vEtEowvwygdDHEDTm9COGJG6lm4HEHBm+P7EbIHPATRHhtl8fqgkrB1LSAF/+VXPCW+JnXFViO1r
AM5yOEZEux64/bMEjhXMcgRBL6vkNqdvR6BCgp29ZByhaWi/6d4vrvQGoO/1YpkL/gFdrjzZfgEB
Q5niL3w51gPUhwwqlpT6dGc33OmhdEVnDLTt27SZz0m6YCJ34s4Ij9NTYKf8ROLVtyX0+UEJR5Ow
Eq4Yy3J/AtODPFnkJkp7nCGwV/WjgGCfZRC4xSRJS46eWNIPRcLR+VImg/MldjF9t5+ex7c9CzPs
iVuEhMkYzrtRyWW7PNanYug9/3lSSTM0/M6HtGbhRQoyizIUCjl9kW+o6ZLFKXhT5nnTRIseY6bC
4hZiVvLX4KL/Dx4P5ENaVYx0VzqmFzYCoJk87ICSN1lyrY5iTaLNAhfREy72CvOT88MxlmSHQnFk
lcyf+MjQMXqKFMOrluZb9iDB9MJEsUS3B8CSnru/x+Kl8Jo1yYhvjsEnPUVWMP3UF6+SwwLibXb+
NCnxglQ9BxapIVDeWQx8OK/maE0OlV0zKRWlrfKeU7aZx3nO9P9eJveQcEVQJ6LTK7qBFldQbwBm
u1moqRiz/Yodl2XZZzq64kbiRqfFjrM47Gui38PR2lR0LoBxniiMZf+LTM2tsv7rpTbxQJpwvYvJ
fNygul7OqiqLBcZslQNC1b/zYaQpcBNiu23vh81dgQxU5Z1/dJTLfJxHHGse2golVTaMTNYRaFNV
uV7M7m3NFTOAVlz7pyiiG63JMJnm3vs1mfRaoFl8aDLtMCrg7MMDEjHPnTxX0PR6DvVXQaJ3KwAP
mJ3BqLlUDdX0Fcar/yh1keRQlDtBSL28T7o48+fKCdkJfFVmv/BbWSS476LEj2GVvYZnhyCqDIWj
9So+bUSgY3SgrrZsGNo05aAedVIGyxmbXaL63f7Ywpma09lU/rn6Q+U7eZvAHrIrTVowB07FSP7Z
4HyDOJZZazZOKTXSVw73+yFkkEnZNVS04LedZifgipvnz546cArIXmYAY6xLCB0JirxXi6lRU+dd
RW72B/JJWk+hxqCae3R8mQE5QL0+glJgSEGBhP5gaD6K4BoJwoLcNYpleXb3ltmhTk0ZsYC+y9oU
rZrkbAZ8cbr4SnUF0vPQ8uF2gJklRJKDBna+TLS3+tq8ol5wrcZrJEKxRfCcPaypRrLN9ZPSG3BP
GGD8HovT9q5T0h7PmIf3BSCC917gvoEQFj1TdUm8RWaS3VL+gcz5pnufp6MNg9AiWwUav4yrwA8f
N+8HjVp5QbaN0eTW/bMg/u73MQOmye4YOAkWrpQv4w+Kfr33K6WcgSbQiLueB9vCX4U/Prt/NMoT
2fKo63HUmTAmtFAf9hJP1HlqY574Y+j9WJDMQdrms6oLgyFGRvQTvzniIsKvdmde4P3jThxnn/40
z5UI8YfGUQGozarImMakIZ4uiMB4C2cS6Mq9Y1/sEy+CSOdyYzZ0czkaA5eT8M3EMgxZ9pfztbDX
1+f1BDW+cf9fSh2d3UVFwzsI2fF3zGeE6M4XdXSHJKpvqadrao3aGldbJUnaqKJ4apUUFWsA9SPM
oKuh01RqYitQ9RA7PLyGtYCksFphzlXIpecfuoGZvzZ6ZPI5EJRgvYo+AuNZr3mtKXbZmr5cG2AX
PA8DxXkVcQTaESFRMjM176mPp3iBpOGQKxi4Dhj7qEGmIjIk6cJRPcHDFSyj5Q0r+oAcNMDukHy1
Dr57KttwwOpYQKYZlwRYGJxNoUIIeOH1b1VmPRhO4CXc+d3aKTYFO+ZmtQadKtnYpPVsFQyKz6Wr
mzG0URxxFn4KQB8zpBUId/afTX8ABRQHINPYsvLhQ7x6EportUVXXkwmVHYge/CIzN4gyeZG6tuF
aqFIv+LIb4LTRfVAGZZcRPYLcw11wcOyyvTdzJ5UMYnVKL/F4nC3Tl9ypTqcmIJjIythmzxOUzbm
WWKj68uofNclGvt1T6ik7Ki3ZiO5/OykB2g70MKxZsgWb1YfgOAr8evO9U5wfuM2sSpq9nI/Trq3
UtSrznKyM1ajANeduPTsCCVgfwercI3Bmjqe7+Jp8x3Av5caUr2UhvTCvI6L3gXcAw4il+o2o60w
BkdEodmhFjIgkvfjKr2NS8Cgkg4hz/bhhpnWAcFAzE6RLoBl/82ugokD2ht9MBABa1SzC8CllPsP
eBRxGcNqCmFNIArEmlqEuL9AUAOgHs6M7DfIRcm841xmjH60GttAFcTP2JS8hM+vLoejivsma4Xj
AVRZ42bwL9xQJIJtBQw+DAB7oNr65rinWDGB48xB6Aab1yy16B3+sLs84VkSxnthvsiO1Q8jwtaL
AYXMy2Ab3oLM2ZPyocfiVSF+3y8yk2ADS60YO6Dk5SgEsGnFlefPThUtrMKktb7Pei5ZexY8GKsK
pbYqCOWjTcX5AcoJD93qcutf1um7LEU3kEc5QBm0vcXKR0ET54Jxi84jd3FzgfvyA8I1Y1Skrj+s
sz+JNVLciNEHAX15lrTG7Uf6lAscA0xk8mGjuVGPH/Qfw/Rq+Gw1/A5bIC58VTBCWSEQbg11lBAR
1sRKfGOipZbqcqNMB8iDfZlP9wIVHeqG5AnoEoIBcztqtzDa4aH/NSqyRXEsB9AkQYx4xh10aLZT
Qcnc8OcA+V2VCjrRjepVZKFUuEnSd7oXjO0wLWFcD7pO0avz1J2H+qRVUNSygoT+23Fk9ujoyG4i
2VO8uZo0DhWXcoo0Zkp8bGOovnyjWLAkyVnb4ljWnmWSy828P0j0MPZZ7+3SGR0rtdU3mlj1vF6Q
MWaknDQ3pRw+07U/+q+NrLUYibhRCshjd/39s4TlqyZIT8nYUCfRrT0cB5vy3pSHCeu48rjNXHEg
I96oS9ENnT0MSy6APpzl6EPJj9fayPxa7lHFltsMbSNwysqWjpYNnHJtrqCJYNfoMMx4uTqbpE5/
/p/DmM2WqGkTs764AWgWGeWKTytauv8dCSsHce2qBK77VAgkMjmfr0OBfJA84WT/SwpwBDXLWDD8
9TExc0iym67ksHVDr5gzFeCmjcdssIs4J8bVfaDAMekyO/9NmWDt16rbYnpmJr/rNep4ck32HWgK
Ag6LBl2SP+XFlG1M3XmZmOU2lQAIXX2PwuuAhQiXgxeU4Kys3O01Yy5q7a+FOa/kN+Kg+/GLd3gN
/W6ncH0Zs93LhpnxJfqMsMJxAp4OItasIrt7ve7Lj2NR5uJN3gu9spmN4GwwAmxT1hbc0ZDabR66
V740ysBED8EPYXLZszQUjV7LF1FDtspJjJesJ0VEYPWFbdjMZt0CovlhmD7QXHOFcpgCZFl4mutc
beqiigFLBsAO23o2oAJEecea+lQHcfdq96SyCxvic3ODEWzZNGacatQ2zuMp+2vC9oEY6fJWwLkJ
s+XYmODxYIPM3UwNKqZVjSlQ7khrMSg4OVDpJt5QxBOnTR2ePxfxpWUf953qo9Wb8W+ygefjNMnN
8ZSJd33kiUiIAMB1FkNQJrrfRNMQEsn1vHIvR2mcqZJABf+demsZX/SeC34u/kdBslvsgRSdstBQ
QuMuDj9ylU77Z0BiuiUlVNBRQS3MTuRhxDfRiQSfF/Hyq8xxjYFhZ6xQtXKp9cdr0HRS+GnVVrlE
ovT77f6uzwkEWBlTKkpMA1RZVWsc3hdXSMNJzl+kO0UpHEOhBstKSxLfe/gXiPRpR+Lb6mvD2bXd
o/fhOEm+z5umt16X65cYxrk0khIS1AAzh7pfFYkQ8vLP9nCIVXCOTVftAOlgYbUCdmhNrhSLuARJ
YmVGcES9xpVUnyo7kqdR4YZ5Yj0+sGKB0eJi+CWLLcuw9bgertgRWSkLVD+10KI7sL7WDh76uFXR
RRRFy9hEx1Lvz2myKl/luNIUxVQjMwqNvBYfmG0Sd1sXrYayaXrhTg5XJySupf2RDe/PMcOtE2Lk
bcV97/K7DLY5b3gxnqh1zH34/w89jtHSl0GlU/JeocdDaCSZkyhEXOGsUmuaumwY5HE8RrINi4DN
7kEKB0CLw2n8RvNldL1vcOoWteH2aNev2pNyLDvMKZLWqUk+rFHbfFKRgcB/DyuKaZ4OjoGssEV0
qx9nbIqwgAXm7o+i6OcbhEJ+3ZY0KoypVTV9UHUGJ6rjfi5StSuiDr34b5Rgasl+7y9xNvMwtkiY
goKaLirYARshITOSuV03bnGeppsOEixwuiJvXTNjlEwCsOAmTih4TG1z/7JnKEU75k+KKvP2ICd8
0iV2W5fRFFN5tgTuMDiKkaK4kvo4OPz0vk1aLtvLJAbAyj9aMK7kY6A6xu1Nrw52BwDd9LBfF+6s
/PnHThgwDuKskxScNV85exVp6RIZr16obdAgGBJ0wWAdy5p+Ccy7LEuvLLsmbEyEdbndEWcAJPFo
EUjDvxRuC0aNMwZ0MUv9rn9he4m9V4iHSdmgDDsRnXr3gJ6W0JGpzybuVOv6rWc+EpecrtrIAyoc
fdnsjII8mRWzwNFrMc/d0dLYu4+HelWqCr4MBZ6nh06cO23M8or4ZQZs/pNY3ScaASXJk0xIJKIk
I0GznIg97tFFmDPqb8j6r6BAjluLaKsSGhH8UBQBdAt0cmIVJ1/eBwVOtDEaDsHjo3OAIoVIHPOq
jxSdq16zfUq8H502hxAadHL4B4HxEDl8N9F+uOBX0OTt09Va/GS5fOGq8nv1TqlY8W1GUqgCoFsc
4iL15GBWBwVIXU/D1T/QRJBGu9wPs3yNpBSms772mlNd4mnUXnWkpzN7Hqt9vRjYIIF2x/LKwcZx
1kYVMnt/jAIX+/EiVVNzCTuAUEj/mPq9fkS0OBg3vpdMVTW/xRaQXK56fXblKDAc86PXaMq9kaAC
wgYKqOD1K3oyee3euy+Q42TnFEZIvvQTiOk3cKdr5ILWDkSmk/kT9lh1JioeJfHK/GiMg2dYnXOO
o/eLUZzBXchsDfd18xbX3EMe+o8EvXJ59KlnznX+5s2Y6LYxwiyXipXwSeBhIfBMk3Q5u9l9TZOl
Dc20aFzPOBvnWCkox5/YBKroyaY6Gk0YDO7KM5LMPy+B62KtP3xcqSte3q2dhTIJGh7LuSUuyzFW
LzVheInVZg7jp4mzlBi14ac0lTrk6DKX9f+1kXrtzdzxGj6eOsh/+NP92fqnsEfpPLIJmEZl0vnm
Km7qYYx9a/Ws/0tpZg+59/bYgFyIh1IT9pM2/VjgPVcmAt1RrtoJNasLgWZztlJM49XLzhl+ixTU
H5og1mo4vsLxfFi5FYiuh3H97LKoC4aWWeak0dfaqjScAfR8070ptNnswyt3+sbbBJFWWN+L7Fv0
gHrqgsITHPWXS+XaZ+6Vzy5y94DpGC4YZrtlznzLUvaybLY/asDigIDrEGeiIBOfcOqYN3VuWj5N
4WLMimijQlDFFLkBWghdyfE9GgrH+MHeVXwjnyr/anx1RCj/GnfI8GLzzYl5Z6H0KFGgnwOZoSZm
M5APJl0eXwz7LHyjEW2O97uHVJimY9BorVnizYFKYc1NUBFr/Lsr4Zc8w/JNr6eKnfkjP4zfvziI
NVnZwASkbDt9mc1yIltGBg24djEA3TDlbx4cB9n1u0l81pUM3nMRsWc39uA6Tw96ZoPzBRxWGDLn
rzp4YRrqfvBAMgQZoD6+AwzxQf/YkLHNS/cMqVlCIuVt8QOZj9tBYmNwfOxTqrHgAuQJ0lsDrlrM
fDYywsInivvBCyS+67jlKgBuGsp0wNlCOXILQSXIW+wUw/gev6hLUDmfWy66y0y1tbj0VoWYvtw/
1+Cr8xvuk57MgJ3ZzFbDA4yyC2dmedHXwg/I7BRDFz2GKCH0RcwPbIxCu5XQZfV3kmQ/DttTkrU8
8QzRRfRUyl3uByQPaOvuNWYnPwy3rhHbaxk6HIGUhyzGzI0hvcaYg/bx/ih8twW37NWd/jQX70kz
mo1l2NtVk+k+lYxguGL++j+uwGbV6V1gNTctSeMzLDxYbF8ULiopROhz/hyoCWOqMIijmK0cYHjM
odxKvi2sQACTAhgncjPaUk2SbdA8ErTFdFs703JSRfBUZnCQaGwwValCOm13cTfpYQbUMdiV6RlH
8TiQ/p+fTa2nSYbBWKlXwPMoNLgce6opJR6IEY/qZq2n0He0myuYuDvwAjiuOYJ6TNK9i+bjCy8c
/D1G1weuOUwY1fZq8MaMNFrY9xGmDG4PGO9plW/D2lbkB550WqeWpipRFAVPFt+1QvEUQ46DaoNS
hfejwgf+KjEZkRZTivDtd4YCcAQlVbX2i97ixcwOWHJl8Aymk6lQ/bWCJyRQRMMxaTND67E/tqz4
q7zOwcdtRkD1hWuqYSEPzpPFDaltlv8j3olJxNrB4tXjEbv3Po9Ap+kce67FfG8W69mPUBFawOWS
T0gvaOoAS1DMkVcAD/tNWEcfJJKujw/+jQ+PyRso5NfGeBgzLjqetZTuSZ0P7Tp3UrE80tmelzFk
1pF7Pwlixk99VVJa596J6USHGp2JL8cj3dpRDuSG6Ib0qEY64zG7uEYFipyag8MfOab9t6ySh7Sc
Bq4ysSpHLWYll+dC546ZVimelPRrErAbXVb2OfkLRIeSiCroTLhVVOYjjdjS5B52vfLrJJ/XyTuX
nEKHPGnKnEh6ZHQvTNGuioPyU1mK/o5sLO3VAlVB8jnQeMAFb9Ct9V8SXI+L9v1X4T3UjXDbXcJg
7NdpEKvs1AvDrXWrCbn79aZ0C41kF749VF+RI3F/18Amm+ct9+lkxIfCtflhhmhyVa+Y8WRHdocV
lwqY92IEoKZGDUYsqAXetzN1yarJy1mkMT7Q5Z14ge7oR6rKthzUqmrzCeqSdCKRkiKvS9L5MEf1
ZAv/yUhUoWiSWqC9N13cu7uBPlJoG4DckJ3VsUEPq3pjDzpwMrx4qQK18s2awj1TRtb4/GdUUObf
+U5Ly28/gQSTmUNrTrGT2LeogvhWDv0ZBhGZ6DCHg41dQDHQWlIFxHwYvHWHY+p+zOCtrZ7eskuB
cR0zOaC2Mp9qmfbcm+l+iFncjloNfZrapJ4Whg7pkL+LDsiTClH+S6xyCCC3SoTFyNzGQQbe0vm3
g9rF5hTZZdiGKNZ+mb5/89nxfmReOZ2chy3W6T8pPhzWAbuX8hk4yUfcfA2R/Rc0Jvd9ZVDz/vJf
qvNZ4BT8RDpuRb8QbVF2dtwvsfvgqKnjppBmBbLpyBzTy792GDTMnN/kwYpR7FWshRnL5Lbs9d4/
/GEgmNdAu+qF8sjG0Fc5i7mTBN4B0FHOvcQcT2C3or3O/I15p3lyXHUiXLvWV9AOb7WJ1mvAPyQI
cvkezyLTgQPr5hbtSJkQRKHGu01G7tUEWht3fvFLNXdfzkXD2Exqo3rxaTWsZl3D3zm+grkJBpw2
B+kRXcss0GsxfQjCWVeh3Qu2hgjCrgpZme5p3BgCuUqY+iw3P7o7ID1c0AEqdNJltZpXgj7m7fT8
q1r9v87l162id7rEs6nNH05NHz3FkljrVlYh/wBnIP9d1lkcB8grdEd7NgvFt7wmGYNmZo10cjnk
s8YBfWp8M8l6dlpUyNZMiC/TgacmHdaDPOdpAwi1pp7M62+YF3EeGiiDRI1u/iao6FWg0p2hSw/d
FDLrnxurj9L+O4ejNdoUxS321cw2CgM2gR+UfHJmDzSnUNzz+efIqAOyE3A/C4LC4yJudN41YmFB
T+4yiC2bkF3f2+REhcUHGuH5OdWk5pnbXL6gy1dPOxTfM3hgcevfTXYIlfO0FiQGTIm8Qc8KDr/R
fasHGFxM/p/UgesqjWUIOhQVg/+TaRPVs3oU69wo5rCsrQI3p5JxRg9ReWG3N4eIZJj4be857SH2
28tMs6MLyIbA2KcsvoQbc9lwc3+SR95u65eBXB32QicYbkLsq5kQaEDwuCaGL8/ouL12ObZa5LKw
UQFErqWr4A9nM0a3vEZhUCgoBr00Ze36SHnTo0SsXBUduHfgf9HaD28X4PwIsnU4eb+nksGTgef2
4On02cKrxXPNGCB7M9RO57wwwDtpAJg8ecrYcvs9fvYpl88dSoXcWCAbKaYFY132HGGargUMsEV4
/5O36FAoBjSZHMOgtBdn3YlsuUnqtF84LdIl9XbCijlDG5MwViMw6QdMbV6c2yam2rT0fZiOnHmW
HzFcl2noZOh+xMTzwd+l9JI/bN1nEyk7CRfLvOJAJ/RQq95lA4Afo5quThYbNvo2iE6ZYrsKgoVI
qzYwjCGkBuHefSFu/M3c1CHXrUBrg8YUcxNcLIdlHyPDnOA6k/LbidXVna1GBS1M9AJC8v5ihzxn
Mg9FW7X/bA1K1cChp86GSaHYIC89pvflLV7AmBjU4oWtTUiG+FI+vbv5Jz9s33L+VGrVI/Tpz1Fg
uZSr4IFqzG2gy1OgK7eDyrINWaeJXKIeyfuIMEH+gGANd9Oub1BvFa9+qe/WqR7UqnaM4BeoxG+0
q7c/peLPP96rv7urn55rGjivJo8gjJr/OcUZeFfHqYm6/qEI3Ghh++DGX4hRvcSYRNYHPaR0gTOX
2J+p9a6CW5T/c8s1Gztn4fNqKBtnJaMKOrFYu/80Y0zSqN6C0By0OKfaaoaEWVRrUIdJA7lXZEMG
VXcfp06hEDPLqwxy2Vg14koljme3GdQAtVvm8YSJXbEbLLpVgGdQUMBthfx9IvthyTjDq3kr+FxY
mI61tXiV7dyEXaX0adqfdIlDuJxayEoQK8HX1+8/u5TM7BJ1BQxU1c+1iymzeZoc+iV31BtZmOhp
xm2+hPllW5NsS4j9SQ3w3r1HyMctyBpkDqeXWbL/Zfxqs65SlT85XY2wd+oXdCHTD16G94iIxPm/
1nd0wMccSKEcgEoPrUJwVVtxeqGuwlprDieKkvlWOHZRa+NLdzXUgBkYCFit6m6eEqQ9sqDICVdF
M4q/G3ttpyiVINLITBz0uMZLaYLusfQ87a6VH5WycUDrcacchKWg8+JZkTVwdIORFrfJi9J9jiY0
K+4HAPfskUDpJySbv7KWT1fWa2eqXVW1ymzTpHuLebn49zk6Dt9t5sNspU4TgNfgtiVHCOR6Pj2l
n9gH9iOpbTYml5kkM5/xYLjWMsevIG2b1tQHpFiy8A/C42KPSXp5IdhMF6aLLIJbuB5BOyJRaCi5
MhdUe1jBO/1KWqM6dXMXWy0u1ww7J41MxRCCcOFhmaIGRdilz0Q86dMgjUHsKGuUcAZXRj8JO3P1
i7KKqRQ9kQDsV8V0I5Krau1PRqgonaC/L+dRj9f/mZqRlNpN1nVsBJEjMi11+67wgVa3/c62Vu60
CYDv3bg7c15zTsPAhVM/CWD+tnLpKl6NPyVKbWTPLBmy9pogWhOa+EBJh4yzI7c5Os/tkgzR8C9z
QPJSUQum32o78zN+CEQVUG0vE2BWc5qAD0E71wSygaEWi2KMewKoTAJ+PuMvCI6tJyczWfP3jlsd
dO+mN/+WiqxJIM5SrHqwfrLewzFK2KMqTBrAtthSIay3RhtyRfdF0DQPq55MhHSsC9yZg8R3BRf7
qeKLDnX07e4iAwz2MVgS6iFHtXE+BWdqjQ0eLM77q0iZB7F8ckKAPp9DxeCM6aHs9YO9TvBRunpJ
mb7T+YpVIlVpsKgCwZnUUjN0JigOoJo5QOVuKt24ZBOCThrvDRPiUQafxbW/pLHCj/e7K0Vcjeu+
UuMmFsI+bOgtrL53b5ShVGZ7z8415+4S2s/wjL9Jbo9EDtE75MNjwYRcmOqSfov8O9au7qncU14S
gHENIJQbkI+IwS1jPMzAD5JL7M8CMle9MeDTCIUnTadz4vWXZZ02l3Q/9FnY77c+iQmYPmLlTOwa
Pz9TwFoLFz8h7Vtp+CvHH74JULjUVrN1Yd9ny16vignrkcfyq/E2TR6KQoEahOOy+5X0gjyuXt0G
bLRp3yGbrjShHlLA3vX284l/L+aIf58CyroYADtA7ZZHRTesvcdHKG3xrPEbAKx//aw3BXwE42xy
sRYQ/lfF2UGTxnLOONf5sAk0GC6Vs6wFdbWkNR1Y7WiOCMlreDsAIXoA2dxpCJ4aSZ5yl92mqJXq
LjR17pjHshEW7RCB/mtJR/vCNmH63WxaXBoHrGukdyn85nkdI5l0pYgYpGMCQSU9QhQxLdUgpgGl
j60eQFpO0dgb00O0O3JJJfzrVQkwT/nRFMSoH64Elk+70RV5TE/nj3ShNmydhg8WCr3BpchwwmxS
WkLnilAqXQbAIP2qJjY2SBqbY7EkcXzeURSrAMWcb2/KLThdCSfYVvtJCRvNc7EFNi9iSoXvkSbO
atC9jUDkS93IU8mkX894X1rItLP1qaSyUQC8CwwciSxk7w/o3Baj7L0tc4AsbqHSj7/kFsTsavNP
nY11994SPFiMEoplgE21QGFd0hLzQ3sD5F4AN1zOCE1aa1Vf3yuNON+aYoZQSPjtJqiWJL5BNw/F
xMLl7DRFnLOVfsXIHVRAqbMB4FRIBTASWvAUJ6hCqUb4PoDuzMdCTB3MTHOB0jA+OGoswTpgflBa
2qgbc3g4S7LyIjA6yz9POXJqX3avfmvG3A4azx0IRNhd/f+gA1peNbpy79tostjx4l6JpQWEfK3W
P+WrwLGIsJlma8Va1DnkTqcnzlf14u1vcBS08LAYRNqkBbQZqVLzrUW8J/Ozo5tp1DH7mqoTPppz
+/BRDhpIasorjpO3B2yg5JfsIBp07PRkRpqs13zun/2eq++Ap7sA6wKY2vSk7wfWpVvixTLJhtNG
XaV/bsNF5bREO1J/LU3kEYePn3DeEzvW2T6o/QnN2xnxVBO1stizfQkZ/NRd/rm2HRTNp2HqzNOH
ZgYVwy0mOj8WWrhBaKy41vYO5eg+pLLNQxt5WuKA3WeePmlni4D0EZLevk8Ya0CwdW/oze5Xg0Pn
GjoH8pVMhQ15NjpprXsL2KRc5QbphPRUT/q4Xujdo5xW3vWXgdnHjZDhNq3K3TpIQ14kQv9JWG/w
gtvzDrM1fbGhQqyfhRHEldPMtCYQtK260nYGdHLcdv/d7+28SmKvHU8uAV5BesQ2lNUGx3VW3Xgh
pkpQx7sI1P1YMK93HfssHzYeq7kmJaElxGn7xvY+oEN252gjcd4o0eASh5Q5F8SB+dF20pv5RtHi
YL2UbGqQDdNlsGqgsY2F0cEt6lS/9z6Lb6lZvvL3Fzreo1bXJEAzN1Z8YxzZQ5Hy7Tw+25BZdpHY
X+UmbVCDNFXGA14gqWh7BJQ0+YWH3gp8x1X3GLsZPHfcuhZQK4KHVQbUEy/56CJo1HwJbCbdqIbq
Rn4nwvAOg47tsTUa9ql8+BdFoEsNv3EPCiwefIdKzLNijzNSZWjA3+OpnKCpNKzp2rlP0Pa3lZac
IzpF8Hs4LYKNJqSj33thXEqOJCjh0YNls8deyaz2/HrL3M4bvT3+6ehrxjuh4Q+CH+gmvTpgqDSM
21sJPnAftwZdJN13saD2tG6O5y0xBKr72qVGCyO8qySCOmhFhCw3aP+uto42gAjaTq0N8KMtmJ66
tDrXqh+RdPZourgB7pTJRAKZNd3FstvZ79uNqFAEvVDANFYVnggJmtB9I8rBZqZRBOR41SV6aOHg
JlmrmQxeVjRXtGsIeSjOh5aTjgbIBcp37f5mvhsu9zyt3rM3iFzpap3hRU1o+YFMIFFrUtCDiS7E
WKt/MXD4PMS3tqBvnnklfXVBy/RmI06UPj3MsUNlbDvhUbuuX+MSf5NuOTc9yZQCDM1osvY+Mryt
/xoeXj+Inr8GU5jeURtEuPEaIro2xliXDd7lfMQsWfuwUaY4w+22k5O400F7bc9s9OKCEGQnEzwF
yn5tC0KHS/Y5wQ4rnXteJkyL7OTt7LLlQYRJFTkRwW/iA9d7+IGI1uVVz2O0lI8uNx6BUZwoRZnH
zSBfS6oxKD4Zjvn7hBV3emtalqMJAuDtEK6oxHDiChQ7I988Z2yMigfAuu17wHou4sqZ3WUYBjWo
EmSmWMYZcODCr53yBNtHjq9I5pQrZsi8b+sBG1G7IJUcGWJ3QtcoZIgOqDu0/BewsPgGjSkL0a9E
E/DHluLw3uZfu+kFIQ4ZsdVJEZN/UTkGAJUFHVqNmB/5hzrAGY0HkZcxi8yOyOce64bs1+u4touB
D/8IHlrfcPZXzgrLzYZyC13rBrEbvqbMi7frAo/B0jNzg2lkDllHDl2mmEH0X/DF4aRJtUshgZcF
cbJWkhauFrO5TYwgwL1SiuWgPB9zUQP2n6P2O/JGCJL1G4BSHW3VFbYZ+bo3KqzLJXyyoFdyK1CX
gJsbeG7POmI4+cr969rENXAJY/jlQVdh/oQTgJ0FE6g7d5CZX6gbtNPbbH4ZXxJbLW5jsGg4+ufb
YVLIYixAwxBHRfYYAV6uui3eRlWk8P1tyeUwhZbV5pTPfsZwoN5ddlNYShYS10SxN4HoLaYbLMwZ
kwZwAebkMwPgIXtHdxHc1r6/m1vLsNGeXFh8jz7osJinWq1s4d5q7bYKY6yr08SxTZSUua/MFzrm
tT4TTyfufZl6ocpzxl3YLig2vLmbb4qbS3gCgLLDAyGZQSMyUrOT+l9PZbu2QMce7E36Jfnxue+x
jROOKyx0iuHBAq/pTn7tudbyRQrAT6KKa527mC9Q9bTKSbe7AchMj/yUq0R2b819E0KRLCzQgghA
vM5VUaRHN703VUPj7Sh0D5RgAL+uQq88V0kyy0y76cBjNDCdkREMxXcqwz/Fyw+Oto5etKVuJEyL
OE2T2jSyi3UBHz+oB7tjnps1ANmDF9ZCbhbvwRwEWZXCp1+lBBSq7XjmiKZdUIS/MJ5YAD73ImiQ
LEUPXFDxlzTafZ+8Ofcm5dRuRtWbKSXDwY27Ta5vrnR8hQQKvAlQNKAnp/p3RY11U9C8FQI3FxDP
GUqTsOn2u5c81r1dfho943dkE3muTySXQepstGqz+/OzkUdQZrZUK2H04LNwxFnHCNazX5cGi6Mt
Lgju+L4KX7Nwd91Lmv/5FjDJHZJEsCo33aniCUwgIAvAqBmuC4ocH6wFriLGnnEsnQ1Jlh542PAi
ZTLqbqTqBzBr25zAbkVF0c6jfJ9ezjNYkozz9ShSRHuwwsflYRHvkE9JOiZg4wZ/U1tRpfxCk5hu
V4co4YcT1EQA4RDVV5ZXYZSaND1/gjyYVu/3PnF666R+tQVd8XvB2nThiWJ4ZPZHRUyenniS9T7z
IoO1IPoTGk0yg+uK3Q3ns0gF2/hvs/LDJdnsZ/jb4j67NhdbXInfVl53d5wiisSuw+vuPfKmcWYj
5flS5sinq4xkAbU/0ecq5TYsMzg1PzY2n9B9wyFp0npqRFotp6hAS0pUT0aSTdeeotoAbt/m5rs5
7gM6n09AhRc7jV1eEWmaIZZFuJ9b+lvTSK+8GLAmGz7cqoSDQ7zK3Q1xd4cgsREyiNoLS8pzTKpn
29pVxhAe+alAfUVDWDqRyrX62h3gF7CzzVk4HIgjcU1GoGG88hT8jKAiIASXiOl1s5qoZ+OlQqqV
oY8evdipzNNSVDOkTYaKT0Mm/DOQ+XHV/8B9xr22RFoOmgR8PvMW3vwccB+DYUvpcqafcn3BHin9
5qeNWjrue97oebhkw0YbBu6Sh4keTRNdUVvx9dOyycQBeRNi91sp3yVpU0eYpZD3d11IKROiwmQp
eJGdKSBs7Qnckvywwh7hQQyYuwd80rbr/M2/uosIp0VkPI9bUhjOYKoZ1ZLZf6mmsYvpIWhxZ6Ry
HWeaD6q4PFfL1SGsgakskTg+c6ZN8lBl9W4uaxVb94CpsBIUUCsrr+X0luvaMtsY2x04beJrWtU5
ZMuTcpgU799T1AOlVzxkj1UG+Yg5bM2Fg/j/wU9Vzn899j70z2AvoDDoJkQ2hfNKR1C7yJCXZmu7
mjOdl2gNtjXdbfTH+kCxcGBxnJoe/4f41nM106kZlahtQtO2/WxrOhhMFgRc86aqSaAZJcdaEzif
YApAMOFktUW8w5Wt8WwVme5mpLl2dwqz6KUDKOD/8hucsNXWCpKXs0HeP6JuEuHOCAAfsfDWtp3N
kM9TSc8u9XvKv25j973v/7ahBoC7kRnNI8R3nHd7nCCPq5B1uPgjOOz/DQVwJuZ2XG5eaQIQIwEz
F9laCtQhMD4v6hSA/D3rcRYhjDsP1ZQf1xyHK+ngs5bnT/HkROLefOyJhHbILM0thLFcN6K2vdY4
ILOxjbP7eSnJU8yrmoXozDoV/VO2rWs95xKeKRETQowQ7EFiuPpHC1f8nzoa66getRqsAgQykcD1
T89qJ1nvdeuWd+sTb5UQ3H9d5hi8SmiNUvjZ3H/FBQoXWtCqrzmu3WC20QqsqDjXuQgbBYOQAVbB
/bX01MvqGaINIHBxdr5IgfmkpMxylYuhFyTXXmYYrgUYZHoxzdT4c574xUnPmyk0okiLT1sB39MU
Fm8lgVx38ORkSIQjZ+6sAlx8ussinBa9+RV9Lf0O7y2A3xuOuQC4URLdncIto4ABETgMURz6m6lq
ePDQnRf4++7hAORM5pXD+AyxgGSGtzFJVS1cOU0JU75t+0l0C2Fo4brXEbTrBet7sR7U2HfwyOWr
I8YX5hfNEtxGNYEJrYZCbcIf2gcBaao10sz/4owjQMFUFzQLKbXQve+zCCBYyDxWtYJsCE7mHeLj
/kKNK1oyfmUK3GhGS5Qw7M87aBLA0oNo5WoHTjL5sIL2f03lJz9DDEyCX43rHMrAOS+sL95gADwr
dbGJ2Q7C7q7tke4EMytu8RRukcS0l8j6cNiEUKGNI3DyyUOxJpuDSILfaWUNkgALYsRd8BNPHqgn
gZUsLKNtYjYMOZ0K6eKwXU344IRYmezlcXbDkIHMVfLJHqggdvUxVhPLh9rVa0z3p6voULPgv+xs
3zopNsHCrfGas+14XFgFBkVAYMJJCQgaZ76YiaKAMmjAMYhPuLTq7oyzqCWyETSKzFgr7xVc2V0i
jL7U7dSvQK1txgAWBBgmAPuXkKGuUFlVgNeXtlVt2Yfi608CG8ut9ctpQ+Bqq++p4VPwnyiv7NOk
KnBH5vH3z3b9Krvdy4TnNi2L3jSj+fq0pgMb+4JK/sjQuY2iLP+fDWAixDQN5TmgCES5V6+eXgkZ
Tr8IxjQPr3VJVIkUBUDYwe0W9DoYFnL3dBA+MTPnZxqWzPsmp9KApsHqDa8gKZFinCdGnNUPqLRj
BUY9Eo5V6KGGv+MPNCiJ4fRKVCHOnnWGqWBOXRmqlHIHRw7RCQZz76QwCXA/n5sc7Uh0RPcBjoBR
ysKOKjdlVFgJogtxAUiFS9RKMMh4FNQBCePUD/ijXoqevyVR3FLh7lBuS63eV2uwY5qQwcOF6a86
SILYm/gegCUWVfiVFPoJ42DWmCg/DMeKdtUI9o8kfTnKYlEeIHyy8hViNZeMh/YgwkLywaFLj9xU
fZBMRCxettxCA2kamionzEJq1sbKDD/7I5w0JiuwQB+zjI4GaxX3DIKqH9/VnQFYEl/frY/A2M4G
nyyh0bfBKjjqXwrOwYYs10FL1tLi5F37lAxMYLxA8I0roJEB0Dt0fR5GSeQkt7sMqD3U6W8OSK5C
hD+EOOowcyuc5x7s13FCSlTLNLX2Dooi9RXXIoC8cRkclguh/tnE8/Qtrxos+n3XIRTrENhHY6dV
2G9Ic1kmEpJyKTu07UgatRLZW592XIFfBfzQK09k9LyOXfHx+3Fvi3XSkj8vtWzvCO5uk/DDaHgU
5RTn8Yt1wFufsleVxax5YMTlj/lF9C5zaqqdN3NJJxOTNTVcfMp1LXi7XFdtznfB290Rm8xqOMv4
yAwaPYZZAD20tT0SVSwwn49vOqgePL7VlT8X/Ftm9X9NieTWXitCpCtzDKO9bEx+ivTKllnsPnaI
vAm2HFn4Sm3lo8TjHYOidJ6fby0ABQpHvPsWNqNWynJUsYd/onN32OH2gjmAFfWVKTpdl+9IUfaJ
o3lliyJQ42Z26meUHw34P7I/tGClgIMnrZl35vzrZt50RtBpn3ojB5cdMXsy/XVIRzVoceRnNXix
PfW9ylnODDtf7+rFEm3FzJK6B0itI+6ZSnzhIwD0AnLWUegJf35gnXmsrxqs9YcTqVIXHgtekfbg
IhBgBGHbNRPQtEhJLWlwJsVtpr8xk9KFCGcNZarkQ7E4AiXJuPJQ4tGWW6j3kXFD8baFE+XtJRIu
RNp6KJDhL8cMFRs5so6phjb+jCMQvarDFmC2bmk8NxpNwPg3h1yeW9eucVdqkIiSDcOiCS9ftkvr
sPrfptdEo8YaXo82CyekESnoVMn87iyhtlie9WrLaDikkxebWSbnv4a5KrDdeytThJG++LKTYtdb
X6kUa3jarF5uwJedybZ0PfnxCMRlpSvGC7sGTjbtkqfliL4I3uvccF9ztc+HX+OEpMhtKSM33QJO
9dsUWUQn6zWbLZ+ngPGR2rNB5G0LyZAEoO71NDud0t8oGzsE0vmlqka197ZHBXaRUmkzrXJeIWF5
OzMOtgMepXALL+PuAbx2tB1DUEnsuNzMDIje48qkwErTrtmH9kRNTXjuDyWyt/xSXIeze9/iSrHL
9vP5dbHX3l5nSqC5Hs/tT1iAVe4j1cC3sqkz8VCFZERsgeg6U7Sw9kZktEFV2iZ1X+StnpfW8TjF
KK76rwDkPKO9vN7aO20qq8ugI/dDGpfR6zcdIQgWWpV8FioyBAbNSXpbYgv9CudYjK/CVmmraDHi
7u28szoUW+EpRCG9E38vCkYkgS7JsNm4Y2BNrILnxMeCokWst3HfT3l00P1nfgJFiYiidvtwZIjV
BT5D3CEvMLUqV/QctOTzTdyd8s1pOOyngkQODSNm6852Pe0jreJL3PxW9IyVhaWakmw8KFHAnlOo
QbtUaErt94kA9vQQiat274AWlrVF2NiV9hKYsKY/GeeYPLjqp4MtLHk0j+b4ed//F+8L/VzfQDSj
CFAe7WMdu0AV16iMTq53qd6N8+JPj3Z1ouXp3H2lPfYSjp4Hh46BkyXVz79PRgV79A/vNTYAu8Kv
/qyxUza62ZEyH0xThmg0KcaVWX7BRWiLmC9zOXc40yCL7JqBs9rxqwDrqLEfJM76V+wUPoEM9eIE
QdRsmaVkS2IXdoKoSLZwzN8BrL67W/HdG2PUJIqloriL8fWpaXSxZppnQxL4mJA+ZOvu4hTfIUAW
DAIaCKaUcOMYCTyxDumXj2PMu8vpqfirbgk+zrTS8nAkWeRyoCAEPdMCeluywrZ09iMrPBgo+Kbi
b7vVBgH6Q8a6PjG63r5HezDgJRP8K2FBQfwRJalxz6B9of/PBHrUkqhZXitHR3pcVw6g1YoILtvi
7W2Yn965L90Kppzt402qdCUWwQedXFT0Z99nDczMb+Abubews12NciZMUVpqZ/+q6qyuzUVkVeat
hFJGrMBDcXROcXUwvhRPkrcRXt0DZ/WfkYInMLBvJq7TEuwF71JxH96DK+guTcABb7XyOJnA6t6u
tzBcNxfgRy9KDBTuxyUpQBRiDJKiI2k1aLClG+gCwA2ZnSNSFSAarXhifPN1kGtyXjunWFv8QJkf
dUQOhSJSxNy6CXzcYXiGskmTKfrQEb8TIJ+w4LTxHelW7/Txbbz1dAc4yP53QTEvxAQT1/K3hivo
1pLPHbsC0qA2fX0j811v/3Wffowz4G2LxzZ7kej8+DzapMAC4iunwyUXphFE/K0k77Q7KEFIyPxL
Smb3CWS5OsheuC3UT1qs9nOoP78J/1sY3Qtal9S6uu3+jxmk8JMrueWqsOPHg8j3rCgZeCwFmAo0
arvG4WbMrNsEWW5fbTgzOABo2q1Xxm7RG2QjLkqUNKMdUt81pASrvGJ3LeGA7+HqX4bFNkUOACrk
2mizq20AtO9PSHEbTyo4/ShFXChnzzS25Fbj2cuSPe2zWFcdr31xMWErFtVYxNX0uchP6ZYCZ10D
+tU5Z9z/TimX6TbEORYVepumwxcDOUza43JmzJpd1V1tZ6vy7E+d/njGfB92oJaDfJQEmlgBEJyQ
chNwkiEA8eSRgcITVZQypH/AbN+abSI5NDmbNVh6vzEsoSWlgv/FRaAV2HzQQecO1DPg1qOKz8Ue
E2iv+f5DSv+JeuoLrF4r3EzwfVdjZm5BrdICuaaihI5cBVnJPp86zqF2bL8e11OWH/o3a8rkeveB
NyUf5KaZN/jQ/r4t7JlfTy7qZ3rNzSghQT1QuLW9Af7NuVgzK/Ykq7qVJpDo69mdszFILMgTgCzY
3R1o4t0X38mJGG93yQyxLQbBbcS5JLgosh9DmvIJLX8SgO0hIh33/UVnGwCMP8i/DupH67I9a9WN
nd+XEFxv+MQEakF6S0PRB2YFQHCmlUOfTLiklVe7lCj0WxpXrephjLPHkehTm2K6+llsHeF/TWrb
ncfctfQ8AbjYaEXOjUifCTxUFwUmYx9YnhXYthnnQWUjFvQAGnX5jH4cGfJerBFkMcDE04cmYf+X
lRiniOtMypBOZW9cv8k3NZXNeDHZ4aVKPRI2DmZ9PefIJHzsDxmM3xAyK4Pgb0jt45kOWQil/kHi
rqZjO5Ghhs3Dpjq6t6IMrCXGqvzRJU1znj6dE1CbRaa3B5qEVqV5A499pxUoZADS+tqGx0Np4RRP
wRc98mmg4erBrZXg4+2eU5x/bVMPbu0tzggQ91LEdizjB4cAzPoHoC4E1w535FQepDsS7r6jNYbv
LfsQGBjTp6wEvgneTK2lNATDZ6yn3yDUkgqQhUlvndMyYMzQp1jE35rSojJxgyRCwjZhkUColdoU
Yh0Lu2cfLoE/zcP/Nlo4fIR9M0fhGTptL0AjJ20JXJ7hwikTvGMd/Q35sY6xcOurrud+0dL79n1g
0VsVrdfhi3YBDBlnyPiRnFylgoV7dH6Fm+wD8g776N6iwkEGd9L3ES5cv/k9S6vIYI3CSQxSVHH7
T+Ba8eq1z7dP739XLrscwwojH7kgIfnnR1/oE3WPSi1JsVhYUSFHQRvG4nJUgXa9gMj6mJLAxwK9
apuXUwHc7vSo3zDG/ycN2lI3z9lqnusGf/bvNc0P1ggzppPBA2kdRjm4UnRNnP0wfctEip9lO3YB
rXrN/gHZwiDfAhuZ20hgxioE7k4oiFVzy/UcWlk/8EndC2sgwn5vkLUCEOIRxUyp1h5NlYq1DjV0
KERTfcSkBae+X2EBTVCh+cuOdIJqOxsREGbXCGbOyOSzXW6gXOyoajiergr3EtniM+KESL2WGHLo
WZyy99E5tfeltwAodUB6/ly2UbdzYFuuxMyxDFVQKMm5EC8En2DsJJPbg6RB3DayzSYNoCm44v5i
OMAM3QVChGOw0zMkwlH2lismq2yWemU6idKBhBy7c9YEWnOKdPCg4S3eCZpOMSkCzdVJIYL2Sq4C
eDiqVorBHD4gft/m3wCjbxXH6h0znTXdSh8qr6UQr8UZHN5mTXMWxcKYlcVlrRpplzIvCadShF2D
WlIyIPqAg0KY41auSHFpKpYQv4kdDjxqyUFvckN3EY5narI9uw0PajIN3MMVDU3amz3qrh6443aG
iy9F5Cvtb8ER2m+D+q+qZ1ZhZSxj7BoqSeyCJprffz8HpQSdImw6vEbDLGeUxsu/S7Yapjf7WQYR
hhoZrKRy9NZOoSpGVVGN0aVBmbxjGZA+2Emle4nAtNdO3IGVIYAQnKc0s0w9M77fmHN67BZdQblm
6D2kL1b5rs5R8Qr8ZZOUmff38I7Q94lXeDXNkzq3fWrHwDchslMoiCOor7GBxfZenie12/TvkHfJ
VI1cHMpYDKdWY/QE73QTpzjkAsQPb00hbakepMXFtXhinVChXgzyE/wLXegOjklcl1lFlh7umEPA
5vJh7uB9YtHJ7yvnax1deR+gMS7m40QLxwVbGoNkKOwDjb8Y87r/J7e48TdtACstW7bKb5qfg9a9
r7bDpNkINbMqickG6jWXG92iMGg2kACRNHdKZjbr48HZVyqBSvit5zFCo1lo8zAbZSleW0LPcRG+
Hg3Kp0UK32ZgkCXfFMATTMLiBq9fbJAWzw6pTRQkzqgipxKbAlwl05wWghiHNoKuBBt7px1cByB0
pOmcA+ngadp/IhWk5oKDAH3bF8PoKWkhd6y81ui7mfZ/N4E5VJJnmryi+gR02e90UViOBV71NK3I
s1ZKo32gXBHovcGpg6Rt/LPnvLMZmsBCzduE3R5W+Vb7lbwRVUmNWg4R3xcoV5kUgwUkc6p65DLz
f7BcCt35RpNgVcyiPRA4+k0vHxGA1D7mowjjpntkwNmWhnU1d2qamrO0ROhQhZjgBzRJZwogdZqd
SoIEIY4lXPC0Cv9lKL2jsM/pwQIcO8bg1UCMq5N61du1tDeEDCdUDcVnDiACde5nn2sJ/tInM8cf
bH5+RqxrB+KG/NxEYXGiSEc49O1JcYlyGW4py4Su0GRMEHy578PStzBBt2B+65JR6XfMAVuRBggS
hyD3xo4F3TA/vQerb4f6ZEw1+UmTCjuei3vHcKxr+BKY17Z8kWdJ+0/XoRFcmYMY4bghhG3GVlLf
0FKOHsW4o1EUlmRDPx+pMSKj8yXj+HZwquYxed14nYhFAUjcE0f1biEg5E/qM6DVp44Dh5BXlEUB
6xk64uJS4b4Bd5qdj9YdSQZkU6duNlcZsL6IB1hPKumqb2dj4Vp+WmiklmqCcm3od/LK62VqoJWK
K68Jd3rjLMRsGAamSc1x2qi+H7oC6+od+D3e6a2BsdXAkfStx+4qvB7IOvHAROUBFmhXfIBxeDPQ
auJPbVACYx+rECQKrKRPbKYs/oa88cN7hOLo+es36OxmTibD2KM0yt1ErA6ne9ZfrpRIdk/zYwJM
vDaaT6wGbllhQ7UNxu1AqbK0NvOAvNH3LF7xRj/1NxMYm5iMjwLIrCQlcGt/rJZthlok2ya1NhLV
nI+XKt9vATHsicl8c6Z4kjcVe5PbmjIoNzVBEjDw8Wwqw6bdfBDP5fAdQfwzHT+ICOkapdtOWetd
cyVRwf4p9WAoyR80vEdfTfna3xr5WY6R7jd/Y3M+7MW78uwqHpBCGjb5pf2aM/CAUCm1eOphKoZm
EhkpOWlKopm8fYXVQ92l5vilGVkektBAl4htyXGT4hOmPvuTeHvlbedXugi13TDMgOohmJXc/ae6
J1MED9RuLxoR1D7au6nO3UX5VDpevWKHZJ7yLWn26ma6nzvF33PLTQN/1JIN/3e6KatwVkPFtbha
bKWWsqYNjv/EpyG/w1fYqEqqf087bhnL+kIp1pdfwcrZo0QyShPMjp8bqnYjZZjTofcAB1/ktc2Q
5jg5l5FuBj9x9p1FZENr9/5Yy6YAh1ha6QbYbFDNH4hRImj3Mdj+lmDxYXJ2IWDtXWneq8wsn8K9
6WEjUog6vY5XXzQO/WSRckAtIZYJB/1cdZ8FbKIQgOydJJtOmhasLzjXz5mObN/PTx7j/rJ5tvBc
ClzACif0dA6vtfWw7px/bjc4GU5o1kd3dnZvVQdUU1xxdtDQtCDC8yeNi3xwpuTZlXLqwln3QocD
/tHVmxuJ45V5U/8b9haWkotu1RT4+8N9QKaXmKcJcIt5jk/i48iox7bR3YLh8B2Ea+32kihUCosi
qhDClVOBObGEwLehJUdPUzHPJlMKRXBvvFWwqkW8pexcOfkDmWxONS4Kyn5mGf6IQq0dJhMziHyl
g73+yTOs4/llBSBpAMGTuMryp4p5X8Wq5qLYHmPFfk1AuV2dr0Ixyo9OVJxcsWNoqysKIoSrXDfp
9LFmIQ/2gVKBiSfI5Mi9JRxAfAd24/lfNU47AzyWbDGGxF8WnHqnwxentuDA1uzFJvg+wOYtnc+9
dqA4rSUBVF+J+MW0sQr1gcp3S//tKGkl1fb/pkIQEFwqaina5sIS344yS1LgJ6a6YapmxOck84hW
d988H4cKc38rzM5AslolV9xMBNwVFqg/xa6V1usy86GgyTmCrU4OzO3WLPtB0RUbmCQbp4jJpqOJ
SXwtwNV6WEgKzYyjj9ubk//3r4jZJzklfhf/F4At3LAIEFUnJxrJSn3M3mTgHbnjkFg5dxGibjyJ
rbtJD/b2b7hBVf8RtfzN7Rky6/hhGHYq1O/mZLN7dkfKDYdZ4mMw7SV9vRLCXrT6YHFHQnnjreVX
jJPrjbny63jUSuA9kmHi5+mtzb09nTTTmG/6fIT4XuXEfMPHk+Ot3LUXkldgfPyyIe1tLrTYZbmk
B7Xm9oEhpkG4QcWzMjVdqsT2ZsQ0nVQlGe9SyVmGP66ZKgFKgGbbMZ3+h7XZkyj3ajdJ4wZLddAC
ajBPjUeg1OaxiZrfnZOWqBu4aZQDwj+KbewZ9StrK36jLtqsroyXc8BHpyj/1mU6BaNi3uku0qfm
fSYrQUsu5ZSiVO9G4G32SlceSk2EtCEFKqpRf38/0P3bLJ0exNDClBQQvdFWeAaKJ/3rUKz0WVcV
A38/FnCmHayVgtuGXLBBQd58dsALLCZSE3jiGtM0nocCtTtQBrYhiWFvw6K2cF6aoE2NU243Yocu
MwGjzIXZjqe+z0C92D19FOoem776U6hTBc9Q5dH2r6ySpEj9rqzWYrbSmgKsEyyIAf9GwsR/YZ18
1h+TCcFsbrK3JxB+AmACAjwIEYOBdhEiWuAN9C9Z7vh2Ofs2Sctp/tTBc3O3lkni7XY3Oqw6KAUr
II7pV4Y2ACWLH15ece97EIeISsYc8+soxQT54ALostpu2dGa7Zc7IsgePYpQH8UgA7cwjXq2ANex
H+AUQL/VEc+9LVJTFSJStLK5hGikoB5c04rgOWubfyoFLTp7FOu+kekbYLaS95xMYa04GyjfVKgR
9UYh/WN6MVal8nzMYWaWz6TpNn3ImwhZomUNl5g3Cygb8WcCTEz4lR1SmNp9nSAG6sxUqVL4vJQg
gtAynCTJhVklsc9P5daoI91Y+ttB+15d6pZTcz7svcCerVWB7MNYvXQhIqDoEhfOEB4tSsUYyYgg
ohhrToXdaeXzbMr4Ffo1Z/Yyir2InszQCsKd7NXWZ/vGcZn+DRIrLUaJKZMjtWO8IjA88e1iikl2
FXCVRA86YuW83nOgvNssgLC4NpD2elek6Yli1zimuLlw4bUtXk3na+FeJTevCZygfVGQ9nRsoY03
Cu1c0WGwnt7BmHyIjtZycoQXOtu07S2cBQDXH7PLG7Gtp6avxWxQwPlx95rgdDn9XMS0e3+B+VRK
NTWhIJ476+nNsf6zNQl4lG29W8AP2HnWvOK3otMbuFAW4QaJOCZrqwKST0V8+x/dgnTvUEb5qkrk
SkUzTRMNm9RL/43U2lT1UonGVvs88Ic02mZpTDKRoK9jAwtxwTjGNz3qCxBTfvqC+uqWaIGd0Ymd
yG9a0fCqIRwVtLel9XifLx+6tvMeL4ZwJvJYPXS1XQ2p1+mRD2p5YxFHs/qy9PbHvGjckqkpz9aI
+YGWAThUFWe1tktA+b3/0DQX79FAYkSRN43Z/yVq4ypuMQOra2XD/cuBr4iittqQwcvjy9ftCk2x
r7XPq61oar0+J5DyQ+jc6lcegXg39mXhvg+0IkisqpDU3EhWNhurVgpXYRjIEQ5O8IIG/Plshe/H
oXx7r9Pg09R0H4wofyPk0IqKGkvDpl7TlVrh23t9PMvR07GLt0VNalFrqBa77ppH62RpzcqHwUVx
V6lWed1K6ghpBogMnPsggZNjtFg024D24c189uCkhtREOe03x/QjAXYLxLWzEQ4smtmCzcgoamX3
3RE2/vZ56L3CbLJEWCbYRaUoQ+3+HnQ8MLIMBkhCCOzClGjpXnTvrxv7Gekl7omj4sds8b6INxas
4IvCZS10emGcUWVO8JRdAD0Ir9+GAse0U6qAzhVbVgkpNL9AU3hGm7vcdAJrYEeWAv+rDlmihBgP
to+XZxR+ym5Oo6rAqmR4Yx6wlUBFm/wO1pBFLbnEko10CV/2nng4IyAgPK/fbpCzDoXGfL8fAX3r
qqINdypOQPumnLZGNXJuKjRG/LUPfXj+/0mb8AaBO+yovVALl32kboKPVXbEOQMD91T+pFi5Jh7w
NmmOUt9uS+GrYP3A6sKVx/5xi/lFsaN0gv/r9wR4KQXS8k4yHjXNsk050DMHIWAFcT8UBC3MlRyK
os2AfhvVHr6cy3YIdroSGd5nK2ANrc6KOFbIxY8X4PmIUPQ5NF/Q7i8M/va+8fA7QoXa6p+dsSAR
Bzhb7MOdP0/MA8LJ/hCfE5okpWHsAzy8XHrEH0jYjHtj/I4Q++JHSjTWEQKC3BG/lDJUtO8jwjZl
UX9ZWm7Aq0BTLsJMU4wNzRJbL/adl7bPmasC0haNwBUs54a67DbrR1Es2jFnyr4/LYjcoZd2QWhN
5rtc3HkbLeyaJUzMqdRB4UhJ3Fg1752rviaYngswNFuU/PP7MnrTju052NsTOBu5JaXCkLoPils3
IsgH+rh8ghDcSuzpa60BYKwX3XPz5rZCcJbHzFrA1cq9zxh74yk5eYM+N4/TA/E7BeQM0/EjzpzG
XESfC+wKh4LjaNJ6Y9TbauyfA5GLIdTKnxWOuUbVScKYRazNtPpDAlF75Dy2BOzqAfcZb8eSEMBS
U16FCGc7dmgL/ptZQbKtcTgOhpEVloBc1DlWLgfr1ICqRc4vK5k3mAS59X645Xe3evEqJLsabR4Y
BJK44dm1vEmcxxzpJWYd0XIVuCBwVkCKOa/39MuP75BANaRt5LcQ5Qr4GjIrNjg7HEn7b4T3xuH8
qRsXsjFD/ylNn2vEHqPhZkAT+Kq0fXg4TcWe9ipcXGrdDnUtHXMD4k7vQTMkAOuBBp0CK2G/jkvU
5nM7Az7QJJqOHZaF3XWoHLQX0vxlLPBbYnvF3wrjpIe8FG4miF3iLQbVpKA47wlu79UW0iP4ElRG
ZDm7UAERtLwctegeERQidx5T961lIyQuiIzQzAZWexAe5NJmw95QJ1bFHbu9H2D0GtAOEQlG44tP
VBFjvW3+sgNeFCGcvT2TrWsmKGCMy6rVCSEOxr/p0RQHWbKVZHMr+9g9eB2E4T+WgPhaBFyVqFkM
WbtHBY9xB/yOn1a2tSJJjEzMCM6LVTbAwN+YtHb4NkCM53ZsDTZ3B2If149E+rsmKhDVnq7XNiEF
aZvHrwFcNQj9KxotCtiHlYUrOO3+X/xk9WfIBCz76JP8QkANO2p/rN5iIT+1XMmc8c1koaTN5jgO
4iJ9rY3EIjVvuVqs1t/IGp9UP4jqxZn/j/jdRSY1HOHOZzqhCglbaCzGalKW4Bb1MHucKP0z5uRx
gbC07yRY7cn7H6qCpvHpTK8zIe/ace2mbj7txWV6HlM6Y3/YmxkIsUYhmkI0i2EpE1JqGhKEjQAS
VAj/RtTgg2nETA+bPAi35aBFC/RHsW09ZL3vslCBXmRxv6wtqufHeUuOorFh9faQJAkrzMP1doTy
2TYaVU3eXRd4MdEmU6ZM+uXu2Us2SCPGjCCNUr93XcY/bfqcgyglPSDEf8S/ZWRgA4PqkCjT2jwz
L+HzKSUxXQE18rC9MhSZd3+4FxRxm8VcSIOI1nEi7fBVs2hl781j4s8K4Y22S8i378MDOlPNNdkK
Sh82KEfHyWEzGAPP2U9wYo6yQXEEj0Kqbb9VbIeCCEUVU1+q8jOw+suAsqp+9R1VYIwkKUkS7o3K
l7FwMb8ds1cQxk/A3s1EXfUzqzylEO1kDQBSFuJk+h1VG4+qCD4dr/nwFl8a/NdCmG10FpsBURfW
cHmhL+/ixOqiDuWBJZZOZBa5+lDuoD1rVCtz0g9VfQDBSs/swQaD9FMuVFrYLs7u3c1KGZTuHcxM
xYm8mB/vwSRdtD42Ddm4YmIDPNHNpHsm3oD8a1x9UXMCpq6baNxee6Q9eEeGjcPDdJ9iFsmaM3Y8
F6pqvL49ZREoTldifTpi1rHdLfndwyYJYiNMJ0csBQF7QA0M2gsmQU6j409fRKVLSNsM8pckyscx
R8A5Xs5KsTl6X8twvFOZUurG3OPb52Tug2xnZRyQrBROS/29kaVA/1MNvCWsP80W0tMF6lHhok3Y
yQHBFjS1ru0aTxXaqu9+EcPURCZSboXn5Ppty3jKAYQiCGHp36W6lor4FQGQND0pJ+q15GGWDbEM
bIqF6TVUtPSKBjYPN/6gKGMmpLd4NKnPB90nYPdSoH4wr3IgDbwM0aUuiwsmSqTyLS6ID3QQ/FbV
6Yn3obzqwHGZxfsjKHublfHCbnsaglLT069WKSGwp5YlRhY9n26vzY8dTv5tdSVp10MrZnWr65GE
oewbFJCTP9y3hMDUh1Cub3QNTWJth4ZAGnuymYg3imOh4DgUfDmIW68jM01XedlwigQDwQ7/nQLj
pTgsIUMwnqysSGEJfBgQ46kThVN+lP6XnFqpLou95Gv2XCTTXUreQQb4nkaF8OuEx6KQoHMoJUVL
twVh6LYD3aJpWnzzdIHVoSZDS4u7HUzT6AjCWEorxE30qEJDCYMQpsgE1WxT8tKMxQ1n70Hcm2qS
5xZPmTig+XhfwYXxZLZEdiY2X3U3MqZzadShvO0ltpA7dr8REurp1kqPndMJIAO4rPQHZwlL1XaT
1DUQKWhs/100NAdVE2rXsAYox9xHsWoYfodLSf3ayBp+/AXzGD1lmrYSIbL6ybCjqFQxZaCQjHSJ
eFuD2G3dKADXahDOJBOxVxT/i2YpXvOuJsNE9529K1MXE7VT+arCjmEFVm2PXE6zS9ldoEdF1cir
6FoVQfcrUuGaMSONLriLpMpil5jkbTxL4LFHHGIqReyb3qWFVkD9Gt+Y8PFpuARpyi9BJiNz/3QJ
szHDdMXduXkI/BR1eUSXXOyKX1SGNFnLzsejA2xIFq2PZPne1FTLzW4c8MaLyZ/LiGtfnlFxJIIE
tMhB0l0a/gT57NBXtHVvOWhUuIDl9m3tFyQl5kWioOdk/j5AePGRw6bItVBaHLKlHP02TxfwqboI
x0TzPl/w9VLy/5OLSd0Zjlf+3+3eZ0kj57+qWM8YuIxkk8CF4CBp00uWMx9+bop873Jx2TtUoEl2
ahZkA8/+Az89sLzvIME7J8RdJCcbGyJ409d7ehh2hRI8fRhSSiSHraDCLeXI5+4psCKzfb9Wq0AA
keU3a5G44tRhGmuBNWfQLlW3QOemJn+q8x3GE6nxZkJQ9q8LMgFwrx16EXRHFnTldK82bcB/lgIN
lhk4q6/zr/PoAiShGrGUUS7WpL4PlFGYLbApHQVxyUQK2/U7UEFWt7LXWZJ8qNSNpx2XpLp2kE1o
fwIRs5xGA+XoisaPU17ZEMk+8qq7c+SFwhGRDX23SQZGIc2Si5QZeyDLroOZ/cW00WWinT6ZSxsW
gGS2OXqnknCiXG/gxZmfn34ncY7WZ+CH02xD6t8UUfnnOd5wGOrVqZIM+j6NMnRGkyOb37ie8x4t
0llT8spZRNyWSnVGc+DAPvZGjgxwH7+NoHO73L5xiK7HCFX/lCpisqBlVp1nCPmS1xPeti0QLO/U
T7HRtoy1HePr/6z7x6O+gSmXFkbs/pGf9ZKZooQ3+rt4af3vLo9Nb30oeFtIJC+3TV24iddmyCI6
EHwMaof4OPE/hUkeRS89i2sazduHekj0Fzt+eBIieUJWNfGdbcyoswqiR7QTP92FwbrlaYt/rPGg
yXtyMvZ9ybRMPZxdwkEd46oMWmP0+fACjxd8ErWEB1XRyset5AuTYpvzbcIjX6hCyWU7zfh11Scu
tP4IkL9maDWbGcy39oO/Xa7PNde8mi9oVaKQUINJLHbxo0DZkAJAEu4cvgFqncVmwkF3ktC7k3d/
ReczflbK6Ubi5KzUp3NQ4UYGdgXd+B9D356nUHiR5iNnm4Ys3baCEGCeiz767CsKekPguzXQpAZV
K3HnhBrWz/I8LIDCYvUXVLIWDBePe1bQrFS4N6RYWoOn1+1eN/9wkZZfIZycp5+bH3UGLyNjgEOI
CVTE5jmdT4e7CVTL2CJiCjz3dYrXI8vo8DEigsJrpsSydVqEm0DussuWqt2Xw/wx0fZoIo5xUfO2
ls36Xn0pqz8B0bZD5BR1rt215jm3bnewLdoPcpMyKUw16QkbUOBF/Cgi0fF4nLaNQv+3D9PqQNI6
NlurAytfDYOMqar552Vl80/+zaXLe0F2cn8uBKX7EQMk0hr2rGceokIdvqwGcCHgE1hGNpjO6NEq
4DViQGSLGMa9DzxOprG8PJkw69WkZWGce0HnDl99VWnk/LDJNwGsLQlVedmxdkCTV47JpkMZmqfR
xq99YpIuWTfR0ssTv6FJjPkojcP4Zp+GUqGRvJPUVPeMlWUw/QWrEjmS9wLhDb69f5tRz4BzU6YO
JG+3VREwmbMLmFRZ3DDacrgAX7TOWqmQEnq4rgQc51xUbPInG4c+8QmuRHvokHAdgKHEVhfuuk/1
isCEOWhq1T65HoxcIgjv9SSZ+xYUHIwl8BJ+COjd3k4ELozm9EI7d0fAoBTriog+npipCEDqU3DE
gK0D7DgzLuJa81DNeMaykzwqTayNhIKpu8P5RpYKAqdNxsKMM7IRx/Nxor645AiKxPJctvDEgXmo
Wia3VPkY8XHLjZTDu2HQhv/ihPg37uDfVPXRErp2QZlt7LUo7tEekfGR8wnUz7Yfy3DHDxKvk6ZI
sFxMADE8YZNUwyB4XxjevOTEGpRhW1SCwHZvfMC6s/Y9spaOJ+cUIq6/L4a896veVQxdzT1PmK3R
p/yRbH7qRnorg/UXacDi90/+Qr2sLlWLJk6SRFFZ8n0eZHzAa6SF/unb2LkpeJLoSdhkcCxR7/Ey
DqDte9u93crGA2tf1UxBm8j1JUAyxq6UcZ+1zeZPRTg3epJ0CsgQGYjLQix7SXcgsGPRhrVWpIft
PZPt8saAgiPfiWbbDqM2fztxAN7tb2cixh58Kfxg7HYhdAW9YYs2+UVxI23tWnOP3xddbgW9cTvR
i2tydD3ja1rZ/AScxavi/O6AWqdMP1EYvNBBVQHzO4HsowRKFOG0Bov7XkiwN0dAnsfykhboXe7X
JcO+a0w135ILENRa3kaM8JH+Ounz7B+/Yc7Xpz5Pjgjf14uTxxnBUT3vqZ8Ky8xOx9WHFpoWWTiX
/X9ysGV1I/D4Y5Mw8cVYN00Qsf207ivXMFxpH6GsafIxw+9ZlJRX5IBMSRUQ3G5IU74Z8t0n5I+9
+gUPhLUoc2oTz8dDfg6e0iZDLtZ7tgAWHyorFK78gWAKoU48IDUml1f3kY8yFgkvwni/UREDjSAY
v+85EiQhZ0Jpv+UABf5nHnRYOVMVz0mURZP3HyUPlPfSc/xDdSQhvIjyJAx2q7iAkgIHhjYaB80v
57TQboHQ6Q6Xd4npsEc759x+j/UD+EZTyBS6eKjL8yPCBfv9/z/Zmm/zl/B1LW7UMrIvpZC+vKJM
VY481NH9AZE2oNtOHY2e1nWZeSQl8mhaHY69l8N02syNu5wwpv7fRoRc/4Entx68gP3YVOmIem43
0tUVKoi0karZi8IP7Bb5cBlsD7yrRHBVtG0Zak7ek19K2LyXT09D0SIxv06BcysnuvWKuMhJLoha
QkSE9ixG7GZa7GqgzyoBbB6GgasYAYr4GzbQdPdPPgFBCDt1nggRtyYLAOtzb8BnvIB3wmPez/Mf
Grf3Ip3zRxeRM1U8012AdShsFRYEe59OUXBq8H3RyRZ9K+XUJJAd9npGlzu+ZxOsE8jUrJRDSqaf
kFiYOMKQ4A4EONzRcLtR2whwevMJkn71g90ewB7hItl6jrbOFhU3smEqfTmCcn53ryuuYb4yZ9dd
gRKRU1Kf+oUHHdwPyh6pWzsb5lwIg16iTEaATypcmUD6dXrwp7O+p9VXFrrNhJIxG5aqhU61TEL2
z/Rbhg9bAzz/y8tnOVt2l7jcZN06L6Kh+Ko9WTClhAHdLQ6eud6ldIJk0KJhBBHIFuKlM5d/ePkv
+n7tHzQOIFs3n4E4mHppWPPLndIrIUMZBAgE47l0WCXPpRR7LFhbxmqqul233323XNwLG4armYgb
Uvyyl+AOwiBbtowJR0GwTQ/Lcj3iE4CndUxRrJwtY5B5ElQoPQwBM7NqzVk+5Cmv2itG0id+xQCA
LcfEZtSoi9UIgbUGQQfK4jkiA1T5X2f6r8UYS/6OKf8kzESvcNHPR+XRXCGRIUGGYonGRMjfJJvS
mRuWYT+QrasFxxYyNQ+lMjaJpoGDuIBVGq41hxo1qAWJ5BpGqGW3m67A3L9o0PTSZxy5TH+Q0hvw
BXB1WUk/oqvNx4q4YIRo5k2wFW9T+GcAd7ZkGMuxAQ5AFZyJ3+GAYxsuzkf7RI/mwWzDYLzLU9On
GLFg0nN4S9ftFLTUedKOWYAAMr3+KQGk9iX/Vses55LUmFvTAR4FSSfBPAysnppzZ4+5/2Iobi/4
weec5xfeyyXsaHEy6PDzNVsmvcmpknQAqH10LqYtwnOX0oY7XFxe1CPerbg+gDPcplSWoCg3ID6x
BwtC0wXq/APXgAqfFkIM6OL3ZOGFFLCfrAffPmeFftCAAFbwSiXTTiyjNgCc4KRtVdIlCH+/TMpr
f1TLKYvFhGahuOl1XgNXC2Vxkng/jkbPlK8xFzVTr1zIsLDJkvwcI4HAs5xMvAqOO0nQbxgYI652
i43FJxPoQUBZGoUCmPmFCeonWkBXWPaePNLz4mSy9HPVOJvjuyot4dhu/GWQdqU6ayaNcCKvgL8o
CCBwd1nHDR3tR4aUKsZBo7A5oJrAps8Q9ca1f6fhUnFm+OslurXSgo9oPwsAztaP58p5XZVn4B9g
v1qTdPCMqWhcyxwgEqb9woR6LMTKBy4PbhzUPSsGPc6D7FlhZvUmUeJbcfzDWbXyGJeaKKaCGN2N
V3Tas5z+c4pTxVVZpmGLMZLuEkOk0gmxDQiLLqNybJu+c3gTE5303KqOKQWwxOxpfEDnWLZb/YDF
cp0e7P4WU6wKpOcxGv/vLjHIDczHbEKZ8fELzdboxEeXhvf2wOgHSumifAzR16rKdHL9OHdzEccw
GiVQeTtQdaD07+RZlPnn+CXxx5SNZ3HIuFOk+9yUD3N0Ar1RwXeojb1Ge6hMMgkH1W0PICfkPNYm
HydF4Qg0SUue/7kVgttCLKHer+A/FxWi24bj+piB4Sk9UPizdLfgNfYtzexTXvFr+2vAaANcYg0J
MkEAhHivxzr8/zI/NQDo1Kq1vb+zwujsx9dMJA+4k7obme/6nYfH33pAWolpItyK8fKhrFOG/jFR
VKKdSLG+AATN9K7dqKZ2L7p9kUygOIeLVlt4hcqI4/DB1ftoJ8y4xOsW32dFWE3dO7rXZSRiToB1
3dL55KbnlF9txlee0qi66SZYEuNrOAfx/87/kB4X/uVZAmfx3ghEiz3dYdUBqer9nLlntD4EwLHJ
ciApeLvZuU5oVTkKCHCanqnfDxYwdHQOU1Vq3rw0QqKI5LJiikTfLI81euR7FkzucaNAKhvvQoJJ
GZnJsDgqLIkJ/gEJO5QkX28mXs8ipRO6fkfL9E8MH+MhRbrFVNShiNsnyUw9Mf3IjvOak/Cg49dJ
P7JwJU9nwhWaG3ia/zXw7Gkg1FNDqll9RwsxbULAU8xN9YX5QqUPoqNc3UYVrPT/EinktFUcuzaF
R7gePlbFcVglCnSxppZ6mgOM262ExHoug/2RiMxEy5Fdll5XtZgIyJDIWQpGIWZlyD0pyJNSDftK
U7XEHf3VkNm4qR7HawqmXI3ohBf7Zs4U1yuty06PKFtlBrmUwG+jCXOC0z+EdPGrzXzKubsouH+T
BV19DwDnSUybTRgrXlH1TGfBCP2e/wLJLmuuQfDijdGsdCEks+Qgxq9iDLgmKgCz7YzLvLbfwGEw
x+9subTuoAjBDynrm88JuzU9dSBQBdDyH6nCjw88WsanjrU8st0DZIOoqOy27Q7ibtPfpYdikTXf
VTgBNExDMPCevr/xLy7W2QASv/vYGIJOBE5yOd9aWbUqt2b46fJUV2vqiu+gPQpj+dxX0tTswoqw
uUwQ3sVTEXLdEK6e5Qnou8XPtIZ/fSnfBjf3il7D5VUl2IndyX2iWDYCF41QU96/1gcVTzHYSJCr
igb0sUp73RsYpdEGhCsua1Q/gXOg2M7VTxbmQQ4qAyQwPNm/RZo3uOBVrx3FeGLy2DaAnEFuU3++
KB1a8nMfsc9C81JsNlNc+vTexVKqHF5GG3i4ycpZR6P21GHpfQBBO1o4dODpGZ4YEfbw+974w/Yx
+EhYx0TiQAndWniQLtdTfdjTIGtRNyHXtdm/FUluduJbRhPJRr98l0R82JBxykA9dPZQnTBQL26y
NiVRIKIh7mSYp+t/vZQSbMgJA5WljoveO4ZZauMJjcixycYRFfVQXpzN65JBixszlanOKdnrD64f
wx5UUQhw64k3aVVU5kPCutcXCjby9CxvATSwucKU4dRWXpZ54nyhr5kEHgY9knq4Nllj3c+G5t7p
alQ45xsj3bfRZbq9rCZmJXdFtu/YmUamYhec2ELTOcHIEbddQztKW4Y8i/+igVw3FMTx4TrOkgz6
u1BMq/4fr8fI9uywwUaNy94ubKKAQn3Jy+byQEdJo7RVAFnMDf9QPawu/Uavi0B/haaYgrObtujA
G05+Plmzn21px4RKBsYDyG7qOyTPe9calwj7A9aSg4MhiRWG9R8CuvjFA9DT0jqbSEojiU70aBO1
YGovHk9RH/w2QA4opScm7FVgPnG199SYl0wVHQtnjjpVFa2YNbcPwOTEucVItAHRVI7ryhsW6vOH
ekW0YGkyFkPCUSlbRF5mOpUZEKcwc08ykVXd4EXLhpPCykfiEX1s6Tq7M9RvVktP2dWGHS4jOCU3
huDlwy10dSNEvBT1D5iz0Jt+UBdWZIn/Xt0j+5mGCe4nDSaV5dc8txMHrS1NzI0fQi5A6CO+unye
qBD3KWwEkAGlk2uExZtWbdp/c5h/eCzSuBwWYGRUcoBUJ9GFPLD9zeeyMUHr2zaa1vApj4c89gBR
OB/B3JE3GccxeBXhcjERqV39aFHKgYGWUXKHThKGzJENt6GPxwExQGS0/H/Rc/mcRkQP/IuNmT8F
x8/06G0RQchHM4u7BuS0QwBdLD9RhwHiDcnF1X47t4tnFI3FVSEoajVZZ8/VXUUsjLwKXDLvB9vK
p5m0gVmGM2se/whD53lppfpTmFNBdh0qWzh+jdadyK8jyJjCyfolF8YH8k/CofjyqwNB6PTok5pR
5UUCvFXHRG+j9b5/SJZ12LalVSJmXr1W8alGRsL7VnjqeBpW7WDb1lsDunyyOAne6fxI7ZqTrsaw
BpkBMmDeMUOEa2fxM4fbNwSItuc7S9QB+dqIUvwFOZNOGBu8tCG0p/jLTiLBvtaJmt5t2bh1c6Hn
FPmctHTxbMC5YysyRQwtIfJA2MYF8zA8dvknNIEXdw+w0eVgPJVyUERiBQ6susMe+dlUeDVvEhZh
FL4GfXU0lN6VbxpZUv7nvyxQYp36mmdSQZXUqH0yAazOv9Mir4QwfWh+JDEzV77aZZJt/GOr1Bt4
DXdpIMZR8zDAVGHtyTfDswb4qdfjdS9Miocc25mfwBBS0MqqyQCLqMkYfm3x9GorWcP+j1UPEHMA
gqIUiZER4jQcwQmmB7s27dvNl2Wb79FrggFqsCYMHtl4fusGn/fELBhpaf29Dhrw44slMZZqTkNV
D4RyJ3Iuk1zPDhVKY7YIQlmxm5yEwLcIbBnOVYfEECWOz0d/eFss84B/jrpnaWvcJ2M1MS0wqJL5
YN9Joc8gIupvJQxQZ++0bMueWBtbztTCPj8S1+2uoh3llnyJeyUOJR7Ozbb5wsB22dJPWGnpqmce
rFUXBpRy00/ElJqSrR8g02g+ECLtlZhczvqhZcRvuczGJkN+DR9+TcTLeT7ghSTKxOHJh+MDKk8C
7ohooIm7NIX+JSK4u94kNzG+yr8nta2d6qd1mKFgIq3Jun4sn18IwOtVyUKRdty+4GatkxFpPKMu
gdJW+rxe/UY/Q1s7HaKaxIUHHhBi8vuE9NS9fZvrc9da63pXyv1IpKWVS1PCP58kcMg191j6i3C9
YDY29mGrHnQ2/zGUALxe7NI6/YwpdvzwUxcNvBSSwQPxVJPgB50yNq8EiT4GV3sv1XJPZH4AA7Jj
WkYFR+eqZMNbMwC7tXEZ8cQnDc4hMebl69JalJDizQQpBmq5rskBNiZyy5lF5HOWGZY27xWhf4Is
5FZHNwucseOukUhu/p6iSmdnNc+xEn2BwW1vjr4r0Iitc9JXORXJdUvvc0J7/3tFeWT+olhld8fX
FSqo/ObMpumCv7tfRQ3f56HNTm9ntXNliMLB5tcPCoBgQ6nnrvkixh2CB1PsOic13dYqN9z00A+P
UQxesnYdsCMEsMBqlPV30AY3MlKh9ck1F6py03f4MxelDer2ac9I5rp9wdCFSodYQM7Oh6i4wYjf
uWGdeyH7WZtn1Iava7YfKOZbx1EG1sSjjQVnJN+wUqHpXbdhJxOvl/72nbg+k23q7CslLgB0TOri
wq3SkS/yhSPmQUS/hEX12qYTUl/C2mni57FkNQV0h9co1vcveqBmWPl0zVm9/s7Ev1TIO9XAm1/m
iWnn/x9Ee4JnJpFuoAPlLHG2uslNLzY2NPbsNahD/85ZUbSLH8VCWj9Glq8BNISGNIFNj7ZMZML/
jp2xguTkcdMtKQtJP6lOJ2IX+aVwQA6SQOg57wD74MnMSzqkuXiWDmFqruJR9NxYJG1r3rtiKgdc
Qz7JPCpmwZ0j4J7kysM8LOwXH9iq7p1KVgDZS7DYEs87EmjrD9YqtBdJ9Mx+MNvkPOBIm9houFul
nk6wDR1JT0LMWAWTTW+3HnrYqFuUlZlUuT612IbHPXj6JyGz0fPj3oWRzKcwEkxVry0bomQXotxQ
fBPx2bT2pFINh50pcnpPthzi8LZtVLgB2kIGdCa4lcGU9PYhYhWHQ6qctxfIE8Kr4ve2Q7ukecgJ
sNUXJWnackjw0FzRcC5jrv0YfGXoY+QRKUOKgiOsPWS954iMFSUEjvK7pDun2iB4rruzZfl7HkZl
riRi5ACqB3eHDj4uchPNeGdeAOxl/obCfkD5EHffu0YbwLHNgKphjcblHHpe6dDy+wYUJpJZDMth
JxVi4kFxVMheS/lVk2/7jHy/jsSmi/RF8NsTQueU3E9tYl34l3WmdysLqaNzCQBjlWDuS0yd1ncP
0nND4bDf96WPGfJdWa6yI4Ryaxl3TXMdGkXH1ER9WmTSvfvGD7sTVd+/P7e4v56ZGM/OYsUJRYWF
jIi/GSE5ieFWKQwvWchzp+Sh7VhkKETxIN4aBJ/PlnSpdiz57Ughx1QdB7p7iPCi3R734P2Q9d8+
6jUVjiz0oxOULBhw1d3U2Rybx86ujpWNAmAt2qtFVwibZsRDSB7L+wy/aXWzineDwJh44Pof9gdg
9jcJPVOEOL54THe9A94BUdjXqIHRjbudPQkRrf7I+haChzI18pCOVU4XUsPF3PRkq2H+ksaCeld1
TAcC14n0knjdcfyT83Fy40yCtAXD6SFurRg/Upb8rUwEZe/hljc8n86/b0pskNpgdYKj52XQex1l
AeH2XKRrgt1XAnPmKkOlyhdLd9melCghvJ4xEL1hecX2gjOcME7z4CbXgTnHnMLnTBKvZs2lrIbQ
johxeR6ugOfPER29fePFKakn7twTA08ANT7+xqkrUwqyTFeZfQUc85POm5AQBsoF9UkwMSfEv5Th
IKOztRAKIwdsIxKjNwlqAmfVpGIil50PJXIVSC+vneqC9Q22nC46tEjlpHLWPM/zfqz0wfHqKL8O
qyrhSrXcMNUMW/Kgz4yKsF/wfYb9I4+bSgNJbwJGIIBmjlQS+3FzY0PtLW0HTsCwVE7wjrV1cczp
EeEH5931w5NNn7gUlRB76hUbcITWa6s56TwxYRwSmU4AnILf14jsEubzc0AKu6zZdDtCd1t1/W72
bXxEbX27lJzSjBLvUhUCEHCOyjl2S/5rj0P2RLzNUiVLGJ4e7Zmt5+N/5/L8Q1JivJ9t8aD6/5vw
ETfOuaRRszz1mb2FslrUHzvyql3Ab580X3NL/1jdC799bglvnndY44XZ5QMulT4ZVzJfeXIBuQpE
S24UmM4gJGwJfiW1+FYk4uo/QWafY5l4jeruBUxdGGOp3WrUOhoZan4Zvy/bVeSOf/2qO9bqLXzw
i3Q08eZGVuh2q5HGtnop9jGteyAjFuSBAHE5sxYCg2rRb/YSBAWR4LkojWPnY7eCpqtAWJLLLZ8O
JzFivPKqTE92ulcCxpOtwlA+Y79gocunu+VfZxBujOyPKMIdHbD6hj046+1dxglJZ6BcnCmTa6eB
tN/riI/slYu00PYdJZHdNxlsLf9cGfnebfUsitK7HO7mWVDI+INFv6aK2Xj7DVdt+bWZ0CcM62kS
5KvGNKsA0/0KUZXClCcRDSdxwFT2f6W9Ndps3UUNq6gjfLuojIcH/e15dsf3FA/WPYvOhXfuE35w
33ZNl9Rm6anfRArnCWyDQiMelwwJ/vpDn5bXJUToWCYOJjkdm3V9jNqtTp3f5fKyDt8KuywwJnAE
Jr+oNYYOS89jwrAv94yglkFzZWOK6+t4PiVBL7r84UwIuR6MvFdEiEu8a40w85CHh2i2xrwzMfv5
52sajXxqeGO7Y68kzYiexAVFe6CE52xEZnoczJhBoaeO6zWa6DP0sOmS/0WEdmn1hqsWFWkc4QPa
vIQDXOmhTUzfwrxtbB7k3jlcRmnpSGkRn6jDhYspyOzGOn95iEviSgoNIikR/lE5/JNVUGcVF4i2
YSX2FKxGFQkQkdptDJGlCMrLJzqPPNNPXYbXq9aZHDaHfMb/9Y4+4YsCoKcDEG7154f21cyg3ZMm
HiD1dKz8Q5orLYyl+anz/T5wgzidnWER18Hy+L6k7fBjayNHwxqP4CQgUntVtOrJ3XR8GChwtZ9c
8uqQ83nO/SMgkSzdM3q1yOwkdsb3LHj80WzhcQWWaCyQJLPR4P/LqgM5RsprWJ12a9G/YgEPL1RW
DVPX8jSL/5MJFZB9JNGjVtZ/psSeM+6T9OGdEYiqc4rGxuhNat/SvkCDfV1NZLtfJDdc0fcuZ2x5
ybpaERNswx6bisdJS3uRvrfgMY6+ImviG8OcvbZFjFzRGmUjOboMNhwro/3pgbv/q0zfl0XTtYBb
TSFWfrm31hxjGsc3YvcnIbgq15SHIv4NdzpOzlUa0mfOYtoASAtcHIh63DHwr/cYuQUIcG54DMe2
5ObTAUS3L8lCUS3mruYNt1RIZJygs3kS65NdhObGT8cOoTEHpG45Yj7iiE5+nO3N3J8zlEeM24e3
TMqJKT0nmwGgETmUQ9Na94mvY+bLfJgbM/G7h0QR6Tt8ssVu1H6WXNR/YJQNtLgL5+N+pPGE1hOJ
Zll/lVlmqHlqNWkFGRvzGoNIUIIFFQma/DaRtJgDGlJ/5FblnCJTZFue1jE1lXiX/yGBk4B/2uCg
UekZWWDMASHkft7QCwx3jPObnzGmXClf0UxdR2+s5Iu/u/MprMbmlJ6zO47qCrimR6wPiCQcr1Qc
GxJpIRpzTBuNXXp1yveFzwHhmxmj4FpUrBNC9BU6O8bfeUP9RdbSeCJ4spxhg3VZ5DCd6BZyr3XC
koy6b3Ok8GycI7HTg5C+ggeyNsKmTS65lINEvvImyOkkGVk+XWKGxm8HKr6LlxXMskd1zMkzlNVe
+aArjtkOJ60oRgpZnKlkwLKwcMqlB41GGXlFikYWIp9n66tPwRGEabTeKrIjSUh9J+kT/VFF5kpk
gGKYEXzC6I5CXb1YyhEo8LLD0v6AbeWrk/+63LpuJKhRYPXF4iQg5Wg+RwMz1eXvGS2fxfq/z70G
vDapJha3V9CsRIYakH+VCqjAwJPe53mZ3OpZ9uwZ2fYakYVixrDjS56GILOr3hOLoXuSTroG+0QO
FcDZ+twP4IV2EvTyTzIgsf3CPS2se6d+s7gi3N6TXgWK61//67juE+GHME+4sLs+gcnl8YsfWbRx
Kicqw/C4XUAIHJCeWrzPMxasCJbT9Lxtrbs40nBONZwBmDYcwxsgO91tgAOROs/YmZstOtQnVJhv
dm6uGDTYwcJAk3QP/J+EZmelzVZp5eJI9ixJwB8ocsCQRPQxtvXe7G3WspFhgNumDnX7C92cex5V
/dtDCswpWE7gdQnzCqiVpdPrGeL6PXqgxR7IhfeKll03p8WflVFDfK7Wk3V8uL2LmdooscM5324B
DEmrjoNNsl19tueWpK1SQuCBTlcC/R5q5sgLtwiHZeHgoxnnTUQziNYxVKX6Gz1hc/s52xezkXPA
GwGj/G6t4Z5chpRMlVhXWWngP0dicWc/OBYqoANf6k3VfQjB+2PtMdSQs/XpoxvLbG6Qi1DcMYBY
6IAguVIlp/Pfucqw3uUnTphCqMtm22/bFmvcVb0w6yqagPcvdn/2OTbei33gKbLN0t2TlXn/NZ3Y
YlXl0e3fDrzHUZf9ytC0hxN+FYSzMs3z9bSQYDbEYsFreWCcpuJUHy+ApaxbjGpCe72ueSs/gLh2
iEVKgO6LK0AQqsZAQfVScAmiQfIyHMB4X5jJGXBevo2eI1IbKmoD4E+E3ymoLc+sqMNergE7MT8v
CVnhoe9yMwtgqxlAVInaosft2Kg/tvVNLG3GG+v4bYdXZC+ztiKS2Xca1iuDrZVaku5z0zTUiQSu
JXOHDM8YCLB8yTrgtcw91JAX7h6y9QptoidQBdnoF8lxSYgkKvQx1ACh6vb85MWU8MSxBAGfsVfS
Jlsf9tVOwY4bTz1B67O3edaKd+nflPEbP+d0JmhZqP2qNf0QiQWM0Gyn0VVxRXBBBV2q7sQDiVFM
uaV+XwPqskuCwRhidd0cp+E2IaSSbn2f4J40CarLwKp6IwxGxoWKJQqAXUQamqAHusx/rAPG0XBn
HQbhkHzGsVZm2poAb3i7DN+AxiTMboL2auEiXf0diKGx9R/FjmNDIoMVAqKaH2cJuuHgq1cIzCvy
M2T4e4uwxfyOZKJQrSg1gMeDFPY5jkNOLs78ExWBXi2R0axU2asqp7thhk8uohVZ8M0Skzp1UIqP
1YDE1FRHjmQQrl6WPfQ3eHo9Yg/mdqCbByd+oNRZA7LEBpOlDeieW+H5PoYJP1ijD4Mfdbb2wmpS
ZUIzOxDtpihh55f7DjCYifmvfbG8j76owqIhjoD7LH2onOtQVXTuvO5vSmOPmf47eI5SdDJM4M9J
vPwzZjP4BIxn2H8f6jM2sc5EIvkEs9Qv58HtALjpSfEVNG500b6NQtNcbN06TTanYzHZ4sa+Dp9I
4bCL7CGuWNmO50rwFL+ARrwYEBWEEgFVG03c3YI1qW1FiKix5bG+KhnYZtga+Z0IEpkPquD9kGgz
pl+vgwxSWMr8erxyuBHcSp0sRI4M59k5NWNf0FBd3ygEtQnKEQaXPByUrwXgR7nO+oZK/e3iGoyJ
mMo76AFQLY9ouRPW6XcUoVW9e7jg7jGSUiaYo13EIRe0KbYtBCyMwj/StgF6JYLA2/eLjSG2bZnJ
JpjLyObt5ZwJfDTnd7aSjC7SFEocJ6yXFdS1fd/rBIftZntGx0Iop0BHBmVYrrGdO9KIhNWJ6we6
JgJNx2OVemUReqKgCJF8VY3tJbYfo9++9J6xbtcQ6Pua9wTHT6Rztxqzjt9+hLEwpfqpsE+pzHaH
n5V+UWnM3NCqOirGhELXS7U1W6yXorKx0NqGM5TFo8/b4VX9MNLocaFtsz3ruPUR2Dccf2KJPUdz
qGlhkHVoldtzbdEmWoew9AVP2MZuAieDK4w40iPrQiNipqVBlhvr4MQLvjyhLX2ENx5HP8iVbiOM
DqBnxeEn3nIXF3WWVDwP0rJG60l1ujUfHFnhnKsTZYmu9nbjFg7LqGfWoIqWDXeK4BHJQ28eh06o
7j3fE0IEb/sRqetgOMviuOlneLM+iR3CHo70xKx0QAUg13QeLaA084qKEcYMx3sAALtkBEZ2q6/B
vA8WlUBNkDQEfq/Z4IViq5VYKqs5qEvo3U6hmEEVwvl92G4tylTm7FbFeDKApitZQkBHsradv3SI
Ig8hForwCnHnzy8QXePqBglWqce56x+2T6Sww6cnk5HlJ6CfD1BDmUF0/gVah+D/ZxnHy9yMXhH/
ZwFAHCOIMEcQn8wyqau3O8Oo09wZqVqL6tDq7k2nnrUys/eSgGlPWPf2qASi3ND/ONtVH9HGa12k
nI3x0Dvx5h9SvU3q4Jl8KxCS6oEO2eOqsXrWsKSFGWUgMjUUKCzgHHqO7FEjLxyg4XmRfY/95NqG
PUi+zF6M1by3NN/zJouOvVm/zi24WPGdz7RVPCrGFc1G+iJKPECu5hgY95W0yjDoxeaeZh20XDwh
I/WpRUQxFDu75Z5yaUO4qgDCG9TSCNW3ghhPmbAz7yp2RuCGGph0ejTLF5GLV50QKp1UohdxQfXZ
05wr3NpnY2cVFC2dK5WnuuUsX192GOB+3wIS3tExZD0wtB3dWNlvtNSNS9m9bkKPbYW+kmKOPFOW
i7X3SaldSmjSt68zXlooHBtmi0PkZNTm57tdPzUuiVoKJwgoNI8eu/lOS95EFveSs3va9juELKrm
2OZM6V9C6zBFqUxAHkJkU239emH3EGIQicBtX96pAKmP9QM1XpHnILkVgwv2U0IRZVhRObhZ15v4
WqXUWWkeJYSJqqxLsRioA7zJwyHxa98Xrjk2QB8D/bnR7EKsp+/X/1G1J98a+yIgsCSm4VELX3W4
uhej00eaw7ggJGq5D35rKtc/aurbWDdZ7dwzNQtOWq+2KebxPrsKCeCN5XNb5czv8111i95FEBQY
P8I3mdQiU8WqEU9+d3rQS9skf+49nU5/VJaAddGKMes0kww0iYdGt6LRXfqfB/Jf3Hn7cwkdFqwt
W06QwsJzARoV9TLWQJDyF/jqmlityCOLZhwoYrC727mJFSoE1hZTjEYmRxs4wyTn2XI9NyIbb7Jy
OUFWmcNaJA9Kz8JebHxctEcst5glPWSCG/hGiMJIN37VXxqlWNUTdFOXf4q1+vHBmEGHeTYSQATO
cuj87HMt6PrgIPzwE7uViOCi3OXEpK1zKfzqLqX9WtPrNgApngGOdMSMtu68GktOeK7ucyCBvr1O
M+rE1XevvRMqZsrYU0dWwRDJgE6UnUOcUsNVA4otujY6mEZzndqES2mrUoGZYyfc6ZGomGMSSvY1
kphtVvf07dA+AkWsVGZv/YWSw9IzN8jIUKGv1XE1yiURCSvbP0QnLlHcAv4M+ibhf8Tyaf9XNsRQ
Jo4GOL92hpNrGSxlTVtpzTC+FLGTAtln/IpM81rAoCb9T2TGfD4HE5455xeBtrpuDi5qahSeiex1
NIOW3lF9ftUFwpXLAhOY/kC58HdCTIhEU99ZoNmvd9LimJ6jh/0cq7qj/c+tiG0J+bVI2yu6UPW8
lA87U2oib2XcHuPSR7MztCPwlfKjJUCzsql0cH3UNNs17lVydG6ldSha1CusM4avzJdODr4mpRNl
u30K/wPWO5Jn9HZN0tIW/boNoJzRTukb/sttuHtnUthh/PsGeZv04QfYnTj3xNazfMTrkwGDzVhM
BNWke0kdnjtNoGF+v9wVqjPGliTT+E7fNBBRmVDoV6qxki4De544CKmhJlq1TuFNFeEzkvZCbq47
KgG8gaNYU78GpF+ZeGyu1r5FiReKR+/q9LnoLS24ftwGh9U0DCU3evEsPRG48KBCVWrUAapLC/xY
3q+IcgjIACbI7ORGiZ/4dZES18mOaGX83xxSZKJ/sJiswgkt0TEyTxP0QY13L6cdvxyJ2UNU+BWs
MzTov9XrzJx8m8K38apKgWhwvxEV4iEmAXjDAuD8EKH/Y7DSL8Y1c9eSqNijRJtRBj7l3PA2rReS
RrmEzanjSJZ1OI2hU6pCGJhqXf6pblKB/WZMRP6Jp53uclZpnhvYpzf/HPU01z5ko21tg8J9J8ep
tiF45YR9Dt9vs8SYhrQ4MLtdc3uG2DmT5GNqwQHcEesnTlia8lpjBflqzGUdxOHg9hke2KAtAY69
Dj0c7WCBwezgAl+zp2+TBH826NXzumdk/wKg5UF2kQQShHfJPppVQPDUubGY7KttfdBAMduI1ENl
+Z+VhiTd3zrTI7ZKVuUIPzH6PGSs7Lh9ZUeD8TlJj3vuXI9Q6FnnrTPkmVk0IxIwlAttjBHnfJd8
NoO00+S3XGg86Ycso5UHLWSVUo2o9wAQcbpFvxLLt57ZN9Y0GShiqkKYI527ainFzphnp4wuipgG
qlSTb8T9UnqcPaeNyEL2L5+ae9MQe/CpM5HDvoyXTKoiS8zYwPsdmgntkX5kjVu7Ig5Jm0YYPS5p
bC9h8DgkyHgkc6HBS+1g/BpIWppTG/+50qwjEFCaRxgU9AnpoST8VxGlK3UoSr21aZBCBVumRkyB
5MTD9YRUD46UfzTRYlgdQlU8kA6k/6BRFAi2q1smULVB6ZM1S5NniHBCTw0XoRVN5LxC+VhIbHsR
AluovP4uwkK4qhQgYSmUCALAMSemcf4zAIAtVbFzMGWbl6j4YOMimpExXNihqGhWvQbbR/RhbuPp
S0AVehanF/jHwdACAWQsPvt9WyeYSNiQXmbHw0AugmUdyRK15jW/lrAIZjehh5a3nVp9bD0iDoCg
7m6r0Hoho7UWOd40YJCO668RX71iKq2OzwbwuU5U5j7tvVHslrEXWLwSI/THN8yxQ3MU63VXuaWE
aLBoiLWAnES66zyyNrkpUeLscHGrxe+E7RYgNGbFh/zCnExrsiu3YqPae2LkPtK/wxq6LhQdFDNL
R9WXe9o29Jp6U4jS49bjthJh7nAyi+QpKtjKcqjab/oLDGEce4B89Fvn7naaq3694zLuYjI/mYIZ
mYb9Nncg4nhYjQq6rGksiZQ0ZmquCY3IdB2A7dnJCLRkeIlKUww7kSfvCr/EW5mSnLLPmaUPlnd+
Lh4JW9q4g/SH8xRCX3gnqKq5hZ9a6dwtmiSesNNbvxt0fjXKPHVhWD1EyabL03r4P9Ph/8R0ZakU
lKMnuLCbC+/4TF8b7EdoeNKBZflw4EPLbzCBkfaG8gJr3GaiEKBwJvUw7FljQ8aCDIkdMoV1xVNL
/AN6CdqL3PnDKGqeYUFWDHPBUeT4PBcC81oo6A6JuNUU22nCEPt7+35uUEbecqFT+qwMBZy+3Zux
2eWxXq3D9RE3uW97gEydA4zOHhFDFGteOMySI6EXvtIsnht9MYH7VFJmTjSmBe/TM/YV5QQgqrIL
Y+w2Ly60hgdPbsPKafH6fIXxM+4eIWcNRxB4aTn5Lp6XDWsZzFLmgpX5vT3yXKA8mhGnXoIHLhWa
aKwAbjTYMe6iNpogC4mFsMoYdMk3RLiJluAxjlCxzDMwIloGM7HfURTKzW1ea6Vk58tFeKhw+/QI
XZMHuo5JPY2LV9LwRDyVU32egSInH5u76nuEOe4z2q1jiL+nbwDfS/bS3d5K/lrPzbWHbw4bMveg
7n7C9k4bRbNvieXJf5xbK7nsXmcSrRMOsvR9zbBxKV0pGFARJraivM3ja7ORoeabOf+PFAOn0u22
rws7fA2a4DVwN+540QpiuEtfSsG44t8j40MvNdl0+xlI5J0LsiDjv6zFEKTmeZssSYyNzDS4L2yK
Ir0T66/x+JG9koed+NYWWRYYZAwIMvkVDzbtOQg1UK0wPDwYnRg6BMNKuqcN5iEVAo14NpB7tZx3
J5jglIFx4YhyizAa6WddrYfnxr4YX+x+NwxaRt55i/pvXUrq9Dititz6Zkak5HhfiwiGsJ+hnf7n
5DNXY5kNiDET9MHjo5OFwIX0wMf0wdjfQ3SXwD9sPT+UWlY7OiVoqLbolsojajVMqvu8r9LO9QGH
YhCA98OYu8wWttMb7DCHJAVM9qHAwZZmWMejz08X/QdZpflyyip2xoWbX9V6dVv+dY8FqcmoYWuj
i3OMhM+YIGw2H+ht5CGEV7+GMGwLLilvHBjc2Byj5Q1Qd60WnaBuTIHBQQn4g/zglzzB+2MM6rE9
ub+CrNSfvPBp4cCGpKdUOvMFAGnKaGdTrJeEkl9MVCrDtcy4PsGjsyJJqC7G87pS9vZUwVIo7rKC
hdSOZ53fpcmJnrO1LNUG+MkGBvQAaO3Hup+AWx+qoQb+YoZOirCoyCf29q2a7JPYneaQnr+XSJ3a
nYTY6CXYbM49AkJ0vOEzbasqHezYMvTX1urV0N5UhUsnS/wRx4Jfx2M7ZILO1akuJv1hadNGw96e
3RMIi1+FRxHnnSiR66SGLcbgayWFyRiWAR66Dlb5Er63ZEvOU9Vv8jzpAcUQ0Hlq5pLmikE0lUvP
huVJYuq3N7Py5Qk3xyxfPVAAfJVus0gdYG6s/F0+igIkLsIy2hdafrjnqg3Yfb4k3e1INrxG6n/c
xSVrLJB4D3sIFd+CZQB2amRpjGnGZ06q+4/7uxScstpN+Tdl4A/T/qYxukx+HrCPGxktaJDWduXO
V1OmfmKXDq7K79HpTkMtj7wC2EzGauDHnFJH3dvCVgD+PAMt4gK2wOYRHxuqS8lbhJEJiMUTaBHj
oUBs8dQQ7njoVhWDHGcyZxFKx+oRupRcsb43QQIJzYEu2G7NEACVOvgqNZvTepYeIECa7/suBXCg
fVA72+RdtViot/EYeNRRdEH7r3DqUiMRd7952sF4xEh09XigdbohUCiEDg1Hmk4Z7Gnpc2PhkE7m
P72fEhJH1uYEYTcLqGJthAg3hBRInfGWSiErN1uM1unD+5VZxfo+JhbGlp5c14tlG+fVtcfibzvz
IjK3qwwEsMRyc++SHHfDD1Xok9fjF5INSNUawhvE5amD/s1Npks52blwr+lcX0AP1eAE5+R/DC+3
FglvXwZlUnftCZX//x1k/p0n5DZGGvsavdXy62Csznn/UoFgAl91aJyAQI+CD/2DZu4piEjIhOmb
tUxMMAURZyVu3z8ibOX/t/vmOmyjVKRsCUrij2XbmtZHILap9hxqvXHCb/QlaRMToa3rJGFCtPvC
o8NyIMjGu/FBSn8691Qz9e8xh3pB+ijTIa8Vk964WMnCL6z7t5E9qdqNqVQ2Gkw3zBP86zoYH94N
ZbjMK46NE3d24HgGu9hDAa4vyPKLhbLZ08qtjgakVD1O3q+fQ41y5Hw6bEDiWSXCeGujVfhW9E1e
c6GyDivKfIg7VVU7mTJkxCQkExQiwcYt+YNkx5faqhV2X8ql8XoiAvGwb7Y36nm2pQOiYvcjAY4S
fWnUpqxchexj7ia6YfpOiQE3UTFpoGKdJwMRjMmKn+9AodRX/En/DTmhOZgLDGofVRScD+gWs+sk
bDDpuFSjpKH2oEbGJ3s+mJyzMsAuhA0aLRNQFghwK9lYcRPVZCDPhdsRCgB9ph4YC+2sm7UqzZHz
S/tIfFcy5UOCX78unrRsxyx/mmdjrkyI0mS2iILSelfXdAVSXA4VY7P38wh8P2g7SupLi9oiqOL6
tUEz0aBq4BQA27+7M78qdQCY96UC6av0rIXR72Gev4jTe71hSGLoXETtFqfa/2oPVhlLWMZOcWSX
lr5pKRlxC+Wy/OiNR25z6ETKdewckYI7ZBwK/0KeAScO+9hw+Vvcup714wDAbGkJtm9sceaNkrvW
Fm0MhIsqUl06FMcR4xlt4YBz+FJH7cPghFWP9OYvaQmHnnZrRE8NBVm5ngpGiAKZ1psLZQLchBGx
9NxUGtrFrGram5eP+JjQgZdaJ9JSyYFrs8B2+yR2QP3iK8DH7Ea8RNzA8GuaWLaiCKUFFJusCqdt
WOzRmuglKIB4vjIdjx+HjZmPI0AC0WJ+pDqS74R6K4zWwqV1B0Wk8+6YxJUem+ejX5Ttd9RJOZFw
DxdtzUDiQxeSWgIJzdq9eDYByPBOjyJ1o7ET0QMzAdn20a/wNfvnUbWNa88MsIj5dZzw/cebl142
vKeslyUhSd6ueyMf3HgB9xnycNfauuYuhgUlaIrd3TISnuIot36oLURURx9gIAApcQ/GH2ZQ1vlp
e+oLcN0+rJrmKMp+eTIbGlS6pVnBIe0xmu8YwQXMbZiphXojS4HdZAwBwqmR8C8tVIbtgPdO/w8J
8D6981E8BZuFaYNVOi0q7bcT0+WENvGl33Gb5rLgXB5O+AIqg/lsHqWHXcSTyOUeWZ+0LyBBQh/Z
Kh8svVvIUshcaCDMuCh6J8HD7pRSCCSjswW/I55xevY/tXO8Ia2PErKQk6HQ8PBlB00M+8UpoDqg
JwUrDJF09ZHx63/7GT765ehKCFo6/ZfY++9myjR06Puqq85pfGAQpj/Qg3jeaZOLkacOnD/ktDs7
ODaolsbBajEb9C1Sy7akm08iPRSmlRb+3EA4+2HA4U0CP38KTqyFwV8qwR6sOG89tBFVGHy+m9PZ
dMsPY7ENU+17WSSoGgQv0B9+D1HqKsaRIynd6hRkEw2C4JfAxROjUhC8ZV+dY85ZpH6JL7mN71Ig
2OY7WSkiB+CmtKMwK6Lc+eWOVJwLScMYQLAFdEKyGGM6GB9B5zmzEdBRwnX83XG07PUD1mbasnhR
rZyPba8oUE70YBDcLSILoLhJXE0niBYGaKOs7Mb7WYiHfNZUghQHOq8mjpIw7cRkE4Cw4vQAnl59
kUeU4W6GEMTzTeqAHuT7SffciMdqGG7n07iXqOWV/rpnRbJ+95yDrj4rPARcT1EDY+ZcuSE2sCVI
x+KAjo9McaTJJhx1qkEXOmTzgYpAYejtQnWTRlKGopSLDoj2SvzPsec8mp8uUI4SbmxBT1SE2Hab
I2nPSybQ0RsT16sGGKtUdwuDZPdKkkxouu+quVsiv14VKcWnCHdKoVM1C2vVm4dzDkOlSssprwz5
CVq6pHoD8/b8+wp1wKjFmWCw7RJpS2b2XWABOhuP2iACdF1YTfBvgyzWZOuVPuSpyOWlTyQQAnwU
OVxsNGmK7P7z0Sw25WDruv0y+kA/U7dF8xEunTYpl1atKPlIWVfY1bChvvG8ekIMp+rc9Mk33sOU
TK8u4PWqps84AMTpIhDDI6NiyQUi7lmOTwxOojF8tYPL7LEqxXMXlXx6bVHG+eN8NM1xoHWSllfC
R1qOZ/2amgIZdgRqyb9iyhbAjcgtnM1QUB4ryAGlTRwIZf5I/zH9+igYoEwvV+dfiiOpXb5VbJxa
m4NkBCSavnigQHhuEGyBa5RDkSbyWHS7PyzPpi9zr5bNb52ENVVR/7qDsfbfXzuKF6mfJTD/l+4o
q2m+ZeRCjvReWUKPsAEUVcLWKM9770hb8Xq64pstvZCqGS3/bU8vPGVN7DlK5NDEZcsl/k/iaITV
kEX9Tcih2KuI8QCVibvvEbo1tbdqH0AOklWPA/5Llziu9FidvEC1xICOghupUdZf5ivXDXGxOYlh
Zzhp61xKXQbd5YcWK6TYCFubpSzko9AU6FZIagABmksx/o1sV81I1q9+88pHis0hEUXJ+rL4fkKa
qn3tmZ4OmmI4lCmbuzda0YtldCbM117QBo0zyYRDo665BV4dmYDpkwUhiChU4knOI3H1Md3fk3VP
61YYxog25Zzn74NjHTU5yUY9M+9+yxYog8qYxFd/BwqDET7xqvt6CBnz1HVVVcnUkVvta51Vmund
KxdJbOSj30pHfjodOVfn6Z4/7AGY64FCDEWPCoOIcowOpvEtjKEKroDVLm2Jlhd8Q4BK/lWOWDs4
L+7xNhiy2HCMsIFcznCeDZhCFYALLUh/F09yqeoNRsFKG46JEdNkx0cfXsbYrJ5QF9ZtCofT9+8M
ZzB9AftKVAIjt96VTq0EgbAsvxJpJT+tGmMCm9Fe/BBvamTtY+sFSnFYFHuSL6FzjjwNCaeQQ/01
8uGrLU0DmzZGS2tsa0gh9L2Pxm1YYq/glZNmUCFkR1ErRcA5tm9avFgy6ItiKzQxhf99IowZMueX
PzYWOIHlE+YKMwXaFFwteX8mRLzs4Wqr01EarOk78kaDAgkwG5KO38J1vI4qQbbF85dpy0cQfXB7
Nyi7asIugj8Db52MmUNjsTFQ1mWFvXLZ93N8gUU4eq5FAKbb4rwgPq/3K3JqWo41CfiweXL6Pgkp
pBlvtvrDK4pFDKuJQH9ce++3d8S3jQYGnUcOqHCovOfUrmrGZjA8aEzigi9OXVP2+kNjFw8gTEaS
iqpaQJyZdhUR1MY8XGb4i75tRNYpk4oejLBHNBZDhNli0zCmxSNQ1Wh75OSXKbm1LOfTyqlhdt5M
Ynt0Ny6GIT7gtj4la7Cp1y/0Aea9qPTPUGWiVttxwA/nOosac5MFz3ZKmQxMsirds5JQ+LTeNajY
N/MGImMPqY3XBt7tDe2EKJGjceN/CRhpEp0WcjcAWmUrJoiZNZIuLBtOmHvpR0Ao95iRslAI2yF2
Fh1p+21EH8EI+ggtXJtYfiUOtY58E9RUxmfnRSepvnlFExtqImc5kfUxhncbYEg737TaUigkEQtC
H3WfK0jeMhTFgcO6aYLI1idChi9I3QEwuPBC6oIqVE2VFRT8+GEoJ7icI50J9xkO7H5Xl754vTkj
K2sHxNVzevCi4ttIompiXlbYRflDa9DBUMWIQJ009QyoKx1H3llaRN3GzLpjUIuBcevXaSjNzC8Q
kV27DRW6F/B6yX95RL8Z9fPBfsCpCl90g4jzaOE5lQwVgGBDloYFgISSV09HhycKXO9mAVGRfr8f
ftkD9qSul2/Ux+MyaimLxtDcSngsWSOpf/AtsJs4raI+8f/zaGfcpMy7lAQFSeaiPyD09KEwI49A
mfQdkscB5dPHhywVMjvJJrOsvIg5u4uYqrnrhmyNE6qamH7dtl5k4P8f8wkBhgO7xyjm/Rvrrbk7
QvZfPz2FX0sShZkxocQ6Fuci5KPcP6SU+kE6SYn/CYd2B68lHnzsrxGus90dYE1kusTl6TruCVsy
ZaDlf/SagG3Bc5k3xBLLGKkxkFwFTMnLmT2BLpeCvXMb3bAoD1GZ2MqQ3o4R3wNXOgq5DBJR+mWU
EPwhX9RLCBXo5WOCWsW8mwvYSvdw+ulgmNe3jRa8KlHKypr+mjCQMIIkVZ1kXZhOUxzb3anzcrj+
ULzC/CKbR4vtyPUEP5Bca1GH+CvVk1qOmudDmn0dRM92UR7L+Sq1PQoWyu6EPETN581GpSX3llmd
Whs191VRMH7IVLXAAV9BzZKyGlZZ0mOAdRk1dVPUHJIAZp562d/sv+rh8ng32V2Um0OyzAcplj1h
eb/xYtdf2/sndbXY5QsAACRBrkkZjf5LKd5SX9G/CXsntNGDjNIuYYV0NvPlj47d3Ldz9MV+Zjv4
tzCLxzu07fo9N7GrJ2XhSMx5KDgaEZeO7HNcN2HLv90EWosfwfN7PSyZbbawtKHDqXrmspBJ4MPF
VdfkPMf+n9oxpM7+n+7pedzYZb7k8OWSw9w/OeSFyuTAFemKHi4cv4J2iRNaeQWLF45l9tFHZpb9
V00JDhRJuovriKcIPTwLhOrp/09h4z4gpMZsgwaTskPGRtqYh9wK6CjVKEq9+aaiVeYdLjpuvEZ2
szQ5gMMiJ9PArm2WSYn6iAazNTJOxLiMElQbbVl2HK0H7NG2CFlGg80C/DObYLjSW9QZNWpugkQV
RcAlfjtsEWVbDtq0A3Cdz8QDFJeftaMS51hJ2QPxsQJRtRt8gu48UD6jpNmiFDiv1DOv+2P+X7lD
LhFWUekIJO9izpSUwxgxoAWRCThBFE16wM09+4/m6RYJWDgy5MDgh5KamtbJA0N9dstEJWjhpXPy
m4k6iC5gPcnU7sLJ70OR5YiYU962YQDbnqRYJh8aupX1eioSTWPe1U69DcN8pzGwejC81nRb8RbS
LSX3slK35iFH3EkKXRz3zxuJFTstkY4/DVCeOIqVcTgVJTq23Xnhgj5zAjCK8XC3Q1n5MDeJjcsK
eXrvHjTThrI2QxQyJjeAFyeA7caqa5WGEUw5GjQoRhEy0BWOR/11OOMVg5OuUjOOfcigNzOCD2Xk
J3dEx/ZEX8Y/2LOn4q98Sm3Z7cDXaKAbmsJCaAEql1Kx+hBOiOZZif+eefYPRecs9C0nJ0NXsAQU
q6eUwzhsZUBuAg90Nmp2qRY8rnqDVCTHz036rGrlBSPMTlGElPaITEi7FY9Y9ioeYEB0KjSabRh7
pjub1EDGeIKMwd7zaPkXkmjBwDRVHcatFTv/7zzd3fRXZjpiIwehb65tbFverHBIFgznUkRA4/nd
iYuJRYDdhglUFGDBVidl6sIeCiPchwn0whxjLCZ86u1wJjhoOprpFLssw+375L3sTGP91WSDS4WT
DYDLcLgVOmfwPu1iwOPUJF0s0ZUNN6fBwTd4YjzEhqmOc/nPpbkNz+RNAfwXO8m5JyGYSYerDawc
oU3XjnfEXnhlGFOaXQCjN1d5eCmMoWyC/SMJ8MMVdg7MrhMzgLpwESJdGMBPcbmAIEX5F1mb5SZq
ahdwFLt1nsE7JRz0ubGQkvLu8vTUHA+yAJMXx/iQI12D6fH6C1+/ly9Mf3Pj5XdXB+rJfiOrZ7zv
PBgFA595Y1t/ViHd3xf07M6anMAgMC9164G6/AR3dgDIkhjQ52WhfFKq+bN5k4TMGOlpGULVEcQ5
FzbdJPMcDuvd8xi3m6sPb23mlI9TfGwQSXeM0xugafj+l09XSoN2tCV58grlYHRGr8lQ2rsd5jKq
0JFWOMz2YXl2f42CV4U0k8KfyYHDwykNr0Vt27Tn3pwKCbWmtc+t9L2uZL2t64vh3hlVONXFiMl9
xqLyho5hdK91bQzlZ6NOsrcnbSH94iWySabXdne1LSHEZHNXFzOhra3UcHnXnpzeAAH/pceD9wLG
V4jeoUPFqai6xYOsz68HNXSPKjaBjU/T+D7ijXZ5GNAgZVEw57TRlPqCiqFbm+X1atwscPXMKXjD
cZu51TH+z/rP26ZX/u4teSOtVR4xao4ClrDgNTPoDI6k3P7SN/xvZdHkTYiWp+HUfkcvScDQTn0+
DY/i4y/B42lwjVz6mNhOZg9ZE72Fj9qsigtdTpapqBbe3xs1MvT7qBDuP+Jmf8ZKgWFKbmPLX2Kw
P5JTvOtxUgT6pPDZw6WxObcgmomyLUNFVG7QItLMQrHucuzDLJbDKsyNFm7NPVhDU4fLBwMQtqXT
ft91PJneO9PyxLNedQnXqiLLCPE+SD8MSeRhPDIolrixsjJPCCfSuS/0Y+JttCJWpEXOET4gkxum
M0Vg9jQnmpZJCxRbgl8wv/sgk1kF6Ylgm0gGRyD8s0vfuAoDyH3bsVIDnXvb9xKSDyaS5u9PDug1
k1lD+ipjVr0HGJOFcC4uOXPPmj8giiH7/kg/4qChsFVPR3exf7Fgn+8aD0EjxUgZ4yyX4eEwbArh
BVkm7vCpVC+crWxqDWjOI8skXrvTcgIyYmlsVQStCSLzwR8/y7kGdSWH/PJT5OPu/RP5Vz+QX+zD
i+Vqhc4kRY7jyNEP6pffVN1Op3zgFUdTH6X5QgjanHDrJY6vrP4+9DLD4NGNxvtDqUZtTkbLe1DJ
z3RkmpOJhNnLvbcv7Pa0D1MghRct9mltMrjCRGLR4+udowN8jdhur2NEcaQ8nDgf8daUv/J8Y/FH
YKDeCyB3Cu+v0xpUTm1u1t9YmZd+38skfJJ3QH6pmGOUNbicSvmTaGumVAwBmx/wxYlYv8cXRXHW
3IaJwlymh6ArGBL2SuMVZ+w+C5yKz0Khl7fx+oex9jiTqV6I+nfWF85P8U5jcf2fpA1/M9gH0DiG
nZ6Juv/F6SM6jwyU+RjFkAK5BKhXLXooq15nu1FPrPYd7qNY7X/hXyhkH2wdCmn5crbXfahsnM6n
/ni2/i/iNrElXQMLGeO6LO+dzId3crCaU3PItx/DvydQD2fxJkTxuy82UV1wxHYFFmz/gJ/8FQSM
0BPLSo0CYaESQWGqGln3EfQ3npd0QOyiqAp/6inu6nmtWRBdzLxR1p6/g8HT0Fu3E6fPm8dd17eI
UrDottmq/ZIpghh3xSJ6eERWdimGEkrEET03H0aS3TEKx0HZKKAbgi+PQT+iejEhosgY+BWMXtO+
UjdppSWOixC/+hBMMcXelDW4U0sc9tDdUmyvGpAFI3XeWF9yIQeK4mQqhoTC3Z7oebl9VDrHa+gE
AyZAQZxGxWJWGVJwk7dBf0BkOK9D2nab6qQh0O2Ugbxv1lhPXABwFBbNpl0J1sW0CFL1vnNKhuHW
MAiH5mAs0WGZFkazY1LhzcrPKvFERCL3dDhJp/DR5bXL5uenRG+XU7wEkkFg/jAYudD+QMmNqly8
VL/li8CpXc5YMiZYvcbnvsJfbxU/4+skleyws1FHlcGwSJUbSemI85LscpcEKY85MHUkDY1mMa/2
QuCCdfVe5WVWTIIdyQ7gO3CVIqBgJEhLnOUbvomGXYe/ZMQCHk8ZtvfV5vTvsEHzplhRl+dQXCNC
qwhq/GvdO/xZfxYeTFs7tbzdsoCIBHeDYnBOyz7sZTiD7M8NeiYqlcIURYHeIgaEvR+bzPW9d4A+
Fb7c40tMFxfx+ES+PGTkpqv1HvZJ4bFX8O1Hwv4TMKRI252rvjWWfQSSg89CmpjejcQEsqLrr5k2
mlt3UFVFNLOcOJ10aKLb6PZKQ+sAWwA8NpE5BF2PjI+5bXezQ+WEqAXEupjiRM59HIRODJ+9rNjR
UihrrEYZAyqQLu96mfJr3OL6eOBVEdoF9QIdRtuay8oYSZvtaZkUcHoBfBABUCNOeQ2SrIi7kUnt
BeGbnv8LxDBkCOmEsbbSwNAYhEmBkChgSCiKCnmatSxaEm80hI3mrv9nX1XGg2Yur94Hlie8n0a2
awFJ+yl8au5YffDYqPBlsp1hniLB0fPK6dNvMo46PWX6mSnw4Bw5aMSIlNjqXGsm1KTxjskhAt7A
SaOgfhNANMDCq2A4NriFNXNrlDpYNLzMS59J910IkfKmvOhy/MrFZLEHJSiBdFtpHe1sdzORCjCz
lbZ143sb3uhO+XGSiv3z1uK8jSn2vHjFGOJazaL5jRDar77vv9Vjxj5uEZj614JyYVbY+eNMLNk6
0yosc/GT/Olq5v1ip5JT/PO/239pEH6h+MqvZkxQEzDg0EFPQCo6NIIIOZg7ZAT6rfUByhssoaai
ZJhpmzM6e6OT4uLLNXPRySVuI7WelvvRwPSeMdLfUTu7wp8IaJD5oEpXeBBaptlEIzMJ1pEJWke8
ZHZaYkp3dZaTs+QFOzymFU0Gdjhh6cWI8FvuLw0erTB88CvZ0t0wjfuebh4w3B1hCxHDmGzjE/zV
piSeW9+V6g/3/P+pS7Xl+dAqvbD00BA9jt9bp/T1dlkUaKWBV/yeT4mkxzPS3RqfGG6yvF8QgC8f
8iVC/RFlFVJlB/HBNnL+BPvejauh4e05az81nNmKPZ5BF4qUllDaKWR6DiRM1VltEdd3CUWb0lSr
qgI1ODNyUYaziTOYsRl7FhQqGfRSXM+mKjJFooOHx0a4DL587p8W8UYIev58SwsJC/vyNevlRaMU
82fexnmeYBasjoT5CMjxCFCVVTXBLNKQuuBP9SN1GEEFT4cdU6A0NZjsjDSWNPQcdzgxg0eHMuyL
IpByvkOXFO8hNbPV/DH5G2FBAY2rknBFCb25M3Mm1X03xTsQQO7098rNUrz0PQMvkEtCONEEAn2K
DQvrgVRJmTjAS2YmwILBOsPe8QFRHwfBFSFpoP35+TzKZacLMyIB0X1qr9GZZ4Brhj1RvR0VjsUh
JJMQLREQ1ddnFK+HneOq+epHGewyOBw/o6m9cUHRwB9E1Wr+RJZXMKgv5jnVCioeHoxdIQgnxWdM
O5sUH19rxYL5lRMqRUihtE3RVe7uw/NYyiwv70xYXkvVtEYg1xwo7PKrsQDDY+RLJQwDXkOYVPi3
kNwTSYcHnluABZHrshioJnK/K/9Ko9hbKweBoyJ9BMhQ3anDY640Wbem53X6mys9yK8+xL25KOAv
sPYd394dTajgagL4oTiyddRIAIRDK5kC5vlemf3oAHk2ldx20U4EpKqbF37+mMnmOQYKZTSxdlUf
lcE8rLD31p4Crhk8GBp009CWbkVAhsHFV1aM+BRJf3bUSbV8ozt3E6SBcvZa1HlfEaZdmk2qb+0l
0iJQWOVmd3jdrES4+ZX8q+51laH3ggR9uxVj9MvtKRHNOTeINICCVllOYyiaM5hDOQyZr2Ii2yrk
zV2U/w8MOHvY0kB9SCx4cN8ekdXPOJS6TkR8dZ//tZN3jvH7e/ueHUWXVBVU5dhJXKsKSjg34MqI
3+TWMGOBp0/HSN+7QPrd22gHm9yMj8cyPWGtvbONYvzlSLnbPLlCvydhgntz5MIFJ7LOfdRLqEsd
qiTFs+7DDOgaWgSPZkilhrmF1HqXDLozldXyLTdUNwzeY16I6NLE7q/FdC3IEHa0AEQ5FXYiVAVm
qgZqxUJj1lyBpYcnQo7fAaIes3dzHldntE0bjWu501J4grVnXarlDfXRNs60CwT1xTRWqJpyecoU
w11WHLlGczyu7TqwVMMztKXl/35hgenCG9tP5SBXyLn14EAVi+OEYT1aVi/EKhapdY/Qno2BecHz
xYjKf9505vEMYya/dVoi0UJc6dBSa3zo/EjxOdvLELyy6pY2ZSM1VhPyZcq+zph8rbW9G5/s3QMl
gAFIOExwqcDztKX+2G/16J7irFPviP23dZA12r33KL2y+0P4oflJZ3lusGtfhznkfbcOjkIriUIJ
6eijfGAuaYy/KJlg/P+w7k6E2iJSUcdQlQFjrLyzxFjf+30TP+D+v61NjWivqSeBZJ4r+rcOO5nd
RKWCbJMYtRUdJrnBB5LswGWJhoAbaDkRHiaqZsQIn9IpGaLB9dB9RwxO1TTT/tnSOcfHgAZo9kNg
W0PKuzvsB4h213DdLDjxhaL0llrs8ixCNK5W9rZupU67pKCoJauPe9YC+peLslds31r24SZoZ/ge
6LeyndbIEK3TfEiAQuBWNPysz8KR85GILcdiS8fuQZmYowHGfkVQimaWP3yen06jk/g76xoKwj/2
albpXnO9ribwv0vG9+d+gDqe3Rnt3Uds8MKbEseXKJtcy3qYZ4moYmFLxGCXR8J4QSx0z1wnbYt7
b1HbRoqO/YnZGXwkH0oajm7WGkfdUo0bFBtht3gic8CQzDwkgeZuaAaZiNSieLR4jRNXHzcwplYH
dTCQlY2lxcp9yIhy/Dv/1TgecZKbeCkUFAu/QCS0FGnOOnKzGDiqImGhPyNhbMw6Dd4meHSwLZAR
nrq/6y6C7RyxIhXVWN/ErGSV8d5idv+H0Zrj1+FYhCH3UmAgTtH45F07VkSSbGb/KjJj7PeYaGBf
+jHRG+MMlpOT0a5afo9stPylATp/dCmW+LeK2uKAvMCNpn+b+qeTbAUq6GMy+PK1C9P8MIJy7nRd
PoAeBos+WFYB9caj5d4LxlxhxX7+oEUft1yGg4gG+bfrtZxNMc6xXJ405dvWs8Rn1FRDyARpWMzt
xc6OHqlImiZxANbUlSOf9u1Umq8e7gmfc/W6Zq8rS/Ylw8PoLOI5PPRA1SHJO7dHk25tkoQlMHI7
HxJo3IbhP5LNjTuR71lInmgOHng1VFcMpUtlqlhDXtKGzztUSMMB84IxvzleqEPqlunQqzhu6cdq
BUUz/9mpE5QWBAUFeu+RYKQlcszMzNlth9nku3wOCNb8FTHZkmvEYhoMV+Q9IGxV+poAIgoSXM+H
XIxT1rEZ6oxxfEhZs6lj11mX/PZV73ec1RrGs4qWrDzdDaaHP4Ohw03x5XaWrnVtaEStH8b82NTe
vHRmd4fbqvD2sTLGT3TrZdkgj2w06xcB4nRC9oWtm6+oJdWQU3V0t2yfaNjuX3dGOVakkdwSNazg
itC49GsUa9FVuF6gn1LEfCirBwBWel4Kw91EQ1UZSIDfd8fMcRZjTPJ67HMCj6KBmNM6U8m4yAzc
JEuSI3FSR5+IQqkl9HqIs1zg5h1VBxyLv23YzIdBH4ry7b+jR0Ba9J+NCL42RolEKP5L3fF09qcF
NxaFKtc9jz4ybAmkJNlXIsY24qzL4kzGZKaIhLLW9e8GNQvmzqJnjPf9gNTtOMJkLqB6kuWogOxe
bN0Ba1p/LykMZyx5ddgyF2hAT+jHTzgzsd6GxZ/qpryIMx15pzu79UlLVHG9mb/6zTeNDAdEDQ5Q
/s11KkmzkeaDXgvePZhmOt/eq+0dlakxFKO7Vxms4LRopplZ2t+iG3g0L1f3R2qXhrCE71Sdd5kx
zc3WtEktcoT5g5LTg4rSwU6wdqhoE5qXb+3FvCQRbC424KYXjIQrs0RlXG8kl2BHjZvG7znBpujE
qYakRV1GCg3fdkBt7S0bQOwbnX689VLw05Z9ULp2XzJLMn4MqmXcIrDlXQ+PZodJI92MGUa5E84i
Kq7+rO8xUsBweKK9Z0QxDl9pK0qNm2Pzd51ZlakZPChTlf63/CBZVUP0RFPX66ZmjivJ9n37OkE0
DA/abYE999gA9Wh9VB74CD21eVguEFfCchgJyid/J3FGWkXkgn/c81LH5TbUq+dLudoowJAX2ydI
yCunJsZQR8DerQLV6L3uMpPgFMv8yhmah8W+sYqlkgtMdiIB2Uz8PCEcE7mZGNfjubdhJGDoxQQe
/SDx/Bh1RY9gzCMxPTrRJQ7ImM/pRDz/LMbiQqVJs2XcTAN/te/TkabVcnYamKK/Srm0k+8Ltneu
OlKfMN1pe3bDepmlIlrfvT7/m2MMdsLkPSeGl/sYLRi6kdGBjyggqE36o9Zff8ojyWLPOZcxIu9k
+jXYqB8cxw9TOTArty8fYbqWi2wZC6M4fszCh37onVLkKnGJMAO5kb0oPNPIxqL/3LC1GTum6TCD
uPtccqmJrsUTm7vRVxK/aSldPrkKR5t+HhUpNBXe3wWF/iIhPtD4U1ecgTHIvigfJDE5ISky0wjn
enMgXEf5lzUUf7b6Lljyahhf6hBDsU4TTz04k0jX4xJlWxP6FbiNd/PDTzBBg+e+EJ6IaBXWHdMr
ATQHsDGimXH7DwYfI8UwCMzZ8yN4oDrrY+EJZkPd4FgEx/9vGlOPYHfjTCuAhK/lVtXQfeTWsH1L
KN7FRRrSttE8nWnwtGk/xHUXpgcmn8oxU7UhJFjJlG5UZqZB09I8R1CNC05f1Mshj32cGZWBZ1sj
yxwp2ZU3I1DHPZVEO2zrY0ziBhxCwcjPGvWNpvoE8MlV7zk1JrVgsENo+evjqa1aVfPvTTP6i9UG
DzAJP5sOktl5Mh7ByKUcwzLmDBg4zuc6QxoKsepZ++V4uBxmnHMWSscLfrxQffcGN96CYG2+iO4U
XlKrr7IfMPc+PHNByaLwQK4oXnsuzDcADmE1O16RIPlR1QFpxkWyL5IgVUcpkkZfdhLO2pvohjzp
1PDfbU/sk3D8S9+1eezglSyMAaG66+DI6enfBpURtFlBY9X+gTg8nfXwTfLv6wTzFKeX07hUz9G4
2ZuEY6gHy94bUHZTK3DI00PDkuBTR9sVevFYbG8OeS62FawW1UNbC8F3y2nZ81yTXMLG/061hHqp
3oz9w9vcas3aSiFBspjiOMAjyq0whI7fyu4ulQlbSAt+0vPSDLKE/DjLvHQgwulEqYsbTmwJAuBD
tKkiasRM+JkKJ5pjPXz5TaPK01SK99ZzvP0z+iTL82bmc2x/nVUA0tVaAf8Swz5h20oAV7r/swjn
5FWHkzNwSIDOIFoPgqRBbbStfo5yVVMQq7QgGZt0cn3tRg+2REHgnwii8E1t0rF4ShdLZtdXS+zr
y5YRO5imS7hyJbtYKaPd0yu5S3hlwsSSOZ5oF5DWMvSCTc3x/UJ8dQAIKq2iOI34Ubv2c7gTTRSD
F/ARUWjQmXzJyCnCVITC17zB1SjjLWiHVHzaqUHNnrICIo6vNqHSvhELEe1jZPrXcR21nFD1wWXB
9Jw7toyWJpe1m8GUd18GIMlCv/bpWGpolFBwbj5Retedn4XsHlxlzlBw4ukvsDCZ/f0G7ClhEe4Q
6uFTPS72eKIycjDuKY0i20YpiW0/I1k6n7H2gQe0ywxujZnWlo8Z+HKsK5OxhQNi301IPu4OhCPT
N5lz366sertBVF0CfK858WbQg2RTl/zkVcZyzScC4ejjsJgvH+8ZlPCwOy7o12Nk7tcYizXBCYPH
qOnUQ2hfQbDRuHhvhvVOJajRK6NK1UATdmv8akw5MwH8jHdKK67efQ+xgrl4BAr8IEd1wX0Ht+3R
5g4bhSKEgVo259I0uHLe/xfxBc0IaAovNYa6FvYvqQKJoNkOjns5Y+56sk3QJlJvM1YF2l04QoLX
p3b8dg69Tw8WVg5RFcyU+PJ1PlJp6mVtWrkHc18zTCNFCZsrc92H2pzn+03ZxNXNUQJYz4GIG2Pt
CS+fbgOW+L4VuFsTeasMGTQbAbcf1uW22rM6nOBn68Z95ayiTY4H/8UOtRAU7aThb6aTEnwAFBZa
Ut6wnmmWEa62b6J2ovVj7iarW15dXBLozHLIecpm6AtRJZyXBQsD0hyPMHD4yFaUAEI/9+rsQ07z
zP+bCl3R82bzMWsyUmyfjJSO85xgUgoaThNBPiKjKYqOSzR09fNeuHdOkv/CukEi/wEVo0dqeZWA
7aXL0hzyfIFK3zOSTaJPbguNXJYWtOk5YW9P9iR3IYVhLUtsThPwaU03r8NQlyKyEo950nd8Q3uZ
Qmo1CfHx3h/hTxMalqfMQLKQyzgUMbNEL/CObwUpmWipZBomNQHUEJSIuiKtttVzYUVjVYb0Tfmn
VUZrnTIApQkRUVbHb5UYMWZ0V+Q7IloX65fVQnYfTlakyRzYk/dRL+4adqd7PcOUwAPiZCnpOyoR
qrSa7XV5EHEgVcfQCgi5Z10/w/UsFjJLtTLfOyg7QIC4Ir26LerzdJz6dVWjwAYdMP8w5j5eYpp5
zIjeRVXNJXSY4GX6bCilazoYHfw/xK7QuHoFIvDic3VjPNaBW/sVpQ/uAMLRey3xeUNUVKkaeuVl
pH0xwmF9vcRcAjoVFEg7Mm1908a4TvMFc9vtiRP6QuNDfVQOw+x8rboVQ8OT+DU4oo5/bUoyJMjt
NJAB5KLUieMSHMNaP1tt9cT7Ajl3OFSgCp0f37dK/weJlYN5iOaZpLW77bf5BMs8+KxRT4oh8yN2
LUU/SqSAOU8iz8PWMsUmPdbddly3uZTUumbyXBSSWZD2KkVbNK8s4QqpczaNo6N9miAGxFYQhe4g
EQz4HtrDSATb/2htP9I42V1yHEgIlXBAgPT5FGR9rINYg9urKqgSIi4la15RdMglp+oH8jVWq0sO
1KF/vJ358YvM4eo0bW5VGyi8lRj5Lti44mv2JkaE/ji3tUGsyXxywtPEOMMUrK3Wbi2RX2XAO4oF
AjVtbRrHC9ATcU0ybeci6am8qkIsAcYF3M311qX5pUQOuSIxesP/ACJRVm14QrqrImDC76UEh3IY
In0nfJlvetGaIZqnXTFVl7en3Ctn0gnqmbpm5hi2WklhTBVFMAiKCb75YvALxXrsjRTOSI9tXB9H
t4pgmfw0y8vAkfZGjQJM6ejwE7I9tlSdC36T3emE5LKvD32PVJ/KhEX2GTZDs+jltg3+yKFdgiB/
R4TxSyrYVCTEPKWTtfe1aeRZTWN0Oi0b158vHJ9ZlkGyIw8joE7VjygnDmuTgPOL7ZHs+tSg5Mi1
CQS+O3ErK/Qvp4fcv3MeOzaOhvFNkXVKBRtDedeYX/XDTpRFMiFQnEAMgwRF9VrW+TkTharoXsEL
8YWP8yhzL6LBqDoKxFcwP6+kB8NHagKnXkksZhDHsehasV890wlQ/2pQgzCTtQlXmYbkUx2yyo03
EKwKIHevZYOpZXw1YYt+lwphqD00x/SUSFokRILKCrqpkOAv4tcGmvsQNAByMcxdfQI8vbvDFhXG
F7WVCTzq8+EbnfrzIn5/OF+j+jh8+HRYNhqU6fp3Pb1X1V9V0gya7Dg/aF6r/YC9lh9ChoiomRMC
ePyiQoMRWKQDZ9QsFZFYPlgLC9hKCia2wktvzE0j1zndVrPR8j7ZaCK5SfriWKwkmZNn42H/Df89
ahiVc3qY1XfQ3dfp+pFqHq0EwU80rWfs9CBMH1u32LfaetqGZU7v38bCDr1TKQWYayMGnt2TUYjX
AH/ZvAAuWRRbrjB3k8GTEFVxBN5oGxJK3JtsbbuXSrxM+afKgyvzdRT2lZ7GUvhI7IOUxPUSbCdE
logkMECXxOGNedzlt5lqygC/7is8LWmWLRY0HF0HAY+G9zwyMZErM8MAnzH8lE9hqEARrQmCqeHk
i4g+zjKanFw+toBDJfybQQiC2hBp/BoCZxI4lH8Uwpx3FvQsKiILLpe4gELREFhQVp1hxApRKsCc
4Sd4MhWTutwbGtrjZpT9mPE7Gg7YT+koC6djj5kUYozATnru2QNKQkYAmO/d4eQrBu2wG99iLJoi
9WTcGjUunIP3bf2Ng9MjKeZRKK2xuEW5TCuVIpihpnG/cGtbWIRtRkbjCIx6zDOr/zZISYS87D+p
x678J52LzebcSSVy/Dd78+8YNKZtw+W3oVS9UAC4KeAi5oMxwICCSg0SGlxTs3ylBjf7wZrZlNeG
l4dcB9Bi4TfktZ1ad/9kPKRb6e+XGbCGjYu4puSS7IcA+7la98X3T0CqLC+x2XwDMVx/vtuQLCp2
mE0/R5vQBueLq9Hq348UX+M4+10fw/+WCFeEaEO/RnlaE52MlkERIYByJpqSCckSNDBF+38do8iV
SqnkJnFRV3Gz5PFoPtojQGWhw+TlHb2H5/Kl1w7hbjwwRlGv20r+iWNH+mJeOMlum9RdEvjhO9Gi
q4W23u06EEAGrbuepGWPpP+kWeIi0E/oMoeg5Sx/TmMiosB8SCWPpFFdWz4YeHmwA+HzTxtFD/ZQ
pydu2eyfpL8gawdGq6+9wi4n9/FzBOSKugBONgi/HmKHAkakMpOVHo9KCPeYIn3tcV8sc2YB/Tc3
qhMQJacptg4ywl/pEf4GdA8/3s1cpo8dAeDzs6p0JoTENboPQCIXyaD9IoXCBg5BV5tGoKavFXpi
N6Ac9KGuC+Hb2EL4P1A83DaLEnYATHnW1npZ8h17Vu+X9UmyzLMHPstvRQoO+VJZ2YRX1KsUMQjs
nmLE7viLn0i6YWC2bBB1awut9z/j3wqhUpPpB/oIxpvOHtpXrjWTNpbaOEZ5+UK0A5thAj3dKf91
AhTDeZb4Vg4cmLsrSHX0sWqhcbFIsO1YV/nwRMkOglv6PHaAPT2k0bACrKjx/a2soqRLxHiC4CCW
kCfGFu+G4a0etMEe03JI6r4xsBs/0AhYHho602jTFRF7GOYCiUXeSCEY5TGNZ6XQ0Xp/wHEoqTUA
9zx5cQX9RSzo+i2bB5me+cnlf4YyrHMXs61vdudYPS0nRMqiuAwe0p8gxr1NN8bxrPTn5fjzU3am
qMVgSLjD2Xx0V5Y8tWa0SYWUBO5tiAv+Ktxb2WhZ+WmxwGdOlUBj17tkqwa6iY7AEZX8MUc0TFna
1rEQLm6FmNeyAanxbwlw41RrUMuwLGl5+zK6yE59OJHsAblAXNzxVWWqyN+AB/mvt6bqKu+Y8/Rl
KWr1t49D+vqsQ1kGAJc6OGKbS9mYciifQp6g2Lj4mS6LKOVS3kZ/wU6xhFn/6xL65ZQJvQQrAaP7
oqUOe7ruQxonTNQAjl88rI9zogP553+fAm6IBdRXangkkFFlkUYJnLo/MPnwjegaE8xo5YLIpo4u
HrZPe4HxwtL/Aw1EwzFVWMlqCpnXfjvJwtLLjcny6r28poLdjB3JJo7ma+6V4afdNfgzyyKJseUR
9eC9OS5olY+JchwbX9X59emNEZmW99hPlQKUjvxBoTN7TIygVQCe/kS4mlmG58Bv2YAKNTBBwV7E
4l3sHUnO3klPTLK4VouAhjSjq5fOZKBb3naN3eEzm3Ktadb4RI7m1TTJOkw/QoVLRjvMav+JxZFx
Vd9dATvdoDzxojq7Fuyz3pxwlQWJrk7C75kE3LOgXAVBRUb6hAooUT98evJNoOUMHnaOsAzF33u2
t6SwgPaiS9G7LvGh7d/I7pG/o9A9c0IPGdJ2o/e6I4s1P6xIpI+77KnKcXL8iO0p/KjSE7HtBMTx
AZtH1Dt6Rk0pe2h02FG1Mu/Pa21Bhkfnjo4PGlq/QILdIsiqDJpJVfckLdde4fixHwgxoCpEDdTq
26IIEOjz/O7/SKeXE1AjNKogn7tGDCaWsYiiw+ltMPtsH+xlYDJQUwjhxctTdTKoPOum2ToJERqZ
5QNQNWpRYduW8YDnvzdQZLQaGMmU1tzSV64WDsmt+BbPKXC40vo8G1Rms8GbPn0xmO81sLkSkemG
9Xhglzzu2lzphbVPvkg00AvPJSLV/CVG8VF0EUHl89Tw/1xKfusAAg8GTquDKuOokmVczIC2Q4f6
p1KKFpx1BizPH5wbDsI6/rAZaBsIJUV+s9LENRnhoKIeMqHaUx2zgok+KHg37FRTVyHaL8SyjmF7
PIQ8gSrSlYp2PDO9nIIuCQiCK9k/CwL1VMvDW8cKwAf8d1T0Hb85cOvivbyepEaah3jskoqDVeG4
sr83HPWH40kyGs5TBMdCr8Mn78pDArHtwqToK7oZ/6JYhyy6TVVpsuZ7qWm/PBrLP/V25jUYCzGS
6JR8RcS3vo5QSqFCVzcRIQ532fP/whri7+7oQsUbyWw4hIeqTAAjw0+Ta+w6+AWYFrpzzbcDTwis
asJKCYsxZVGM5OgDJepkD6ZMLas3yh3xLo2uR0x2FWmp1oEup57/sfHWldffIhrjXzzVrbTceODq
4P9kBt8N2InSP7w3Yj5jVex4UbCf4VuJpjOXqAiWrb1mdnnOeyszVcOdF1gwdP+aYnEB8T1VbOHZ
biSoWlCWRh2+5FLxMmpZ48qw/NGPdi4mMnb0F0GWQ8YkAdBi/5A/El+5QMcLg0lNz3zM6ExWHObY
IHSObiWO2rmgA1r/kC+jSRK6zbC2MJaVeFUTI+NEvM3EBr4fuUrDOX2tqIUFmu9ov647Iw7O6e9V
z2r4lN33+zZT+qNcL1OQctd8Zicy60Ae5EHPYpXKKMxHjGP/5bFnA/gOejLlGt8lz2siMvYvR6MP
zEjrAN2pMFTPz9mIG14E2wOZD+dJ2m8Ay6hSflx2KketCrTTpFRwt8dJKLzKtpbHE4VpukaFg4ND
jhqYnK9arXO9awNe8Je4MMWpknJbmN6XGcydcM0GG9i7j/fBojHQycCJ+50pZMyqM3qEQDjSpuy0
FsQh1Zgb1MQXckYejBL8Iu7hrm+tIEbAJjSE6MYPCXNBlkYdjKTH4QDTJprx9BjyVaaUS0mCZfrb
UwMoKlYsdmwW80nJ43dbE9WFq38ugOc/O6dNH6DljBWOTkyNCNp6X1hO3tK9m+cCWm4LDXmDbt44
+CzI11uPxaW5keSK6EffvZhmFOxzvzt/vQzLZJ4y9ExDZA1EVi8Hzd9xNx3rcqnPl2UrUQFzmvfR
Gj9enW3CrQSHUUKbrlSseOupdao2pf6wKPQePjxd3A7+qkoAth6RtZgaYSdy1PkaYYeYDcrOskZ4
iBmn8Ijn38gV7hMsTe1PUrSXRQhPuroMS28QYNxkqS+8/OVCYvkbBUz4kOMDi4Ptbbo3WUKznP/8
ovR/YAgcEb4UDN3HXmTTIi8Db7/0t08I2/pezzmWACpVhdZCFqhm+DNMnT9ZWlR8UP1VfYgahVQZ
TyuMJH34yNuCVSPp2oe+WSmsyvbRqdHr/TFga0TC6M6Ra5LK3vZ4hoLxUv7vuD7rR6QWvH74DVgd
GtKeM5elWja4yo2/FCFqKe3JuP2jgaC2XzcxsOtpGN2vb+VKFhR2kXa2fq+eHMnBEpgijX0r4wjH
67nqYIFG0H0yu8TdzGgAebm/WWeCcYKz8swTRpVZlJMmat7b7Xn20DXbyjRduT+RBk59SVhqapLH
/k8YgRZxoUb0E+Hww7I7P7TQ+NUgjoUzoK7LoWNwjb89JVRYT22zte2B3Yaa0b2m6p+QQtfQAHun
9UYYpGMAudLwGGFhZ2wlsUGvMzGOxWbm18gx4JcNXr4+748pc/2qQu4sxscUQiE9i84CnFzP8LYh
H9jveTCRgDp7E9TgApE/WSvncWS5/R23NG8Kpx1QtOWSYmbNSeK+oITlIcxCr4T74ofcZCR1jHd3
iwx2vOj7nOC2DqQ7rbN7Pgs0bhCVoMG8VOGq3P491l+10M3mGwUNbll8SR9UbBhI0b414PtlwsoR
tWllUrLHQrzsozKbB+FYz7rMtOQ/NQy5USToIMrAaCi32QyDZIAWFr74CfyjPWrikKlKjtQriRw9
3oyvrT/8FZOkkgka5iRIQK45heTHBNOMB9G37gfMAVfPFh0a9r/vwV2AXyLc0wjcP/iC4BT/G3Um
oG6WNlyeSmxLRgB76KlGOmbV2Cozpva6SeaklMySMWf0rZYN9FdxlKZDqJS1ypjVY/aTkuqCUYjq
1o7LftoEL2yx0zhpCWVcRO52JiLWqt78VYmQCpaldY1bSm+hAMOMsmcfMjNEFuiclTvlB+gthI1f
8SUJEs10/Cn8XYHeKJxvcIROXIyRbQWMi2fgvijxEyhGcONeNX1zwlN3X6cHE2209MrZ8q0/KbLb
x6eFDaXqlnxCnpkDRlPBZ3zZSjXAhhZ4lTQUJ/ZIOk5zppYGjfRMuxfzutccNXXgzpsAcLKidifO
8CSK4ckvqjQdAGXdgKIfW16hl8XVdLfpz8jdIKWtrJnp19AwNlNblaR9hlG0zNDCW42wTbOuhvf+
Ii+Cof+naQ5+w2SMMqcyf0CZk7kqXqYwqL+hmoI/XMVFFhtSMZNkuYeKG2Dlv9J6FHp+uBiFQZtn
4VTRxYscZUTkduhrR9QWh+5WzhqhEjTFP3DokvoT+hlgaAJS94t+ykolXxxNI+DDw2a6BzJNeLfi
tUNpGTujw1iHQi8h/CbK0QVGa42YGAmJyn6XdmCoWCd6xLRukzPg4N5Z4vW+Cc4NsncMmzJjfdWJ
Hu1PbMN07o0J34NKwRrtYc4IqiiAQshdKI/O0GUWJOE+b/ZbLVz4cqJHfKSl9WJpame76GaitEZf
vVKDVIItmULlGK8kgnWZsDHl4seRKW+Uhr90BjoGeTnJtCwXbd9RN6GCfzYpUMDbP7VUa4BnhDsi
VQ3/0sys6zJgL+RgsXn5Fn5LS0tInh9Tm6unh3vqnC/tgY6fTs6gVgFhVhkcNO5IloscqiFpIG/Z
s6IcMSDhpHNfFFHcP6pymEfMVRN3jPHGZrI6DyGg5ccAmAuB4goYHxjT2D5IcJVQsEYNVmNsXFFc
3Z8S+4HV8KFwnDlogeHV5Dqi/Bb5VY1AJY5vZ6K2PbV6gV6J4PLyQyhe4NGPzrtb5Vx0WqhJm5pv
iNWGDVTwPE+h8S3UrMlX5zRkFaBihaHUX4ssByz9ABsvxIoVmAfmCLBZKEuXFsolE9u/ubq3X9W2
FbHcrp47BB4Y8W4kAbswH8upXcxjKk6jEIJrJbPxih4CK3YYttedakmx4CSXlqgE/WELhEKKW0Ym
gaBC9xF4RXtDZx0zIQZxTx08QJHcReqDENLR8hs8Vw42831/23F4VIY2gfivLdjSWZwZ2PoQExWG
cZjB66Y013XEkpYZssEa8rY+cCSZF+iuj5shUtYEb86YAduKvHaidbg9IsJQB6Pa7LDs01auTkRO
2MI8r+EuL0DbLdjoAW8xSe8WKUpvNH0dP+ckZGXQw1p69asgQTFq/QoKJu147V8Ld3VhfBHtZnf7
aPXmY0IBseut0unIZzAaD1Pv0hXwKUfZ9Gqtc7hqJdJyAOSlk/tlx93fEeN7XzFRHItbdnHRqXBe
qXs4QvmwXM46TZw/Db8Wj2CsEXGo12A4bnQ6XjtPA/B/4TAgJthkckb54F0cFjy5Wsjf1a2lp+ND
MxGpN0kMSonqhdn/lwV9NzHnoxAaVzPduGSEPH/UlSfJVyN6/PnUH5FXT12+f70P1SrADJjoau/N
qvX8pIUTGQJ6GV2HAT4aWmALZLPs2rOs+J1bWU/WD/jvmHE5blTk5kxq4Y4z0Uo6P8Z5TNOYcnRy
hNONfqPbCdx+Gp9oRhkz1mZMVkjoVcF4itK1HlP6s/pOrgnxf5LrKHvSb48X1iTm95jDQZCxrWRk
6fvJ0owJ26DQbu+Dzx81mDXe5kt2iS5kzXHUUI9r0qZ3e81P9yBGDy7EifiEr85YwsnZnzoftG8P
i+xnmCg4w8h6EWaZ8nVHPAs7I8y2iMp4fx5UC4k+8tltPVWOdVD6ekPHcfyMUuQsiBMNo7S5/X7g
ZbLTrv8HprxlpD6ZvuO3cJIOp+HIEw9nBREVA8jCAHmBvP1xG4nqGY7Iwt3uRaef1aBcaDeG24s8
7/DEIBJxcCcJYorGLEtQ7CXpzFvLrybweuAL8zF1i33wH4DJf1rolK558ws9Wod2mYjDSeLPXncu
iL1g7wcOaDW1xLBipWXkmm+nlKqvTPsPFpGmrhmQmylij0wMGfCOkrikq7IYiCR9uEcQIqJZ64vF
leh76+QkNRrUImyNhA4fJtMxnawBVzwe5Yk191ABe90MAnB4MkXgBmAiBVa/I09pC0/5yTHXy9Z8
YBZ6rs9w54BwYLfAx5mEAxMsMW78kmGIDRpPcKKgSx5McNZ+jaGtUT3eSO7X1tpXYI1RgFVHkkC1
IOLWKD5XsTpVdlqRTjzFm2Nu84M6DUu/tFs5uFWK2JWPwEmcoplDLKhZWClMK5S/NZ09qsI8NQCj
Sw4N13swXNgvidpNt3ugHHEQGnOWG3yj6fb1+8SXfcNtLjcXC0Bc+gdiZ7OsD0k0Qt/ViOqed9zc
NbwRNEe/o8rYJIuuSEF3KEClp1DdfpxqJZelit+eM5MlHGd4BUW0lJkTDjsrFX+Kx6sg8Q+1qo4a
HD/GbqdOioGpRW+r1slZxiFL4LhrE/eiiBvJKh4kvDLDqp1WzaImQAsTQHlKbjbxUPBVi4AO+VoR
SRQoypJP0HQFYLfAsInvgqAoYcWHyK8BQjC8x57bKjvBWqx6z9JRDJIpGWqyxauP017nWtHWVdYm
kC3ltDWoGqzvI9U89yQFeypF/KK6MfOrfAzmElrf6AlGM01/08rdTl9e8BdJf+DbqVFpIMqTjyFz
gvR5z0LhGdegyeb+QV3UqB7xCb8jCYBTg4STyAT/CB834h3W7OML7gwLW/3l/nG3SOSRTPwKD4Tj
UlyqUZ3/bDG10KPr1FnncTfag2BpwGhGMYF+uCdd0eiF4rwMXq7+3ekPUxg3R8NpMkvSDXL0hkHP
nVjPf7ZwwnDWcd5wS/1XjYJHv63bglxqGRZc5Q2Ahv9QxLfrzRp3XyCcMLzOr7Wi1oKUEYgagVgy
jA2QWCjoBS/AgbVU/GQXQsryR9oF7+usNgpq9k/2clcJD/kok4+e9x1DUClwF5kKhLhvafIgtoXl
owwEFVatXFH2xKq4j5cs5rcADSNUP3OjvyxqiiJ+7ebN76QmVJOqv0dUH15spj7seYEcS43jgyDT
rAh1sj1efP6FB1OzTxg0EGjjwgvdnDFTobHlya9p1r3TqrGmzWbVKb6tWw53lG6VoSyj/bqjXG38
wZLL9JpnFqMfHPdt/LN8WOym7Pn7rlrQgmbxci9pEtz6E56/ltcqhkCdRXUh6/7+iWJWkUgl50kG
4rTlwskHquiVDE557JwPuShCmCSP2lHTLM5m3j7uNhdHNcYOcWCmJNOeMU8cyrQlvXXDDHsNThwP
96iso1X6S5VSvlKA0OLZHyZ9nDRJyjiy57VncsKPUCLx51t3nb93sJBOL/zwl3MlHg8Sym1X8RCu
jTI6jQbTWSneVD+95pwkKSi52j+QTmtC5BdrhCci7QVEyqgEPTs8wliIkmJ9HgIvQZZllomD8Cev
UjENcEZLvZrxFAmycHSzYyLpvVvOi0y9ecRMvZzhkWnOD3UMSyyj/Cq0jGXDLUab6yeC3ArGagZZ
HRZaAcNlzFXtZWaHMJkG8icPmpMDv2xgZ8Or+95lqKyDAlTBqbtam7W0VXyI49hY0fhcS/qJOEgX
ym6kdIe9M4Z/O20nBV4+jJPXe9sn9wjYVdswlBDXr+1sjRxWWy/vXWeRY3/XjlSbOK6yqr//dde/
+BA7rz3AaNc8+NgaOBLygrS7QME4CBuKMfJ7rxsa75hnRcZ/n+hNib/iVUXq02V9wWqyGq7uS51t
2NJkZyKXTzpE23+VJ75vc4Uo+NzsoPm1r2GxR7AY+g487OEh9qZhtDUNIbV5/Ct22VW7+8c2u35x
weNomW9mmC4vpUjMCcmSq7/Kggq9e1KTeW6r0RSAg10kpTFFPd3gyyDANJvq5f5OLobEflEBOrA3
jVmBFbAnjvkc314vMA8mCvvwouHPFP40O4HBC3hd/zRGczW3xQ379AA6zm/7jh4BgIakWh+s2yhe
uJVuIh8p3r6blsupIi8U0DMET25B2ZT1XEVlTz8gJBIkQ+1F1YeSSwIgyF/mluYP54T6n4/VX2l3
iXjzoeqLnGX2RfzXSP1y71O6aMvIjhhvxtxD2Xl28WcXDM0lOqcvI3oQCh9LNkz/Aqtz3ohzU0tP
sHK4N9tR64acAG//mpUK3oyQoXtWb6z6M9JgpJcl2ihoWCYwKK01NfDZjAt1qDaNPuxPHG1ewxqt
M3vRmcXsagBHeqmUzKjfFNTp+gaj8E5cMyR8LroWwJf7csRSvS5iLYr/5heC1daOg2b+iOmbq5MF
hbG9Qtz52NLqXOtlcvbPyi9QEsjqlGFMMMaB2xO7t29oS6cF/JR5rUAEyFPhQyrfvcUEJLorqRnO
GWGBMGn14YUhv0CZMLSpp+3qUHaOX+5GtmT7qUaAvieYuiboZjgEV3opgFtLlT1etKQI4z63OIjf
ReyGVyIqH/RzGTgT4PUEe6mjrRfZASbjtcpSb/iudUEnSU+iwkE89g8nhPbMUSqWeZ95CRxj3ipW
8YNeUPD3euYTj0RG0R4k2f7AtidxqoXGdCv8gQFQTO6EbahE6D/sugIUuXdYDMsHdiC3XOEIeuI0
bc1ehgqYD0RAKo8wUWpHHgzqKv0iAsui6T907UF2L4TW9pUiIT42rIuDYtjb7so8NFhmIe/6uM3K
UW6HxTO9pg7i5ZiQvJe1jDDlS3dV4Kha+BFXiiMQ4QkZfSYZPCVP9u2gQKkYyd3UYzhL5++/TMnD
msTxDm2ZSYQnWbpyNHyVuIokbql3Jc5OPEhyxLwIeAWAOFl3SHeLurwKuUi5hcQ5vXrhaERPNiBo
GK8tpje3ocabEWWfzs+mpuwhQxLbd0AxZrm9DSDH7uQjpvVZIk9Dlx4vdC30JxfrXopDqVvetAIQ
Bqr9s87qTUTPrCCPb9enNjeULtRICcgWZL1mzphbmd6rwHLIDyLm2AjjuSzip3TdjQg3sPG+TOJi
5uLadc4eK0wEJJsfCOnmR6YrTddiE4miRIQdA812v6i2dNLhcCwanmw+96HAzEuPVh0a8FvgA+rJ
LVe5776pSpXconMqrl90RI2PEV9rBaMO4CA9NBXkbhRqYvvlNJ8c/YxFcBVB+wL/yGD7tyQLede/
nE0S+rnPnOrM4lTiT9X6UusrMqfGyML/F6p5C1XNGBIFyn6Gbf6JzMzT7+wlhqE+B6OTGhnhQXME
jbFmzSH0V0HIdJVMGJGkVSCDII/tCG6YMm/e5AjdeYMzbFLf54pdGm1U05p3q8qutO/Eq3kWd3DJ
oiMMIPt5T9o9xaXYFlAT6DoUCWGjCcaeFQW4GwXNjVdlf3QttbHjal04p5Wr5pSBA0vAGWBgLMf3
hVSpMC0mE2JHg5JV/h48bJ2xwo3oIqrYyIIN9zQzBowkZ+kkC5ulws1JajqOMmJoIv1lVcbL7lcG
YGcMM/9c7EkUkOJUCWk/OcC3eq0hJG86vOMW6y2EOFACL43AjRHF8dNGSF8/v1xV5LTzmxPeqHLX
u9d9Zrj3jHDaRedQWEm13Wo5vbmFH8/ILqfilbtLV7fG3M+M1X98943hUzjyiMMcpIkbD+YciqCy
dIcySxNhJdqpcicW1cUzvsEzKoKAObdTqBMnnbJ/iyC1iloj6bxLqE6EP5IDbh18kHZwPVOcUAhz
XsOvGQp7MB42WYFpiuaLzj4YOMLq2EiKd1/vhwjkNsYqhIYrqkhqS/P9ZNAUoLB1ysG05Ec1reuG
kP25ywYEN36h9NAWRYG3b9toozbvl2W7OvWLGifCQ6lODebGdqdJ7iB+Ml+a8qDpErJqxxnfAg+S
N/nnCf7t6Vzg83Aph1iX2lV2lwbUbzXiJG1V9K+ceJALwW8TLIILPgU9GCYX5A5JvSk32VgPm6aH
tSXEGY2yoJw54UTg9+bzq6gv/P/2Rs3fLtPHRlBLGKeyvt6Mbbi7ZzxH+eUxLK+vrYnOl8rFWs3V
z0xeJhR1nUVJmRHlwkBUTho7hTIOGuXnpS8go1B/tchmNwXlqkjJtAgQP9M3wzE/5cJxuOukubEg
fJRd19AGkwZTST7H07TnytoH7obmORT26yH5P6+ysi/BUTXK0xwZz2A76eX+fnKgZCe+z0cp5w6w
ML0UinmhdFAj08lfz3axrPKmf8Pjsy9lf4hO1vuDZt+m2Ya4xnqUsaw23eBg9gDkuK4l4SkgNZF7
4UQq/MPYCzp9LEbJtAJPorqnu5bhupXwch45VCvwsuh2Qjp4SOUqdQtv9vUHPZTDjIlnKmL5mUFC
hqXPfpGDPuxTZZN/3Fu6Sfshqgr1BY65N9xLI5tLK8k1GXwrQF0H0Co70CbX9tffVBBjmKRzvEBg
Qd/fGADfLT9rEzNCkI/k8XOtNpV7N8t1TJdptO5gNOihq3ohS1QU1TgIyvAuutAjJrIECmUStPtA
OEDgdG5+5D21WVOz+kE2lhoJ7ujPNnnEZk1hMMuTNqJ6+spwU6H7e1BpUzro+eA/2cHXM81ZoaWX
B8HlC5sQicy5YHLW+s+DTgdLiUsTKhrikFzm+Ug+zkNeDjsNHQkCdppJ4F5Lz8ArmAZDhBGOcNQ6
TeseeUv5EgmpKbsRalxWsjoe8avdz5nMH3nIqBFvqsJEGdaBvtugewnPGmo3YOPkawRxq2LGbX5t
bNWu36qywNWV/ksnIuH2tKn9xvTF7asTF3r2IZRY8tiZWhwgZ1L/8dN17a8ODwRRNBoG3NsanwFR
PSVBnC4cQvvbyrBQBu0OTcVj3tzHWwTy2HlTM+APIg+y4osOjy4zgU0olp2Gx88BTO3Xyee7vy07
LqnATsOEvuLGowj6IzEZAynp+eYrpOCMhjF124wUyyv2wgp00iA/75FSntliBe1UoR+VY+ko4eV+
zIMbdy7m8Ep6FRxx4jozAKnlojlS8IEu6SX1GHzs7uxhZ4ZNQ8pUwlNjjrW7q6K9r7XgFwOFYI68
6BywuVG0r9UZCLw4d3zpmDC5p6mOtEpFi0G6r/M9IKzQKojIPgFmGWaPB+vNTPgAeXQG43Eg65NN
fkMYxA7mkZON6AHlcfod4LoaDodYygjeH0D+Mm4o+TYr50PExRqBBN/OwmYYwHT34G57qQLKrJw/
Nm6zaXPTs3mgma9Vex5PfE2CjAyRiOx3wUCNmFbyWZHjr9QbhgPjZjBmqy3+Fk11nEHEX9qBAN4b
N0t/maWsoCO7dyCuwYSCZDXI664Bh4YPPAgUmH8Q/SCAA9zfl0sQURgxuQ8nw8qjde4FUUURMc8z
UgOgfg/Wf0W1g+qyHkpce6gigI4PgaIlj119I/agHZanifm6GSIeuYyQB+L4zrHzcLJ7n5r3hlDf
lOdePp7NzWe+DihgvRL2iIH78nknSyuKm1CtsLlRMWqPLJJn0o9UsjSi950Pczzy3wzCHsGOCZ22
RsnjFGPecTCrgf9AxDf4cURyjnuf0Qhkjlu2jJeBg726Iz2cOjYZ7yXMC21A1icMdrFLVEbJMPMQ
XdgSdbXZyhGTH2VpcNDAvVVkXcHiozxl/n94X3bPDqvlYaIlcKgbK2PajNUlAtlJR2qEcWeiYAMw
T98bOHGsUnWfJOal1ZB9A8OsQj33XM2Nca//QT25DvTAUp2VcPyxJEvLXEcf0D37MRAYWPM48y/7
kARZa/k6UaUKmrRnZCGDYoNmk51FBcPO/+dEpFPQ6C9DPg5cNunBkpJsv4DdgUeb+GHbdK9Lip0h
YSk/U4Cvs95p7bDEX8wSRObg6/SwbCphOytcL0z0CMe4hmOFUASH0hFeOikroWxMX/aIcH8AGOiX
qRJ/RrlubvC8QPbhuAvsffOMIZ/c3MLlDA/XzpWrcX0lybebP3Ju15PmnDu/Yqa2ECHaVYnkIiwD
qJ9qrOi/4SnZq35rXsy8j/3w9TMgZvN26SQtuf8ZagdlHBuvZYeX2Ugo6NkqlRNehoRobQUixEiU
ar9nuGWdcwwS+1Plqu9TZaNK53s2komC3z0a7qoaCRC4PuiISyDiXPN0r0aTd4JAY55AKouVSG4M
mKzZiXcZE82HtsGO49+jJuqFKapMCI2CxUJZpS2S80bLw/tJfOcvtId4ilURUNudp/zXZfeDVoNl
DCp6no/TDilp+ZaVAD2oX1+3q5ZfaWPt/Me5M/tpoX8trclHsQ4FkKzEcHxknNss/VRGjcUYl2rX
AbQn5l11Wz54KZaqkSmfEYqn6gPkyHosMgbTKoNWk0rjxLJWkN6xIlAaBRSev9kah4DbVqeqGBX+
nB76/pAmxgld0QRv/5E3n934tK/JITZpxUl9heKyYxflo8O9/ZFOMfgiRPUAhru+Dea2HjvmEXSE
6cL8kCLdj+q9hypZILTb76blqOC50KM3dfdI/canQWOEd7kvb+O4eVvcIuP4Cv3CnNVhCkyCFFhX
mpOi968URMCvLjLWbqO5jc15zjk1EtvSc/9G4DqPkfGhLwMeP8uJv0A1eiHxAwRcEzzawyHB3oIa
GJNdA8Llt6oAjuM2WLJCtcL5elfZsecs/EWdbXysln6NVuZpQS9dvz6s+g4Nu6MCESQG3qM6nirk
PL6l61LShv8SWE5geWsz9glbfoa7lZ6JtdGAhLvn3cVuxTr6ir8Pvbc47/EcSIe7MpP2HpfeJrT8
B1xanYkucLpvSkqVMN03uxJ9rc0jsGAHL4mMMeyPCbxzjcfzrw70h5Z4aJ85b2Sw2r9aoW1yJ3/5
Ep2IfxWdYekiF2dpvrLxrwf26DHJyI7Ww8IRw+6w+aLKSJWAKMZvyeOBQ5E0+1AOFS7D5mNWEd7G
yCkNgyYtW+UaA0nUIlHm0nXFao2JZSuIIutSjt4O1naP7rTPFj4mz4K3UHbaXxyTlJWpW7hehsII
DMf9jCruINeBELJjkJ/YAVmDlUmd0DQMWD2HqkQSi2aFF+qDG3wWS1E39/1aT+y5UaFZQZX1TwfL
HIOaNR/s2DQ043m4KHjLeRfsys90GKa/yHQ9P2zRKJ8k5i93BNXpX1DNkeJ2WU/otc7/3ElP1VGr
kMi69a4ddsRbkM9F8GLFOpx/IkUXYPIY6CIEVxkzCZHFHmEmeFKXOCqPZV/Hbwg5bHQYzkTBv5Gj
XFOxCeL0vStqxveioat+cSWHX3bV5nlUjIxNzsLpJTVWHsRxIgAjqGM6H6kG4Nya5R0cmnxTqQPS
0X1gDyrGH1rP3sqQ9ABTu10pBS1iY0FTRm97EkltGSMO951zjH4lxloRxsJG7D5p1fwLnUJZweVR
sbljvSNVIG33qM5SCDKtVu//hGUOvdkCDpD1Zh9SuTJ8nL+cmKUocFvCvv69eD1GNXjA2W1NBEWk
4ZyxbUQP85zK805OP/53TOLEV0DrIMtx3TVXentt5rcilI7vRz1NmYNjyJhSB7jq9zNmTnD3gqYV
WXZusfe+ywB+Fm8bzQOrIKc2+HXwPEfGJkkHnMNp2PNCGNpcrCJiYLvQ+rvtoH4DOzIneDwM6d+P
CS9ZL4bbPprkVYi2Ywj0Cx1m5exVg86+T45blowg5O2i6r8wJvmqBDuCRA1C26oo6vJCCF+wWshM
BkW/29z1d87extIZECRLEtmZud3KHCB3i1+QHI5Mks4y8qn+kNr2uUbxp+ljA1lAvHmZVnKbDE1C
Hj2R+GuY0X29DWk75v22TGlK3qZ+pLIy8g/0B2IjGHpXHZVgdLC6hRofeK8zcB2ckg6eXm+KV1fi
nMI/I3iOluzZp0NmL8CWgliGDZDSJYOD6I6JL1QeUKdCVjfb2A6V8AitzHQppHX1PWyJ65XSUqjU
cN7WvldriagUOugmAoyLq2yCPct01EUp7XMa+qgW/i9zPJtuB59/WXmNAOjpPwUZ0q1GIK9O8Q1P
xsM7WbDWpiGSzRaAZTtd0KtGX9jn5YCQjI3cmIkyMq4Q++MdQrJZj4Cl+g0ddPayOBOy2zPrhF4B
lKrRz5YBHBdyaiaOGD7DJMxEVX0SaQP6hf+EbkEP3/F9FnNwtmAI8dWUsjm+PNfCQe264adsabyF
SJ6C2r4mR3QvSunxaTLXpLoQeDZBRcSb1mBk2jvODdUz6SiomHF1mYlHy5lx6OSUy+qWJeD/0uCd
Cpuo2eveaYIQg3/Rg9j4gljF7QN/CGXTOqy0OF+Hu4sfiF5oiVA/Prijk01WWEyi13Co5xXcoZFC
snXQRgCPtm8Rkk+uapo1EWswM25deV0ahx5ybDeIUczZ+JaRsQ5sBvA1mO/swueIoQD5MYhVMuPy
2QzwTPd2gsYNIa/Fw0wqSX5rdPeQWnrcc24zY9ENCjvX4nDi41cUc928QAoMgd2DaNhAHUP3yZsJ
CsijBF7lSaKsm5Q1s1FRa61/WXNeXmlKrIdp6V1+b/YrtKdT6gMsFV+PB1BrtepIkPpNBwoaynZF
0g228pVaO6y3ag8eWXOldqbRXUw1ImtF8kCTyrGDmq31RV9rSpRLl3+TrPzoNGcAubbLQKeAcUCe
/+JHxBBg1rSI/EVehmCQp/RnKhUsSNd69sONHtEvLbDlmP8sWNgx5MxzWVx6DUA/rXeMi8Nm06Nr
VbRaqhTJo3y7J1E33R0mvCE2OP+fMHCpDOLyDmZic8YFWqShFdN5NDNslGgICX7pT2yarKXNwkkA
zdr+FzLvHHqe9c2fvdHoDdegh8yQEnWRXaspVUO6MbgQdpXxee/pDmv58+XBpZIXbX2aXo73FhpJ
ViUv08reHIVZdW2FS+zACE/0V7nC7h1pro8TzEvVzL1mWlg0YUA+4T0xRiMEcdQWdgU2TfugEsvO
ok0xHF7tKZh/IGitEY8ZFI+RdgueB8tSnGWL7dDxK0umgNV0AdSe9ekX845p/6y9tfjLPqLJf9Zn
RK1vdTk+EpWNaeSzP7YEA7CKg0tmVUtss+bgZ8VV8J2bzy4Mn4yAVyE8APOxkr8DCuh5SFkgm+Jv
/l9cZXzEITTVio4EONws1Sq7IxzdM5HrURCwHp9/qh3QWiRZwAuMpw0Tj/q76qWOqOxnk6rdszLh
FF3igFZUaHjxcASpCDNAjjlPrtT78rnA0JBnpuTUwrtX6TmHhvd11B2rBX2YoXm4HwsQjcCbsCTm
nsD4eReQYp7yyqclxg6/MzEbuksrBdppaApavmTVnQjZuyK0oMPg+cdZVDmUpiiYoJk2oW9sTp02
IV3S+mxsEmk3CHcxsEJCN4dM8H733SlWqIfIB/KwgolJbm6ajRCuiGqfwlPPUwfJaB2VALK3TuNm
tkpA5qCY70mc5KZjOMgBIXC3jhWZPsCX62mjVE6tgKvVvQVgevPV2tXBcdOEX20/eQpiwht0GWAT
Kw4tqZgt7jM+I66KJDL1Ovn9SK1c8+XmBF8PwXJymmO9dq7UY0VVsk2fdoApWYn7sJkolPFHUkpj
IXYihKUOLthQU5dUSHKkK2Fm12FswFZfQNA39mixvczMekSRIt1r2RzVopfg9pkrnqeDYx7ljj9y
IrgrUbKF1zBPQpc/Aur61I/s8JBBWH22+xWt4MMVy9lecw8n0DAjcuborm7dgH7NHe6sMmx7em25
FUivc3aI244oeRiZjfmbLYmH1zw0Nbt5U70TK+FqBDqJZ/WlPjjmNHXpvkEgh/pi/QkFgQhYMqwS
+fVS/kQnRG62aZ2HON4beVydo53/QjcCTXcPVNaXa+rL3RblTqg+xciCIeBTRyS4qP0c4OV+q5A6
sdW36i92BGPmnnVwiR7zPKihOxRE//2fzwGzsc070QZgunYYZs8wbLvv5iC6oWS8HiMuarfM284w
sxjb0itsQ+9piepHsSYT8ATqRIrT6IuJmrv8QUSDGbTZr62QiAk+THo+aXAIVm9ZswFbKz8tcAEO
9uWILslG/Hj2a9jbaWapOPnTMAisJvtCZhpQrrhjDhMeZljBrh74McPT8wtR3OToRs9sDQClRDkQ
evzuXZfCvT9895on0qfa8MC0Kysz3V0JDiCXCLF92Ab95aCyBJe/S2SVwlmItXbQSnpAbK35EI/R
AVEx6uFbPX+byv07yYlkdJmQHdgUog8UQvds28LHeeThW/G8jz9+VyTwm+D3BXjnaMngSEXYQE9c
1qA92YfbedJ4TpyoFc5RzKQ7BscTu1YR99uKZT95cqkX9LY6ICulKYQWN2vnPOlLWqlOCaleg2wO
0hVB6tQsIctKYYwvg24w5JChgFNPQ4MrRwTjWvoouHpyQ+GsEdk4xdrq2x/vAy3VuBiE3u3znnbe
RRJYv2KmN57ZU9Fc++LmzyeGCe6fFhkA1cXWzWL8tZ6yBba9W5IYiBtJOggvj+CCNt20D0oAl2ZG
8uyK3V6D0lfGKUpyIz7Zo3MMM5T7c1MzAKqc0Hg+LcejSpml/7Wf4MH1UIdqwufmiM3h3KS9zJog
KNJ69lQrWLhEj1YUI4LoJ0znS4GX5t9YiQEewgzATf+E586ui91y7r7/63lYo3c5jnOa+IEQGbD5
YDndmYTB/uEbv6296LwcbB/VfKfPCN49cwzRzhrdPBVCvenj74P3TMt9lwPxXk2yPNIfgSjUbxlF
BZw/GYDppNIJAngn2TTsGkFKE9ISzvYvHSloXFMh+YoXjehrsptYoGpGFGRHHU65zuGDYm7eX6Pn
HjPzgXWViY/vdgLofEVeR8NekYzK0at7NwkbYYxuoq25z7zg6Dadmn9a0U29gcFso7ZoejxaJhwI
t5FJw3l9FaNsCo8QgAFu8c1SUreyWcecR0bR6KEDonMLASanp1Sv9VdRqiUUxV3da/NY38UARDU+
jC4mUFNhtigh+VESYerWl47Yj+0YHso+/JjO4gRqcxi0Mv0DOgC9kpABXdKB1J5Cq1AfsKNd9bOl
BkQTNRL7EduN25UrppqrO/fv7qX+DRVT+By9ekMDZmHLAdlaYO4kaPGZjmduct0U2ud7LWntvvJd
+ebl7yAT33F4w7HZoOpGkXUZcVBfAs7MEu0LFE+5/2XbtrYIL+OKGHvq9MEUCpsYvEr/dw5F+rDK
MRfUTcVhbpE+7ZbHkGJgAv2hdOQkYuY8iKnuPQC1cMMGtMzY8qd0GUquA4v3+eK/DWLxZjuHwnfc
felnjx2YQcm8DvhdZMBElQNffdPpOuEBWsOpHdzgrTPOOxvoty5zRh/n99SBcSoH44T8da2XQvVg
/7O9xVbkR4dfOeEmlur4O49qAhShhmZ0XNSCTwcKdWeWK19exsp1RU0WvUxc84KtM91v36QxvGEo
OJJUbFmjvEIeNo8SgbkwHLguCD3lgcZDOiBoHcHydcLNDyZ48QDbDVqF9+6KRpSawsO5rahoU+cg
JiRNT2iCrpjNloyHPJDKp59MbjEu3uwOHc09HJ546OLCRmilrJYxNFh/xdTjZv0pZRPNmkyudFG7
KkgEweQr1K7EAeSvioShM2DTrqjHZ15jnrKbTva9ZKwo0iB2A/eMeTOxeEnzi7Mcaw9IeIIArMZ8
GDHbEHIuKc7orljwdQuCaBSpYQZ9GiKnWF6SxX5YIISHDgSzLx7vIlTSemPOT9kX9pfR/8D/yPuX
HXbS1y2pW/uEWyxaFdMpKOsUjHj61slGkPM9arBDYQXvxh29R6tUZgVwuN37gnMc99gqJ8Ik8Adj
rkfmvZh8gdFvdhMvbS3UXTcLgCiN7FJWP+DRzTmXq1W9sibhROhE54Y1hxUEUpz7JLwXSLR7/e+g
M6QcObqrOy1nfXRlTfYMWCYnKdLM4r+5KjWz1NaBqrchUonO0eYKBhfpdsV8QhPAbieijdNcn3wR
AeX7quK1KdjKBifwHm1uvAW/4nqa8OHT49x3TjYrONijuh7KKvnuDT2Xf2slAfMM8ZYFhXojAAGC
zd6wWAMLUjY+fw1TlYxq1NF/W5buw1Fuavg3hlErgCKTAVHhjK2dnBTy1FfkhvZpdJ+57adBdD5c
lsWw2mzvC5uR0fNfD1WitaxFvC+PO0gABB7EoPN5gcJkO6sBrW6Lmz50lGPfvA9T5M53ABMf0AOm
wQe4Yg2LTnVNz3ns9cOvvmUeW0TV1/kEBm89mxTTivQeBMOsnCPqd3IFJkPxb+gFs9HuPqLy3Kh3
u0ckfsRNjVSLJb2xy3dVtBhRWGUrycTEjQMWEgdU1e/SRwNqlLG74tlHnaZHYGSTclqBYvWBaY9l
YkzcukSKiLTK+CvK+oYPU5FZnC1+RokM2oJOuQja5WmFItZzExZfdqq39QPmmIQ3vWKIno7SLI4q
FAoab3o7IlWt+zGgbP+9xHRa1BnzBlX+oni9qBhFY7Gm3THdA8i+7EtdeU12mwBNVU2sgRMkuFtm
XP8k4vJNO6JLWT/h04iGVqmgRUVEjxttV6iAqcGTGf7tUO9X3X723cG7q5f8yNIVzDh9Drhho7aB
FbRmKm8cbsHhC1BP73Oyy6Ib2acjkfwPG0Sl4OhRPQhdBUIEUbVBTa6R9YauXL4gBCrh5bC6+z8z
8xl7IMj7LOuAG8A6cpOeuIwuJhnz7KO5aUJ8YQa+o8RFbk5ckpy3vuVNuEnr+/vNHHwy3jtlUrZV
l/xpUHaoDtWDEiq8RVPbVOgVmLySx4gbalzLj1va8gfgGZBjc0Uqev/eLFdFApIi06HFXo43vjQx
PDFKaxRK42YMCgzA+hYG2r9arvo83/8Ej2nmsZar1UQGpOUqnKOLHcuaMX94hsDQ11z2ds+R+qR5
QspB1+8PlRcZSaJiyuKk3egAw/Npq5/03rPga4Zdx7XZuSQ//f+WQ4JpBvQZi+bSTXBS8KJHMWdi
DPFLEn96LYFhBvYqA5+rC3vs8fglPsCvYSLV6Jy77mDND+EktyA1vRcDhSfDwWMtr6knBiF/rek5
cRGYVK2+Fo5LirfgDXQG++dGJ3wwZNYY6xxIZtUFRMljEdr8zj2qaOQ3dC9OcGtKR1je6eQ0fgQn
HsI0Rr7R1yVglHFbgGlDaQB/FiE7ltWbOx5L74Utb0CCDreEJo3L07AQsJ6pU28xbvRrpc4Ceoiv
XUmFgjlfOfweQ8lkwRtjuBxPV7GBdqvOOfY3eMFOMKQwyCyLmnoxvjtjx/rTxGEsY1sauU2EfZrc
+GX3OetG3qc1R7eA1RkzG5pHDxFZQIsoPkADspR9SMmHS2Ag92OxPF8+Y1bqW9avIzrbUFARVyTm
eanPvMQ8DyK3UWgZ3QEfJT2FaMtM1L6mKvritjzaleCdwullZ7FOrumqNqxpXcrpM99Sj6QzEwA/
DYurr/mLpuhT3ln+fcASHVZca/rYhGVMpCdWnHFYQmbGzrX367EP0C0bFiByklGTInJtTV5EXGbW
chjn38+YX+2N2XzsqEOoODFHz8+0PEmjqSBCjlpoRGkere4PXqd534U0rItIcx+eXn4qlSPGcqpU
rhe57A6uTNxXlKzrIRwtLr3O0zkaIdGQvh0elCmUJ9pf9RzVhryyiJhB+/pfEEJLC3o9hJsxldnS
lDQxm3Nuu+8DkHdmeaswyOiokV4x7lHJ/SsmKxanQ0WJRp2Wkd9gIfAFyLgirBGZE9EvTPomk29P
se0wSNYFRe82515SScclmBUrvT49tCrW0JZYWroX0F7oUOwUnDlxSnx+4SkEjoEvY05iF1J/jm5d
ymhumnFIMAZwWkyzWRorQS1JL9WYalAlW/0ZOxExKsIoVMvsNMvpmjuRG0uduMSZE0vMYeyszhNX
c9EhUblS36CtX96ZqliZaDMUXgyX9S71SNY9Xpig8/LmZ245P6vQYdW08qRbcMxjERLg5CnuKGlq
VlY6LPrGwoTdtU7eMackgfwWN98AI7mc/x+dDvhPobyWGI6IT37YVjCFw6l6hV99xvmAwzqn1D8f
Hdw9Y7+iEGmOVlv2ceafOrHNsw1BFP6GJmC+0HhncY7tdR4X0oEK2faS6/jQWvcxDz/G6SkSek8z
9NAlmZADuZdvs74XvpFkV93A3v2L/9v6CYhZs+kYqLD4UNT5DzjneAP9Y+cfEENrQ2AX/Gdd062L
QKAL3ruwVF7KNhLyYTOob/aLs/UdufB4NG7Nca5T7cNVPca0CwXiRaQ7Q5Sgf3kXPxJ7ox95rbt7
aX4YlWYYJAtO1jJUKzFMvW41To+YS5PeKsnHvAEtE9zbd+qzZ+B7Lt5IkIimNohDZDwTWP5y8O/t
Z/NvHIzvGGFTBMW/rKPSvQfln2S0rPLnMkTkPY5TwHgGfja1wJ8ag2fpuw4DpYOvYT9kGMYYIQ3u
IZr/fR6UEOn5JmA0ZhrFOOt+Q66MfDksn1JXpct2o7ALsSFKAzDR8NcTe79LZj/EGDtIZEK+QnPN
9v44dzgq+oU7EQ1jyCXPTL6tdF1VONNuT8VUqg11U1Oe/jq+rngylC3LNnenR/xEf2Fr8C0N0tRW
gIlGBpo2UdBc7ox9f/pDRleN/lWVupMSPmjDEpA5vequ+cTPB4nfEPg3W5YF3lWSaLv5R9BDGyG0
Vkd2ZHS8RmaZ9/Atp9Z/zVI7fCo7RBcLeZjQkuAyZ9DOG0SwwEnLFqtZDz3oDyx6RKfBK+0EhKzw
FjoQJdMdSdWj7tvfsbdIFj83A+XmXbqt0Kad/qeXAyglypRoZIxlU3Rd0UhEZ4fg87CnFlizN+Ik
sAoKBWPhq+LTYNxJ0Ouu5IjLfzlM546XL0iyDfgZSDxDR2SLec7cBvj/bE5APHvxqjXLJdRJB6V1
hC+sGtksWYMJHTJGYPV2ycEKySCOp5+DAwnKzwmdEueuDvLQ6ZX67kTTPdTKzhON5XKgZ5M4hRLT
QLTubPbwreAq6A4WyIUdlDB5xWQPQLrUn8WyDHrv/uJUWkL8oCATSwqM13G8nJE6Ky6zLoUvijmH
Ri2MmBC3WZxkyNvnlfd74UbUwQvm35A+Kny4T8GGAag42bYRrXfvvlYeTV/e0+8nePBpF5LcfiE1
cZa4ajOTv464huYbNigT2jGlgwZeWtDnZDaa9cfsgcR6+WP5NQgRKzsSGWxLEUjFn7QmLEyybKfH
qwxTZ0cBdf8plXBt0KxEEts/ZZv4IID7ZL9LHIOi0FsM+SFsQQGL7VowLvJeNvrnb1LluaSpP5Mz
CneNBaPmogTKCN0c5SFO2RVc+dUBHiRO42lvrBoBPGuyl9RvVtSpOTKZuKuYx/sjkvrq4rMM3VBV
SBG1Hi/yueQUOyindpMerPK3TQE+4KRvo31RbxrZYShHiFYiJIVAbZ6ZuTBR8658EqLMgSenLtt1
Wg7SgxLgroieZItvc+R3v7lMtiDm8RLP8LoSQ8e8ofzESWY6QJtqLQDtHVsXseYSdN77aKJy3tuS
ea2pwRYZipjqKpDxTzIyxpbA+dMN/xDewESGPzXlmKKYnNmPgNypBujNWahUTsSvmsu803DnNpAg
FCyylwYjMLzGaims7dzf/N7yrlH2F04Aqq4GuKWIQQx0TcBPRlvr5sGwnlQgxQC0drc/ufYDZgRX
Slu8z5Y6jcggPjofwvAEEtvh5+ZEnWTM+3zJZiaRAQc882sFhBMjjNdriPi358VUpIxaD0+CHLOU
M/TEUZOX7RqJQEOsZeHLqZodTxRQeRQMzwNvEwS9tlc0uoEFotx1PLPIjxHiLQE2oVKLczTix5p3
279uxe0N1Xego84bmwASHN+XM+gsEfz1/AjsqB8KtueBg1wmQc/B5D+dMjDdP1Z+3kpah4D2aZS0
AuWcwa2yny9L3+pyFR8ZZkRL9A0N3pQVkCC0LL/pguqNAAJzk62IzuQEBB5B+Hq1xoJPwSzIhpP9
5nu4oSziN6dETpgR5iP2Ff244lxml7+/aFLzuHY+Z5FJli3iLqNN8jy8rzyA6kLEycC8oJb3j9qp
hcU+Ea6muMGKZhGiL27nGmv/yDok5D5i6usGpw3nQQ63EcuxxpOux2HWWKFzmM/J81gwd5w2XMv/
ZhXcpZVajFdxn7+68S5F+kNncLBYIi15vk5iT2jTkYCGTmJafx6/Y+a1Xl47fAhCTC7TrmPTWv8E
0ve0Ee5c9EF4SHsfoUv9QrM6SAY2grhjM7BMcPjgA3GraJnNGCzFGY5FVIxI3WsBtsGnn8HkMdia
iklE98Z/FC0E7zF/ZErKIZqXKZTpMjIImIFEsRBzI8xLVOAyfm4dIznVt5XZ6NzpEWqYi1s8nX4F
nuUrf6P3si7R3Xdwqbx201jjRrelPcIwzefqtkZINPACRfcajal5h6gDsEo6/3aGVMHCu2yHcy18
kzPWJINMVxS460qLDZBzVJTdMs2XKXTW8kvuHL//6D7lNGxRSUZSRXvwwRNaOHh53oP8AXWZR9mi
8kx6If6C9L5xMly+5wewmttae8/vwFMkhVE2P8FqiBGkt9DsJuiSysX3epE+6mwUsrEkDv7drXTn
dLaUXQjayNsOjPpKzZUlyh163nqkTD+P1Bwkdp4GAqqBay3hN+wzLDDQFiQN7/Qm8G5bJQA2zN1F
Audwj3ueTFIyCj168xkgjR3Pjan/WnCrobME08mjMGp6NPXjY+gLuVL+PKxmSkWsizHDnQi6I8CV
aJL2qjETqiDiFTIJTCWcQKXFvkZsaWNjN1ce/HXWFkMuxZi7kywBWFU8sTq9zwNS54iaKssF+Dp8
ZOovmhscLocJRTeMz94aetRKYsXbMfX/ITqlG7HT/ZT66AzsPM5KJjGnEz0hQ+w1oWTVnuCg3pud
a8UShDdSFY3N+YhkmwV0nQk1dCHbtdXtu5CIFr0667H/t0SATqE2iEZ8aDy1sqVaF/c6IObxy3xU
p4sYQoNqK1oeg9tcC6JTfLcitUOiR7WKnP7QveABdxvqgmBHUcoaQqewVtDAEByJmHSdIA75CqUj
rF63lZ/SDZSgJsOVJoAVyZSDD2J1CdBpLiLJLfW5rdJ/hRtMGH773SAoNWU5nzaM+EBxo5UBSpIu
X8F610XyEGSzFPZ6FEopHBi0V4zDsEQYoRvFk0IOGSYmY1apiNEFNww0PwgMjqC1Q/WUpGkyKOh6
Sq0TTGDP4IPwgc+TlWGXTZiIaBQpNb85q9AQzEqmJ1AQHrTnn3N1gw4uIZ9scTS9zyv4iMrjngv6
LVDNz1YbAJcsk/Y8k3PxnX8WZ6lPgZ18oXG5p2Qu+TAAfVONunAkFfN3Jf2PM5mScIweMl40nrHx
Succ8gpHBceHJ4XfhbhY+OMWZrlePhksQHSRPXemc74JI0tDRuibd+YxUpqQV3KTNRM9oNUUgl8T
hcLO6o+hQNGd6t7tpxGrq7YEFozemx3c+AW6SZRV1O6glQJ49Nk9t1WYx6OSKg7hTl4tDAlMLw+R
0rKiTGPLVa8gbf65IUeS32c2x7AwICbU9FTIRDakkj59wwzBkpdMUvRUmMbHPSxscwdreEL8arMS
GIJBcGqwY90tyhC/ahZ8leBqPnKLJKD19/wVsbXubGYQhqXCBSUe5iYH6p2YgeU0dXaGRVTvA+SU
cPTRWVsnr6m5uNMA6YO0nEVkC/wQz9W5elWnakwupk/EFF2HBOjQ3l8M197/gwcyLKXi5JqoBLFJ
EjeWFb1xS0JIlzh7ukq5aLbLffyFB13ca2j5rLEySMrEU7Eek29ieShVpmXB1uxxDoknaTi3KxqC
TDZsNXkhGZLHipFzyUDQqdpocAVjXir5WP4S0Grq+hu+vG2naBLGfjTKX/VGrKdA4KdGQZeu0Xqr
exh9BicV4P35xhNgox8bZRSWLujpi85M4oMpILmk+2o4v19SD59nUf4l8BsGr0pBFvFU562O27OB
zA2eruTLNSHq0+u7mwsZvNQ0Pp+UBeiQVotpb6E76+pyXscbTGexCrjabDExE4Qa9a6/SNYgicMT
zfVCqE48an7Q5OdP5pk/4ru1DZXdgIw2JKsejwZICJMfgJYD2UTXFVEAxlv4FCehUPTIVTIufJ4D
p6h4MZ/9Nrwabg77P5fc5GrhhkqYfBD2jeX8JynI/7VQStKgwYceTT36rmIoeLglNouyJqI3sjut
S4YGXBRCH2wiF5Kr17XongfzW0HM4h360GtQehKBP9KwWvU60gPWh2abhsy2UE2jh4CPpbgo2RFB
ILEevSxb88F/BE/gOiscBRa6KoBq9HoFLdt37z+wIyMaFRf3zaNVSINwMjGfAUDbJbtd4QBG3jrO
hNP5y5h7ijW9O9BOGr8dHTvvYNEv4tfXGmDYnFjmVZ4hWpNXs6TOD2sdCyoMuzekHzdDuM1Rnigo
WCgA1zC7h6jUw53YviYgXV21xRef0rPzLGKP/oW8fx9ouGwFkSy5LFWMftO5/g5n4k3elNmYqxbY
VruI8sO4xMKRESdaB12jui1kBIHrtZfBC0TOb/5Jjy2bLhI3Yf7nVVVo5sZWLDY3pAlOVyMwJsmk
0eWHCmkd6KwLM4WBQSF7tsCaauUb8oh4QJwxNPjIxLLrMtLa3WuiUIVYvcCunXKm7dQeWjbs28dV
P2vColHlsBLxUiv1ym5zkrrqe3r9nJlKrDcLmAZ34hLkVcjVqYO/aR9R9S0V+pzcFgolKMaD5gLp
5TW2M43Qxs9p2mENHQHP6091OmTsSHdsGyStyU1bpvr5xY6rLMhOwiZ2Ppz57CTkG/mlWEVClPmq
gSZ3kqmGxYfsyp2hOrzTt9IIb6IursxKcusyFp1hA4hrAe0bOHRTrZJ736C3XglJ5T7+OVn6VB3t
JR3NV2VkqK9YymTFwHlgaqORyJXS3jgiRjmz+T1+LBtOR4WXgk5cPdPuRTVCTtdWHcJKV4T2NZfY
YJ4TDHae8kTtl0krNRBpivE8ASOrSC/USAnyelgUJZUB5jvv4kxfKyNQOOv6nTTspOS5A3SihS8c
vBvEZo0HnUyMxfAsyjWzBTY8R3b+mqDHS6erfzQsZ6Hbo0QRyJzPl2X/SSS4lY/4CXuyn4NRfNxh
3koQ1p+EuWU+OALQH+F4iHdVv52/IzkhF2wrAYw3nV//FH1Hk7KkmmuPZPY4NXgI8tgWgZJYEone
TujooD4zlW7Va0ZLEnurFRe7bPJfsS5xOMqbYfgGdA0oZZZtsLmPleKN3zJoQfcFImMyxndt0C8u
fwXnxjkseIbTI8fyWSYQOaqj7LC+Nrh77wbMAMmuQQ6vHED85FkathW0JKfs0PqpcAW08K5HAt0+
+Ccxf4Va09vNRAS0YeXgfPCjBJz9h+j2RPWMcNIEaz1e1FV6zcBOMYluPExktQm3YA2k0c8R+2Iv
773J1Sqh+yH/nTNg9Xm+XEAPmh85/9kT2lJtWQuH5sy2H5BT5m68xa2/WtArtLWQYqwNUlX89VHR
5UUyvtHjZDyH/G1NxN8IavX8WRX13O09utwqmesKJvz2028jcoYd1jVyc+nFcuNeDQidnI/J2f75
77YHL+Ad1WmJzn+iTHCudkd0nvJQnG4PzY4O+b+ZfC2vT/JhRNmiu+/vADDOTEkn0kWVwbQKm9T/
sHiDWRMqlTVau9vhakoL6yi5uISYx0XoY0ku6nWJJFkp4s/GWe/zB1J3abfMVPuBejX9KCn1jprY
pdGkHl8byz3x5iKW8SLdCbaZtBTYxJpT+qhcJi+rLRnK0a9Yky4fHcd0RVMwNvygggs9RO972OPg
x/oYBehSNDRmC0JrENra2tYSLUZN6xYCdUeJY2g0UHhm2XHt7mKw9SG7ia9tjOZ5LYDGj0Nkcu8m
zwkcNGye8bJ1XA5wtJ+J3CPLC6R0Jg1GjIe66vnOSM7hFcS2Pf3z6m+Mv6pJvTQgeBr6YdmiteFN
N8x70sHFjxaNcLQtR2IcHo0GECm/FMgHC7DIuBvr+B20AtAqhlCMqgujqBvQ1w+R7M0QaQbGZJUV
fktEhbA6xV66ChyIMJoU3e/UX2uldEv+lC7znjxQ+YoXACR75aFgP/PRDxt5CDaH0yXdH1pOr9yi
XhFeuoQx/jFKoKQLxEdezevRl447Od0GMHFXD8xma/fM4gsvrQT7pjanaCgUbmjn9rbByhAt4LmB
rBqJC0r3do3Wad9QIe/ici3hqvEUOzLEvi1d6J6x/TCG+L7A7FTiQ2WAXW4iO/j+iUmSRK5hPdcs
dFu4pmXV/dxMP+4BqVYK17QViNZXZ2LXsbSrHrbEoZWab8LBz3c52E21CZgGyE/w0gruLMDuTTb5
wJsQSFfBWNi/Z4hqH5KyJzTja21kYUDjkHhsvRBMdEFVic1uhATnP2rTvs0prxYk1BwuJgFRY9X9
QHzEIdoXkmSuu+c0ef4ksXlxKCFOLbFfI7v/i1CtvtM3HAXVGoX6wJjgsKvz9bi4vQNRQfO3+LKS
67nbKvXE/K+X08oF+diHTF7JebKYXwSQvaObjDqDtPaPLwzR/2yVjJYMqsHEg2tEtWyfBPqzeV6S
3uDSvXfPI95Q5GreNtFJ0GuzyCOANJuxPF8cJBHfkHW1Z29zSlY4d/ZSwIx5bYSGZZ6VbyD0NWjm
HvIzVmmBEaHWINr/tKz+Hk8vj4jcTgo4D14mW5Zf6tzjS+TBOU/ei18pX9B/++7VkbvdDjbrYoxw
TO6G6ZsrY2jfFBBQOsYfG9MmZ2RnB4Ka/Go5zEDncMm/DRdyy7wk1SqfJyfjPAQu3RJ6aJdGVzjE
0O3OWxajycbSD4WRVX1ZJCg75MG8DP9pZSTH/tkhsrPo+OHUG/dBa5CTdDY5bETSKlXwMzp8XeLj
Ds5zFn2OYN2d86EfGVjW3puH8NuRPAAtCrpKJ07lJR5qaKB2RFp3auIHTUsasZWBkH9loJ+/sFzS
UzoYBVzZ+0z+op3oQ04u7tZF3qjxNpdvAWeLYBVOrLIFGZKQYY+lWTp8CQu0Nbl4mOL4+A5bOO4C
5x9MIalyncZiTRbfbgALFglSWQy8dpgll8khNLY78M6O2QNNnyxYyr4xr/TLPr504vPIiSlbJRtt
C+acYkT8wX2XlyCQBas52j6eYAfdeSes+X2asMAgy7dskVFsfajD2pRc/cTNTFhs9111GqR7aPyZ
dEuKNLkt3AarscanXDQYKbU+JzY9oWNxP4Z8dlfq1m5TWetRH+N6LIVEHeJtmnVC/7STgchtJfvi
LZwNJjbrejvDh7UtObRgDo9GUenGfYw8gDKsunibZYW7u5vgDtc9JazAbkC93ZYKb0nRgCqwubjD
LFR6A0Z7DGjTpCTINQ7Kpy8p98osrFV30ivZhHxK1aboZXh3yjuNJKEZx7Fx3w4qVCZCVl/DteIj
FVo+chqRAd1KuqZxp1C7aLWHOCiwwvCpTzJrJjMXtMOlg6SVkKGfJJGuRBtTiLmo3qCBLsoW3H4L
gcv4WvVMZcou/9pMPGzznT+zAX99neeOUzHx4Lc4npaujwhSu8FyZXGhHk2+fKtRXpz3nXJXWB2f
jVr+NE8KOgpoSGUEnYsxh46m8+JSfJuKanrHWbvTjgl74KGKWh/Ep4NBXNZLOnjjt/x1Bgotj+Cu
tiY0DrB9AVmPhiyvzhmOCyeqiQhHT/lvYCPzDEq+zi9Qav+4DxzQjZ7JI/lBn7aS/FzJ2p4KTyX/
23gVezstsOm1Ci9+mbb4mMBjC0le7BMgrS8yT9JXZy9hyBEaOZJvMHXifGLp//CjZHYuGPX8ys+y
jmWTfy8YdiBsF0lRk5zPu+X1nAlZHMHHVEH62gVx7R4fd/rezXMlkimSUdN8VDzv89ccpHnRLC6u
G6F92RAr1M/IeR7YM/vABJnOQt0KySpNqaLhnrex6IeWI8HiiPsQpaJ5LUHQV55tsUvCk2lJaDJO
IHOc4kMZfiqswdni1fmELvXky+hUPVELTPrvG5cmvwocybcKbUkwZ6EoD7N1rAVVZyb/R5S6mGy+
sIzfv0Cd7YU9eOYP/vD2ryrW5f6Nrn6fONlOiMfTTdpn6g29eJYDagQe9dKjzcbKVyC0zL23goZi
fpv1j0VM5fj+kSoBaYf8FTSm9IlfcnJX9/REFxs/Wsfk2LqwQf6s8pco7KX07nPm8kKmKjxREJ6L
s3vXVfvqV73/mI/DY8T9aNrorPz3EPGJQKnDyREMhy8Bi7NNR80q33KihnmfQhuBEtSRQ0odMoId
lmgMY29jrOSmFkeFuHezPi5WEpU32zWj++TcyAX1xLpbvvK1SSEHfPinVh69way28xXhJgiEo9VO
6CBNZSx+7CtHAdJtG8trUbhnyvGd7cNu5TZwcQNV5OcqroUwaKZWySMqgmKrGLK7qTrlZECFoE4a
njata0E9SLdtGnlmI6A2Xx1Bf3qyZ1T+7p2JEPHg8ztu2LXd9lvmw3KewlamIPLZkghAkIkI2ub4
Sf28ClVjxPbZVwni99G0RJcqdlmvnzPBCxLHXXSjicc2p1hV6Q6SJC354kovzze1pclCl5W/fCmH
s3spsnWm+PTwcL0OnO7c+5glvzqsl7FZg6IvTZKB470ZIibA/D65DzTzBZhh1hL/Q1rBNZFx7RdS
HyooVAtzKyDRUyaGG7Y+5/FGbS5ADIX+1t6TehaBBcxBu1qBmgnqoN9Q9HVi01ENvNABFq3aLqqz
JW4d39ubpbyVS6trOUahXxX6KmBzYhZwPsDiHkoxmI7QIBZ/MnzShfSt4ZwCCBLgMPXZ8o+mgdhA
iRv+0z3I3KIPj8s/cdNrTmgWb8MCvjtp844YJiDYVKgYumehb/sPBD3zyYbuVWQS6km47zZmhPpi
qb2xhk0iajSAScakufFRjDnRMhvQghhtXX0FKNRaFF1YugOiw1HtA0ugwoxD+KBgiuRNR8Otek6s
pJuuDbcxqiTSqSjvxHZ0ggghtbX7NlrCqpO3sCfYRlf8/YZSVDlbkviUmnbmBmF/vZ4VMIT1TTSH
4Zy+eZ5N20yOx49cIbtu8gn+mYrxcZZ0sdUARPm9Br1GpYMg6sVzNT07lTyR07NmLb5IvOP5CuJ+
kyBQoxu6fAVSofKN0iCUbHY8ssnlAF2fPWEKDOpE/tCt023+LsrycsyLJoOXV7zLKmtil2z9Ru8n
iq9gTFjMHg1dWGWBRU960z6JFwM+8j5mVVWK/tm1vMhtXvAWtoPQFfJF2nNzCkRYtUKM8ga01G0K
J3CugCMSgtaqkAQmivGhN0yikO93QAazhGVfNlJjCx756Q2IOBfgHIv5XLK8qCy/NAF/L4qV/ox9
tryLc9vEzMEC36sEXzBVJEZFfRCv/m6bXBR1NpClXQwpkEyStYvZL3osI7h+Wom6hr8VPbOSw3Yj
UXK+M+XzGvjjry4B+wzZSXJ4RWeOt0WFE5emaoF7p62AypMIV/fLU3R0gp8LFGiN6V0gAsp1Vj/0
yjXkol8lRLEjToznjwy5jAkgpuxsI39NuD2pUcF+F3iv31VTtxOGF6wLah1xHNpekjSs0cZ7qNqt
gUh9AC564aaBH6LwB48BeZDkNTzq4mmoZWyqTN26Iq6rBPcOrODQ5LATNQboHqlyyILgrPxdOojx
D9DI9vdez4UG4NE9yP6BNHDyCLpZZy410yS7DznKBIJpHvwE/O9yZ8Y1XDpoycqmC/PHb6M7vd7K
snzGFTF3mb9NKkK08N8dqK+PmKPc3lIiV2kEVYz/+TSYYjinpZZSx2KjzJBvHxXXfXIqM5R5ssSS
ozSrHVsWR1yIAEdcIzbkHqsJIC4ueX5kyRcN18Xc+R4qv9hbA1ETpk1FWuGxOgdRfOCF7rxbMYmW
XwRcCAwwLn+FN5UsT3lV59qnlFd5wjWv2Bh59FxZ0zJI52uXGNzaPwmg0K2LYM+3pW5+XWm+8aSP
XuiS80l6/gYbhGBjoHeOS5wzxcELER2bU/x2AjbxyGfoH8wetOTP7RbApqo5Yb8iMQFIBcvy0HVJ
zZGgPlzJX4qiB+Ggv5YbMmOtkbH7lHAGo4zU2GsEYnB1vAGCxGo/PA/q51fFpg6pt3LlPU0jRklV
DD+7yv8bq5Os6hX3qq/tBGjUNhB1VaH/QY01MTUhvXLYp+ySVsUsrQRdF8pH1GR7s7q/cxoEu8Zx
7Z+XAwjD/oCZtgwhxGBbn1g1lJV6wJyoPFRrY0/G4OdTxkYPF1+Se/YC3y5QGhIFHBptMNpoGJbI
C/9GWNd0bQRo7bf2LvzXstdMenFEy8sVPu3Me2E5PsTuG75V6zIijYXpVikaW8necMDxC6WyXC6H
k85UTdQfgMPcN9r4fJrvs4YCFae3MIlWZ6OBLrkmhNGaRNUgny2tt/pdk6TXqXXKANs+6+3f+LtA
YH98VVNjZh63qTXuN341/8grMZSFZg4Xx66c1vxvv9avC2wU22GApTQ0q6pd131oPOFHvakAM4Gm
wp899JtCuuGHCSzVhwRqMq5283Um/0s3ezfXqypmu06BHBnJFQ/vyzPxLwkP+eXzfVS24PItA7Ex
cFdJGhJyqcCkrVr3GW+ZXjGCoMH5KsTKwlsvb5W3/HZJoi+P7EMiN/vj9uxFd33nmXtGRMYa2Y+6
IcbrzAsRxMpHN6IwAI3X5BwrfXC2IilSg5DTbRfSpKz2MaLTbgX8qmGOMw1Lygj0ykNtgZ4gHqMG
djOJ3/DjpwR4Oi9BvBN6rmc61IvoVNQt5do1YpdRvvtFf5yfmQ7a/tdyTOU3YQdm5aIkg/MIQurK
mARFcYEPsvzC2XZ3q49BYOHmpdyo9pehw0EcA7E1S20CsNbu3J7F+psTz8z0jFLJGncprvKbP268
f8Z6ynEXraNNQHNsyx3rVIFFc9DuAWG7OJyAAeNNwkkVyqOVk3ebAxWKdRgACug8ykDIsEjKPz60
2c7QnfN2s8gAEILphvzpPZIbhewt6S9prHwRnHDQhZ6qQ/8XpXcYuDj5HaWpgjBUsVa8WY383Vjn
u6VcWAqjrwxdX0ONxm8yUIRtNFDKrMFrQPtH9rP6s9xgLMVTlK5k7Kb29dFt7S5uOdBKkbEIj7zu
PKJmfldRmwMd9TugxUDo1rghTmYAn9Tdeic7QIbF1x7qmcqH+514HcTkmUqVxFFG8ueJDiESiZ3j
l2LSKn6bzqS9AEFExxfjqgO/wDCyCOJt4FcpPwCEPLmbBES2k27uMMWb9guaa+4H9rDDWKvGKkOx
p2zdpnuoFS9qS5pFPblsFp5xtEMhYJvwZP9MKtmZ09he80jjGdjT/9f3uNWMewsIxA9k/gMazXzf
axT/c+Hqu0mDHKsj6HServoefYbCV7NeP2dpsTDFxdTbq/Z3cQB5Jz47NTGLHsiiwf/Pe4Kj5oMJ
Kn43ggwps8FC2wLghwCmJjvEWg3gbnN+f4RFtf4waeVXG5WeqLPrsU/PhDrAVRjNJpGwzJjeGSSs
bjzEumUBEa+aWvV670iz6pvfwTwGOcXWQnpPUDvC4ppbl0ycGWg3X37oQmDVKq9ytRdCUUp8u8CY
ei/wZviCiN7SqOI43bad2LWQllOvYg9ruSz/ImA3T5eM4DA0zsqc4uGaqZKNbi6CWeQyCpQrsGmc
WkbQL1JsAG+AYs9LlXEkrrEFWS1LwvI2GfPbLgL8r4ocoauAvUJotqwUtlYdgeuWlsVOuM7BCQju
CuIiOnzO4wukrebcU3r9qiy7rUOpv2v4MUfyxza/4APbSDgDOsQKUXq4uo0lfEUD0M/uQiSTooME
wqVn0mqbSkmZa2iJEeLnaxKWszeHJ4xmQpX+H8f3Cii3EWudDe/6vu783lUtODIOMKOUmLh4MPvr
+QWSywu1iS2IGanCtd3TJqryaN5tMZQ+E72u0aekTMX7FrrU99TLawhFqpsDSbX+FKHYgzAXN1TU
sHO0u/nyzJrPk0iczIOoKAX3cmtqpJyQB/z3HtBWre+wk2ujg7SAljh3RUsC+uDzgMDHpmJ2XvLE
fGxj+A0a0+Tvoa162VttYGM+vW89qZPY2ZmBzty6+1cXVlZImyotQlUaHhmG10GAcuqm5FHHoQ6E
ACNklsi8MxObqMaMo8NBF1caVgxHyXjSDDwrIQPyhLkzs1y9aJPnr3P58yyVgNPJCT0Z+DlE/eUV
MZgncFxMX19z7GYD+UqSkmWYbrAql4SujmKwUx+nQL3Glm7UGaoCqsQ/H9Y4mmfgkhn5cvu0pbxj
bHlZW5faY5bDp7DY8q5pOcxrfBsX5fAuyO38MdjKaL4yTv2oXSPFiffwTWlduflEaI3TIzAA3ve7
AikAJjU/Ak0OobDWpa+FzLflJuIlGXJo40CNrOwatU8wUqZh/b4b+33Zf+Y5qGxnYqfbvfmUzP/S
oM6tUU7ZycmeLKze8z6B+jv2Pw2G7e339117pYvXw3UT6eWbJX3kB+vMau/qVEcKuSLELHkGGGBj
0DbfOVTlIxbv0ANIL+1GzXueuWn2sb+1/dpBh0VjrvfR1BRE2WpF7r3wycxU3N7EoPXEnEbpl54C
zAsu59BUaBZGhZpqfjGoV9r5dCSpGqcbbzeM4tYJs32S1B64/X7Xr6AlnBnMCFAw2P1KMp6dbUA/
lHFalZouqbrFNPNftA0u8HUllWbsDvcDRlkyxMWraWLuqJbKAAcbjVIE4w1l6cilibV4HUvW/Wfd
wSijydQWjQMVXxHd3vcg0V/H8C19rrZaBcvIER7ljjpJvEOTlHsLqtqOF8PkaEEDb0tMDBOZDCWd
vIpheCb2ppPs7bOtKLNYHTOWwwETCxYZ/msWXMO9Xzbz9sh/7D8R3AoIQuXc4et818lAVcwdFtL/
6ScYA5uZbvmKKwYwb29nswkJIcuElDb0YNK8ko5OFP790jAsMe0SeopnHnprqARL4qu0RnLr/bX8
Hm/Rv1F7vp0DcgoWc3XHK2rFW92JXgrwV8oK2tNtxOirBVITfxiEOO+syvaMLU2/U4ps0QX/Hqbl
cmAa47aBlBQYhCyPxgXunUUuj8idzUuCCD20lFJEzoN8hV0IyBq2BmoBvlmWpumyT0Imlzx/xYo8
eSNHVUybH7gYfpLBIWUNys8/0m08imP/9I3T8loFB4HXlWySj9RtR9p+s/rZ4iwNJVD3fufs6VKN
ULTnQwKTx+nVJJRLUJHmppexpPQBtGsbZ0XeXw9P6jvB+GZdq8x24NuV8jO4gRhzsMBcdyjXqOiL
ulhAXyeGKgJ1kBJxXXr7qtEmmu02qeG89vtc/4g8ElElRlRghHTHm0dKBEOi2sj5Bso4Efub0wS3
ThxB+UYDxgS2Ry2HyTCeyDxrJXB0kaY/Lt2NEhmR7SMs9WCMvvIRHh5nk3/naInw9P6XFFnW/AoF
AYKyu/3M30ONgZrg8yEXHNd1yrHCcYesKrEjvsOHBM556QiXq5LBMwVNKw9wmhSfYXXKue1Ura1d
6JU2rdK+FaqdSme/emsrddAk0vJiDXjL3G9f5YkwxztEwi18DEucbgNuQaluAJGPupTvpgoc0Ekr
yOrMDWyDfEA4XCPlLP38uTvBn+s25vX4Feilh8/DQsum6i6oAbqCCBFvpMuhNUEs4mTt5xYT7s4m
0mBTO3iTrpuqiYXLq09VXL8+UZOdEbcvvKK9Yl1at0gRfVUvkmpAHs+re95R5mM/XBuSLOe0Tb4A
kIPciuZz/X2D+B2bCaFuSOiFompaHv9RjQ2IzDt/PTdmXG0Ebxw5po7pm4T0DJpWK4mJcv1JgxGg
0GGLRf2R/2z+Dd7g1T8x4+MT1o8LDnRBKod9qoxfOeUZQkZswDTV5/GdjIh2+sjwEGhAQ930ASFY
hDm+ndMVuJsG8NNDSKy449ttFOnw9TaIhrKtYyXB9uK3jSEl7sq7Kg74znuPZziqvFuTcpCbgrjB
qrmmetkgu3V3k2JTwfmOwEw+Mn6c2hcM1qM2hzMsiB4FWs/3bGOGGaUaxUCp8D8baDmX6hd4g23m
xeY+tQSlcywNpxmc8bej7Y+xUhbvHx8Y6LTooyv8LnJpQmPaUNdNRhYSNMOcRTxyUWrUuyVZoPZd
8O4jqFAsi5jWFD06jGss0CNu8n7tVPCj1ghdHgk4AwKRK1rS+ykYH1FUu/HAf4kt/s2BV97phIeG
+VL7gc4X6lc40OKkIKc09dGSIKsJudNUxFAnleyza0mR2j1r4tDf8buC9wVXcFhWEv5ejBcN+YGa
adLNlpTe9Ttsxi1oQM/dmpQ1GOrZT/RPmSquxJY46F79aJ2gGLWjPJPgSPpB492P7rXV9/QDjVoS
sTI2iTvCU8HCEeAhYBTRwDr4eUGA3+cSY92uHRpJzx+SFmdk7sLP8Y+Dk/egOvK6bCngGPO1RIRQ
T/XzoSNA6rAJZOue/s4272dfS/vqEmz6AMgLzXlNkFy2iO6OsiJjZFWj5Rnim6PrEyr6UdtecIZ4
yuFTxJC7trbyhs10488DuyK9oFo1CoRohWR6LDoC2nQapcXW1k8KTnvQz1y5697SKFruCyxhwU0j
HNIUrkiTapoNB9nmAWPZ71UDk86J9A/VetUVNT3Wwh1sCO35RSpCc2goxoIIOn/GXuRkbQ+5MVwz
MOm3VZE39aqPjuJvvEsVzGu1ZgBOCfzCMA3v/S8nN04/T8dTImDMj0RrFUlgfRsRetINWfHyoTCL
rRXlgEDVBVzejCTLE3fRtU3IpPkeV79DMZKPJmIDWQGxULOhZdSaLgPTpMsdV/N7CO18j2C8kbV0
2F0YV15O5Y8zaUQqBqVvCA0kzG2OFiKlZYR2ncc6Gv6S7TNLXkcz4vVSArslQJYdNRJmsmkNjBIU
iYx1+Z3coCDwSiHgEm8+3s1TN22ReTQROX0VjJJ02X3S8NW3cbeU/dDf9SaIoBqJcQ9EwfjtSHyX
8bCW5e0iShawNT9xfzmaugu3q6B3XWNyHvOavq0gbT9Lldnv63XWauLa1/FIUl6SIvfG5bMHIJNx
qE0HaKr3rzV3dJxlyXxEPsKoKie+u71u9ZU0V10OOLzQnm+A3GjeBA5Cb/5xAnfI7ki5oBxRqD9s
Wwx8ojZgg2hDNx+clOB7LpRDA3m0KJEjJN4qZrVCbx6Ncb1RafKkl7D4R5Dh3q/1ShFbPNPgY8L6
77gKk7i13M8s3j6aC4PZ02C9k2Xnr2pdAunSXo8iqc+sUhAGr0cEDtYG11aEmsHTeFVgd8WAy2nk
gVXTL3O0n/Wdtxh9hNaPX5IML55upEomhF6NnbtUs+2X6LDQG9T/BggqruQjL+iH0AjYdnGQ7wgP
FT5qy4BZI7Q6iHv20WOWS1lO7EyA2n9ls4OM+LUTkPdh6nd9M75qIhg66SqTpYEGnc1+cvpQ8vtT
CY2Dv1yhjs7K8YiVR3sfT43e2upgepymrBBCJ5x+GAi+wZNY0sbzfeHJ5RGa/Z++z1VSBSsGySB9
zAOG2mD7exubbFDMGxprwpVb5Hhm/H7MWPltAE3dtDwfjuacc1Qv5WHm3ziqrzhVQR9WmFoRzKdm
ZX3fwjdZIZf55ouExGDGQaYk6EV/A9PtbF/4UkFxTPa+f15fI8zZ8eFZ/3Xf4fekiNHvJImUwyS/
fPR810MU61wFy+qlczAAozivPxVmYFHA/A1gpf6oAUfr6umBTVeBKS2OGVKe6ieydsYH+UO5ZhyR
khzEbYZO+KdDFwMdFCPiMV6S7PxrB6twmjKe6jik5Esl/4lq7JLMJOonRJE1zn/QNFMISQy85VDN
9Pt0rTYSAiceg6J9O24CgZgw0gKHm+jBgyZ+Q8gnvJbm3jD9oX2mvMZQwk0ZOSMCMe9epIW+OXCs
4SGukoV27gIdlJjA1umDthFwV5Jlhj8Pv8Ue+YBJdsrks3n6rnQFpH1Jy6s+EKO4RZQtriNFy8fS
faSeMdRcj7gjphbFiLGZ5IFHP5am3eKU2M4K/2G/aOym5TRS4qXQJHmL6HuUbfWfiiHc+n3lu200
kzrY+ZTOii2PoNQXxP4f1qZWpoRZjfe1ikJg5qNJHCr4OxYs9lfwWQACXen6rnsqbhHsseZR3IOy
xOa8P4+d/3FJ9KDeIqzDjLQRPDJMyh5Tq67YVA43xdmAvTbm+bctKlzEIYfo8RGz93WMV/tfpshZ
VKzYrQhjyf1V8U1B+NWvP6myC9AAhJBRNyEJ3cULuNGzB0no3o4OEY+P6G803imVg5i4/UkixloC
wQWc8/LbrSBJJbNeg8pONmuMqbUZAFa67Yng5gumzHKXBq9WZlOce1pV8IW1iBykIV9GggadsgAB
CtMaa87vwQxrwtiKknq56UTzNEQF9vcf3FGd+z5Hczf9fZYjYsv8xeNNr1gHdP0TW+tTx7B0vfkg
Zx/xJH2p9dt2ET9wqAi0Gh5XvpyjU+yt+cFMnxAfXKHOP+lODfQvKWKvD1NQ187f8V5tuR8yjciN
HvNVV52w3WmWWRq6p/J2iTlqYGdVVKztPZGcfMmhaDzeQJNGBHUDFzy0s/pyPS+JDLxvgOO7OnLI
bGfXDucqbV8Ey9a3HGJ+lf+pYrDeVbufySJi8AofChWd7kMGyIGGAkMk4Gr53SAbbfJUVAgsn9Vh
Kg/CxA5B/5nG1N8txYRz9ldVh5cQbFxJrh8fIpjKGMy4cytTC8TkLozxkZnnfK5Z7ydpVwtIV+yH
CevCsYS83wKTnhQKO1EdO4M8KFSouuDnPuLaL9cO+RPRpvX4gDxCD32BUlGzsFCSb+WIx8uGWHww
TJ0z5Jir777R//QEY6U109pO0724UoBF/wg0etLV1YzxSlzqQRaeLEUDKRFBvOoNKf/NfT/lX9PH
q5K+AkXEn9MoIw45ykBAxgN9zsw6WfHa94FpesS7yer1oaeTdpqKVUX+PoNVQ1/SFrl+UHveU33j
pZyawttc70TGtQOBUSqwqtC6BmdQaS2xXWeVJw2kLnhXRLPf9MybkyOc1nuz7n5oZ7v2m4Wdz9Th
7Go/c1zu8cDTXFrqo+QYZnqPz/NQ5QBRsLMW9M0DX2uH+1GHNEE7uCQuTOYqyh8Nd/SnfbvgMSEv
TCGiSASax7tIcbmNzYcctWhxzPGOcnry0aOd+lqSlrQkIMEb4uqafiS4EtlPxC/JkDqREWVCh2as
bY6Ulg84nYtmiXbQbiESuSnqX4IN8TUqpN44wee2BIxjKxqWUlQBFcAS4xd1q6/Lgsf7qv2W87cM
eRIaqFzugh57ywd+hRUvpNB94+UMouwoJsT2S2OnRjQR+EwO91wGE6aixMk6TPEmrouw2QlkSx8M
omk4lYtAMqp9InHvy9Kpl9FvcCNC9ysIDCIWBjb+jy59ZL+MAXQ3O6DZ/lo6I7wNid0NhmpHw2I2
n9tzFzCHNAA+BdooiQEdgQOEPXCjzH5N0/f6/d/bJElAXPMluyW+KW7lXrOVVSA7uMxWgkRVPQvF
sFWwwMB4AsyRc1Plw6aDgbutZSjDfLwkaAQoMqtghmslHwPY5ams3L/hQVR8P9lBHQgzSZO3cMl2
GXV8hw/sTou3W9LoWaXfoZ/AZKNZFqkr6TyeE117NviLc8nVnUFj9DbQWQQN9bejHHtip+Gm0VlI
b0MZu9IPL4tST3+RXpJuLNHXaaDrihqtbBjF1bNXjSsC9V6bHZiHFe6TSAm6YVXNK/KknwaWspf5
v/9yED0EWLQCTWHR7+LUagxj7V+dmSNrhHiFtUumg9AJhDSpJFAMzZVp3RhIBOdNDMv7O/g3VwPT
DHwVaue+mEhBOG1PbxmDHHXbmcPn8l9Qsqny1GMwU24fPnBK7OedvZ7dIH56kP3qercCrQbmx01i
qcjvAD94ZAyt7g5CKoZPt4fNu65uElbyLXUlvbYBCugWdnRjHQIIwbebfuqbH4dqPLf5NoJi9I1I
mbap9VmrAx01jM6Syv/jb3QtjEfzFl+Bb8IBjs9mtwNlFsD7eBZHVJEupc6LBZ4IVuqdpU5gjn55
aK5x+aXCjtf8Dte4U38/lE06URlOd4S0EjqyJzHP9uhjKZAjYMzsswuinV8vUS+9BHJuOSE0OSx8
C9GEpFkf4bgTFaDh4BL1M3x5h4zEvnj3zXZo2htBOyHUXlrmviJ5CE+hzJ4WpdICkc0F14N9u9PA
YREwBtgdvoTHK0c1MRIxHtUsBVS6pUjdvLjpigEEifX2cgAwkCF/dfPM60GEqHt0PmNnvzIr3D0w
nkelss/fQPmw8J2pOf0UUxh9iwfwABMe3SL/idBTHVmB07VoJDEv9e9KT3i5oFW8QZMkiYgiHsLT
fjQKq46ZEJhRv/OYgNMYn6JDmDS5Qru8NRSBJo/dKFt6BxLmiSDRHjf7W+0h86febhzP+Gmil7/O
k78FFMK3Y5VFWoD5byjpH0FbaTdhxg+Az5MrGc5nqJ+8NFR7M1OToEwkyB/LnHySaYFl5PgJDi5c
6i4q5s+lrGWa6iJj7KW7rDaS8aFnXVPEmD8/kgOh3peOZDLgizsPCqjIXp5QPEK4hdL2smXWQ63J
KDjhAKSbFx8lX/q2CETuNkGtVw77zei5T+J2Lfkb9TeWug2HUsaEsYjcA2kuM9b/NYbkU7nv9C5y
IM6grzzLIT4oF1HVvWG6eLeBUFqmLc7kOT2Sq/+t7AA0hiOX2H18fOFbsyty0NiJzXQICdQ/cEfo
NvLq9TiTlJXvJ1WI3/84PBmTes+0I9CRXHnyo1aRLpPvegsgILBDevnSr1+d3+EIN0rocvh4KPhb
pwQt+FMoPxOSYa1wpWkow5uEidkuAmoU//WZ6V0hdnq47MN12CSUZgr6ybK0nc8Kkxua4bK3HXX0
VK+0+E2HHAz7W5utaukpxgaCtTTL3erDxNSEJQmyrQ8WFdZH5Mw0tVgM3iI/yHfkuQPuPsvZUZKP
+l3trgFDUnwjzT4p7P7uo6WGJ1um94KYYE0xtksUscNZuVeiJpTyBUntYIyYgyJlpuwT4BQEAm2l
kgHEAJO5x4HwQfD5oiZ7DKrjglX5rxWFHGxVdhlpkmuLdoMoHsowJFP8jHpmtPfZgi/4wDCWpjdI
eJpbxQf3d7JciJljFtKO5UZlcnzsM+H5uNHvAVRbV2A0CfmJB8lVy6YuGUEpsULuhh9v3dxtXex8
IlYotBIeQVrhBscxDKBMV0HgH6Cvje1eis8/YKjOMNSvQCm7JPgI9zJbqiSXBwl/0tW5ucYNpdP1
avjqkpM2U4WKK54zic2SvyFHowF3PY7f9SlQlvvr8DTVAaq0oyLgfTedYsk2rNZG6hZyu7+vylEr
iH2gYiyKdlVpELJAdUHdM/ljJRuPFdQxSJ6H2Ctpe3iuOHWn+SREp59mq/fhroP3ra5Pddkal4AC
W7DRpReHQikrdFsJX3hq7/X+4+qy3FzUZ8zFjV4tFBE99rEMiVgOFicsZJ425FWTZk6RTZcPpsQO
8N1KxDNHJUE3RPg96Uf806FwYUfA/+nG3lBYjMNdXxW8uRuBMp8rJkcO+J9aIGjwNPoOGIuK0TVk
7+2zI4KVur0nw0j2rmVz8okW9hl5NblvCA6fj0ir43LY/mC5XiVOhYF5cxVEpZ9YDBl8mD1mdw7L
rVVWSUgsLN97iiz6bQ3QfwdtPZAQLrSIte8m85lN1GcTSeZYqLuYziRQy3huD4KRuCSGtzq+F4pa
5xR0eucHFo8830wlTmN0fdagNUolEiwwHETviBOihc2gszZvUrWM34KoMl7w5Obc3KE8gIZfKn21
uPX6gzh232rNreAZNvjYvpgjhDvtOM9GO3mcrZk4XU2ZNPO6fHTaWlAkBSTmt1dpn+t3YMy/jbYd
riHbJS9B2O+mdAbSAm2VtGfpKd67Z4n3a/1dJlI039YWb9uoe8T5HhBWEKrRTQyGRdAYd+t2vJHO
GfDv9wR9KTSJw844zWMQwZHhW8iFT5iE4wukNoDAjm4Y0xU9GbYjzy1+1vh+fvhRwb95y2tAY0FR
7ppPA0VH3u4OjCk4qiXghXmRo6ihoYwDLst0JbH8adCZdZvNNwMmubaCnltITGfRiSt0MNdlAqmB
8fvrMpP+km8kEjcVSjgdColaoGr8i+xMNJ8gMgeLMBdspYimyTWhb+DFC3pHD3+TI3agNWFME2rS
Qn/00KK4wF7nzOJPTcA6Eb4zqfh37bJmnv/G3k+I/KtI3Dz2WSQ0sBQfOJa2xDbcZMjPSEp5EtS8
7h0P66EP5RPr13CuYOUZlBlOVGuJ5wRaYDCsYGItUeLALTHOMDYWLPKIAE0nqXB26ix5h8lLhkfu
uLHx/v8GL1fhb8nk1Wsuq8H8lH+3DoZO3mcw/K0xvPqu58zGHm7VfuI6TYssYw7bUZYEe4DdFRl8
DmdzphIyuVLRoXR5O0tpART/54VWsKbU/ugWDuaZlLzIXZSQ6lgY+1flj6ScubwUwMVVm/EzTMr3
jIajTUr0YL/o0plfh0frXNl3qtdvnPtGQdm4IgdGCjDdUF2qZG6Ue7Y73qvJb/bUPeKg20SHHU80
fEZbJmi6VPoN1IHUaOhO2AlmsbGEA2jHsG3s1Cu2gHvt+SkESQSy1hwf65MxJodemeXONzhYhJRO
g7qkeKTvLh/36pkALGVfjBbO6Z+e/1XWn+9I/iTwSIw8bqd0QJKhmgdJeS5A7kNvT4q5apqW5i8e
iT/fNkWuR9sROvpSD1l18O7HgT9b+aBEPQLvJ1HuGGR6rMgXGCTBchLkSfq83JiK/6ePSJVeZKf3
948I0cA14LQBKKwb57LnAeAmXT76bMtpSjUtN5MNwZ4RVrQctaRZFN7QFZnQ1VdlrSI8bAmhrZ7j
PlQb6LI0vVv19ipTgQPKMVrBJu1TjQ5PCajpPX+0ZVPjZs2/MIzgSLu0NSFWKBs53WH13K3ir9EF
8JcKycpq3fd6sPK09swx9sqp+zKkH9SSbkxXuZRY1nngot12sz5Va0stgjYOc98kseECACjzg29m
nZIM9gCpzkxt4TTSOz+GdT/fFacz939TXbW0oGFa9tUVlMw3N0grbCza8MMGP8QxL7g/BY5FHmCj
fFrbSUzqGAdPaXqv1efvyv5C58NZi3xKSaUpSYjK0SVet6hGNOTLHwaNjf+aCwMcjPy7Xr8Ac/RZ
Gn4YJ47OYQ0RTq7hM849keSnchRnRuG5wy3vpKpZUo3EBQIeO+yUzY5RotrpiMhWeyS7yLELFWwD
eTCn1C2vLWQOExdfNJD4LHlCRFf0LNAwFrFbXL3pv8r2eS1dSiWNtrFFgC7ZGnYSLn83yYdgaQrv
9xL2k0gTbrlrVskjniwEKkchIxi30diXKp/6BltaLlcrxm1td65v8J92Myf+Xco6/eXGnGRlvTsI
THbIxyzrTkyyZ7RYctk7zK3TUQfRbbb5gtDhzA6H0HSeqYuGL0Q0yixdG2DG+ZNy0grKTv/6eukm
w+lNzMb4drqHGsU3xFuPg7ClJZ/k4Gv3XgCLE9H0ow5H6pqiW6+b07QpW9k+C22CZvdEKssNPSA8
LhHnMpN4sHn1zqRpB1B/L+bABewLxzI+tKj7cMqZdvg7LiDHtm8TzTZJeAkvhqDL9MqFrVTBdgqH
ZFdME+wjZBp2hErdzLSje96bVRgK3/aZrybhX2u2+W8altpnmXr6+OLtZR/sPgywFmqUvmTU3trq
oQoHXf2iXFIUW7FQb4Q+DH1om6sNr0CUE+3sO+hxEfzryDibXkiS1ZGuQaB2ThvXnqNjAxTOLivK
AKWFUZavdaKtSxRLd1OOx29e1LoLsZASDTTn1iDGrsT3PhDE6rC9KpsnA0UYzMQ223kJrBSZEpAF
n/221JJ4rpm2kRjHl0uXp0V+818WRCsTXw5kPX+z4Jykq6p68FIi7F0QcqBE0c8ABNaHJA7jhla8
M8ATm/hRDd8K5CdLgg/8uCEf7N/LaFNyQF1Y7ZMuQp5zvmu8f/w3O+A8kc9g3yixJsmXiTxscOEf
r/NnG9eD+tQw6wuCGzHcNJom1i1OOeYvFXQlKZ8ED0bMN0ACd9nRxfYz9poWQFrF84z4dLFBXOHD
v4cVq7SbVBh6y7qCYUEaVGnG/OA4R5pC+vIvLHzHfFSBZMbJcide371arQxJ99/CVUpYyY0Dqkr9
hB/KiJRLkEtzVTn4ZL574hxOQ6o31wftv4wrWcqZGkIjN60x0RhqaQaa7HfbPAXbmGM5/eC2LtOk
Ar6HFB0L9GHnComTVU07LdYPhqFaMOG1CU+ej6axm0sk3GLa/mR1sS271T9rzilz7fIxjhW6L5nj
tPGlpYckZCtfoJFt0OlNXNsk5uOTWBljjps1b9fxb1YcpN8EuqGPYw2mDGljyanK+h2ukcpNDwN5
ShmriR05TplDS87crDS0qXJyQby4pyR7guChXuqt0Wtq9ANNPG0t6oEi9BAZj8A1/EGtas6dVCjQ
nCskVVRVS9LU97/+gKdfzbKG7JGFAG+PevcwBKaXSYhod4brqM/KfG2lJ9NzkvO+I5TSWvDkpMIB
VvT9aX4lrNZfX7qchBHWH2wqr51go80/f401izCOmfhs/KTNWivH4uZjEONbkacgbGIGv+VvrQbE
0FKiBCbCgPmxDrCp+X566hMwrLPzLqr+AAkeCteSi9zOxliB7QeOKvYtXr4HvFYE7o9xhGFQsbzW
yLK8xis5ATxEi+WwJ3mWMvJew9V5Snu95uZUojNjRd46fneQ4BypxDoSEmDlWk5aPQdeK+M2dBs/
qvMJimSVkp2q6sXBryBcFhy5ELUdd4DaUTh9qQWC7k+ycGPiLTMBiKV5xSHh+slBN5QPKXLf9Qx1
hvs/HZWfhoEKDmg2MUPvQliRKiB5ADuT6Fa5c0E8lmDkQz7zMdUdV8FIcnmxR86cNS7kzWbO0Hq1
zwkXYJzwhoXyIGUb0j71aqTi9m3HamnYQRw3uM47TZNfpj21t6NQW4HTkOA3eQUXHZouZIyBYxdz
jkQYGI6JyMEXjVrbTgbQIh5i/94HKUbSpLzlvQ0PWhOmUuIKDf7vQhWQgex15pMI4uNS3d3uh4CR
BMmrYNYUrR6TN9e9R8jD/d8mmsO3dFNRW8iqvjnWwRqVMYdVRV8vYQoxmt5P/mdHviZgcQ+/faJE
TeUpXHvsTIOsFYnpaqAn1fAdCEHQ7J3NFAokWsJI2G5jSB9lNxGTMkJjpAzJOKwY1ykqfwZj7dI1
CfDINO4IMuip+DhK9K1z6MP2uAAOUH9PwPHAm+bIrHq//0IRwRR3RMvAMqJ2/1ENmlhhzPvNMK4c
rClRQt6tnW3NQFg9ea9rPRwkEXzNdNdvRI3qalwLqJkxhw1efQdPV+d5/VD1bHb8FaHUCerywLQQ
1tLblH5LS3yMa7v2Vhgz4DFJo61DVAilhLqHaWa3yuyF/IeaJOa60hrKF9KJ8kogJWc+mmTCy2f1
q+q0zNxBxbJ99mU1JLNYXcjFFMl3JGILumRvSdT5Kh9IvicyYQ7KTxVgr5pDF+mV+NJqPDvR9o4w
k4waPlFwXw3H8ZrSsuozKOHyQo/aS0lpdB6J/AS7aHXog0khIQJPcCa7CqWJcNJpJS99ZNkNfHdQ
k+cmyNkbl2t1Qz+ixM96UdzeHJ6iZUlo7NtxvR6E0e0yCYHtMM81TFRXfmegs0r0dL6rPwXruxQM
4Gp+BgYdD5Pd3WIVdXMZ/mCI2UYwPPJaP9WLUGHQyx3Gp3KnbyHKHYNIodtAg9of5RBgAALY7j2R
jCIXG4Nc80HoU4BcNl1NQSwH3dyDiQ/PS3I4EEoBSTMVA8bGxpSX6q+yTjkM0jKRWpHr7iOZ41mZ
7VBhmxXy791LSkp6bNilwH6WEVME0JEcqjovqQJIS4Ycd97PyZEyaDeNab2zKjKXfRB9o9HEZCT7
28JzhGD1yYPUzgqaCyAmPLIpj64qsHt6kA2Fh++A9rYcM9hDU+OsrYkGmXqx6Vvdfg8GNuvEusxD
/Z6Xm452DYEXRhu00eQR9txcaMOs2RsGmE/6tQNiKYt25hLG6k6TM+PYYD5LnxF7RaDZ0GxI2n4n
0G+sXC89dsbzfOV76fuY97t18ItcpGBO9R0FIxKoBpkpXmf3l5cGgUs+52q1Bp9BybzdQ+EMGXSK
PGqVwRWKJ5z7cJ5hHX7amh3umLh9ABdEHrJnT1CLDDfblTxQQ5E1WOBZQz5vMhkP043z4DXOFMM4
hckwNmLncD6pbYZbnPZiXxOm/gg2UQ8kMfNrYh3A1KBvTiMPif+ROZBcUyWim/iayVPj3IsP21IN
RAj8xVzxagyrQLpmYTOGO+uHq/Nz4FJtCeGP6oypY0TTbP2NVldI3TNHhQ0U8gTW8G66GEwm3w+B
iqocmNdEPcwrGH3yM+hOrcqTC8dhEWv1EnW/9KM0M5IG2a7ovPmiXvnGUdAYw8MDPCv1DQigh3ld
lSC3mU9hnfdTmP9Em97A9JvQ5UdchDnv+TrRo87vepHV3ZnsJ9OwCiaazyfquS6T8ONnoW0JWM5j
nDXPhb2R7fnc93IrVzN8RFee3VM0aoHt6AMDwe+CWrh8XFjr8e8lYU3mx9T3gyZsKcNuCGEPgSbO
PNC+dwncK75Dezg6CxR6+crUxwNqKDa0sl29cw74GLkxrg/AbPg6/lCwAO6VORPsm1GwGLUqhTrn
D/PMYCRUJCYxSZPUVQVSNBg/aDQ++mYGY/s4WlfdJaEPT6QNb4e7uz1fQ11BNTw0oxxx3tfqVXBY
aX7YwCX3Jv1a7Madp70SesdjzCqjbLyosr718GfdRhxI4kHDdrdNuujyK/fcvyaF2FLWd1NXdAPG
NpiEuE0kVFZVgAeKUjeAoM1mA2Y/jeHPDDq6ASp7gsKcAKNkziFkE81+CCm5DIVbR6ygF0K77D2X
9E3ZlvReI4TM2WWvf3OkXvQeLQRo0pSlo078cBvJjiPMTmTsfCaqELCoZWWs/zYWO+yN2tO31Zc+
uRyIunflkqxygnfPRLBkhCvS6ZlmgEgRs1DyqWMYFIkN1pJK9GFc8A+fgXcIk5odgC+KpFQtgKZ9
+CYWxjeLf13mN0xd5Eu+4xzd9dCQC1Fg/rxUDTlYT1kIr862qN16IBu32t6j0xpKtD6F+zWM1J4/
I4eyipA8Tig6qjoSCXqMFNcs+PCS0HIPo/NAezIIA/lyWNTuUc9zHF8LKKOCMo4hZceBHpavmJip
bCTQrNTKhsFfwQVVm0R4QUWitM/S7VPQewx+FX/+0XQ01SsIAeqOGk6ZcEhFjCknU70FH6/+sT0X
PJtQI9q7E5MfDMs+3Akgu4QOntoTDH8D2kp1DsWmnz1M7mS9opzfVV/2dNshroMLBLriAWlzBa8P
MbNUQZAfyylUXcKiPn9z0mwEly1kMcWjTaV9S2nNURsBzPrSIkkWqjZUY42EMYDPdGYTRzuXLOC2
yTPY1NFllbsbM4oGitANM04JWlV8mIq4jeFtqUreDvT87ja4yVYPTMcR1ty0Peaf1LCTlnfMxWuK
PKarK2uHMmJvIbcWGC1odty8JS6URiLNA6DW+cC7oRVyse3UFAl79FOt/lR5WgSQnXJ6gf7z3GdC
DOG1GLsVzl0dONrv68mANwGQ4p1mD1xA5ElRjntbC68gvNTroKBDTQnkElY/Zwf/tQQZFOV6uOu5
Ny74XwwM8KkLqomTQpEV4hgm8GcVTmqIfJAF6hI4JVikWxb7W8C782uAorQj4bB7UIyQWoHfpjqv
sj9HJ9in5GdnTq1wfuVGinao6JLzbrYGBrZA3vZrmjo57LKbKQhufjqdlqmLgI/uDqaB22aGYtL6
nKrU0FJ8zpjua6GypclbiHBxwbDSWBG/+S1XWvZFJPQRvnNRnhKYS0EwvV3dBwBherdbai83IGqU
e2aXOEILONIvHxGpiVsVIPicIAAzwVn2XWxbImgm1z0lv81qc9p2BAopz4LcsnOc82OK75eMYqS8
E6s6psVD+a5Wj3KpE1R8+XdL/LRBxtTu4DYgPKq2GpjgZv7s/YN5u0LrBKvjrGu4egOx6IV31uzT
kYrSojNppaBpJPVJPyV/ZwjbQxGRGKQ7kchiyRHqxma8iNp6JtS0fgBQH1GTyaOq8C1ENw3p/9BH
9jl2Or+lserwjpcFXJ14wdhmbbry3srhLzOgTMBPIQ/5EaNPaZ1QMm9WMMJi8E4tgEGs7/XiyMVP
lOGoTu6OaprKzDe0CWU8v6iCoWMPyz5NIWE1KdS1sGM2GhIpCw2n98xdu+3gIjIRE1XjarOL++lC
ujKIq9xlnMjo1FLPh51rSTbL8OSYvtTeE5QKpySymTqEH7c72RCerkY+dpXiG9eUEsMCOIMJUwBd
ijOIi0hWn+0ZLvGNkyGDzddGubf2+cmmvvdcMDzA4l0cryxa2cJqgh4FhokEI39RXljb9kTa0bv/
nksBAmeqILoeBpi4urBjvpHlg3+A7628eSGrErfejSZZTkkkM7TVVKU+kd96L9SsDhXECw4fq0Qc
+IGkkEKFnOChhtsva4+SRs0U087Pj4MttSqhFa2KN8oyJSycjUZAteJsbxb/Ob5YsmZcqs2Vt5fV
7cAfesh3X4rqRlKiXhCdHJsa7f1utj7IXOhJSXZ+tZzWoPbkXjTVW7ri6cLiYspHof4/GhJMgmp9
tkBCyhKoPaGaeeaj7wkca5pbosjpCU7t+x0wOUGnc9k9+eGrd/DdeVha0KHhrYG6jpQmCWLBgdAw
DtBErewvtXhkJEoOyhM+Y5x3+c1HXJmwXFWVrp0P0bGU8nnsHs4puxUn3Xb6YNc3z17Sc7GiAlw4
WWINLGaeNNvGsATWZKT9jCWNqDgoxXw4tOPEAvzEoBPMvrA9XXDs9iguljNnXaKn+XqtATK9bw4R
IqtNGecyZyGBBEIj9xMXUSD+LH7n1ANHwN7FT/ENpVxivY5EMyH+ZNjZVu48178GS7OLaLW5WK0T
e2bpa4HFzCr4S8kZ3FCp+/34LMnkfth3glxfsg5hN81ysBufahJmuM9ra4X38NKIy6XFXSoRsYDw
5JLHcsTN8TT8rki+BTnxum53hMlHWDRnTMPCDZBJO5jwvyo+Om2p01uVU4TenJr6javC8ssQ1sEZ
HR/lm0fTRnJHr8yIuYjByjFahITFwcCLh9RS4O6VbrVz3uqLN+B6HCYOwH+FYXc7i7/5iTjkt2Ql
TmCsWzhImeWhsaVn5/UItgFicsPakBjsQxvO83KvrwPYJhbCs2+Kdtj70U8WRW7c3TqIMSVb479z
11no7N0BsfCO0qB9kuqTMSne1cJZr0iFWULxdMSvbv97XGA8bIVM2l1f7EY92toQY/EvRSEwhPWL
TY5kcfNfD8OrTOXfKQVpoxMq4RBN2pmXjvbGJstnoSO5BASiWEWlLxpwlT2T7Pd24oqlwCd/TSLH
pkJ1vJaCJC9d2wL/D4ShXsRHtWP2ys3bcrmH2tO+FqjlY4O8rUJBZqWWvnKLHDMpik1C8uUUHWuu
SYg9eoqzdY5sQQngCHsvprinliKxwriRlI49K03VTIRjkCuEh4/a496XdgOVCbjdiX/C9Y+WN+lK
aWwZYogcmtBwHexyLM0g3uB0Ng008DOqwNKJ9IBESUGS3fVjpX8H+EEF7kMdTskPGZJM0OtNrRhg
QRM7314JfYG8yTZSpQcBSCbmg3/Nr9tMh6DqNavVuRUnqmCYcgGuCSxS9AJkwri3H7ygpXFnn0UV
k5cuW1v7cNXswPuM1k8f3kdB5gXxm2PA2jsIqtSUp0UlIQ/MK6Epk7oxiNZ437cxaLv0b3e4LuA8
GPkqUi7hNXB7k3nUeUwoT3BNBkMQfTdEBzQlSVQ7lQnOCFK8yCAwC6oajGawpbeGnjGzN62yqo8w
dyMZ20Sloxfmkmk2tWTLKHKacXKD1psvchH+L8ELWZwe1KcqEQEeM9RuLqnEH0sggg2R940My0eP
CrUHN54QoJep8RIP0o3CtvOd5RcbqORasifxtIMv/qTmXoaUClKRIoL9lv8ApmJGC4jfipWa/DIt
IxW9qGgXsHXrBhk/5JMoryluG7yhGZC5L0lNy4gddUn4lVStcQMZ+X7TaogStgS8yAl3bDkPB90V
WYEqeJf5Gmh2EAWuJt2M2x0DtjSMczZ97xYMbOVAksxkd1j9cQTx/FYSJbAkS/FIl4sLIYDCFAx+
APByjnuVOg4wjy16QShrCbPlgFh8P8W6mxqbdvbhkAes8fNgHmynSR00FmmEIbIYk/14gR2ngh13
1qioQJpp0/k7GGRebwKqo89Bh5NfW/who5xPEu+xX+TiHuZ2syZ4RrGwJ8mFMwStG39+DuAYCQsB
Bd92Sot0VFRvdQSa5Sj07Us+sh2S+Py6qa8Z93JUk30zUqKeV+1POZqydvSBp7W9OP55Km0cMutH
WM1Kk5XT0mFAR+8fx9jZAGg2nCnS+7Lrk2w8TMFtgCRONgk3+86qfU0Go0sqF1P1VgIiVOsc2MBN
fxXhLv1qtN7Moon0gnYdFK7xfBWj++Ls74iGkjJ+ueaW7Vak1Z8y18lXx0W5TMHqIKwgkClJn4H9
xnSwp0d01KHMzGshdyx1sxuEYTgYSbBGpweOEgUOcOD/IvGnJSrjMgkGiwRKK+Wq38uKeTYKyS+v
d8uCmbefLlXV3hn7BzRJdWPdU5zzo179x6Soyy6qhgb4qF3IyF+T6bKGbMSZKx6AhhyN/lmB61Op
cq8lRc4C4NalhbzQqcH76Z6qa0nu/lBL041v4sIlJgaL8xzPMj/7420ffFbD8D2PxAQBq0tzv7ph
QdJWxEfSQNDF+EbXHNJ8793XlfomMD8PM9lPSp+N+ESxL24p2iWfIUW79GQ7+rIUHyVXmN5n3k0o
UyKcJ+zsuy/S4g5alypXSCs8CUtAyUFbLC4vWaB88ijV1bqzsL5RoQEp7TlgEBzw1uAHuhxGwEk6
IztPVnfgOq6MnSPDlvQxsPiq5KdQFUvL22aBTgNK15vxe8d/N3MipATayGb1BbgCmanY58d0jYTw
rV0SFJoqKHEtZSs2AUPnRtfptUDbHbyJ+0Bu87VGTAmGDSvVhZKIzkkkZ1/35vdp4s1MLUkfdVKy
ggnnadqe1Ub+AxNQzP8JG2xpzh6IM7nHER/9RsVSbIGizw9jbeUTDKEkaXsz4UpWbeuBbGQppz7Y
RGmDzh/+WaBABGq0C23OwuzJYWLdeAF33uikX34edYnLUHcF+BHkrYwy+gXUS1dSqvudscoU+r+S
k7c87jd99KRFOVkDDETa0jtD3NRLHAx8tybL+u2ZMhGsWUk/NrjGx4zGHZCjbJBmULUsFrCzoVmR
GpO3b6+0CwTi184NWYqADeKP6Me4VaUWH6aLJL2gL+hSe0K/vENtu465JzCJjpVKxf0gou2TBunm
vdJ99GDIrLRrTz5oyjnI6+qGOBEDi+0t0zwvW4B2IcPYWBZo9jLcDOT034UNcdxrr9lcCQqREVtI
PtXm2nUfyNC4ebu5xOoMuv93KwLB/MUSxPXlwgla7LxwZJBOaYoj33o6UQzAyyxNeQqf+AB4S41M
hDrgPL8/PTBIp1+bSsap7PMfj4zlNx9qF7VmZhw4MYE6TUt2Car1eah9g3QJHrFQboGPHkqiEl+C
/mCkbLxqqNTTgw9ftIx88TmXWZgc3bR7b+8goNj9tIyhVIqy3wBr38wD+UqB8FijIE3Oh8gG9s8D
QZBdSy4MPGoq0Gqg6woYaf4KwVJKfF5W8PuCF825AA7N3re+cXVOdIfGfj5SF/oDjDx6V4rAfiNs
Lh9B38t6D4EnTFbnu2ir74LZXYhDHc+qKCzkm2Wp0B5J3biBgI4reE6IrQm4AQCS6xXqDXsTh4kP
QEj0u24aW7pHqUotWZlAKBg+NV5cOzVEkWz2VZ1VAZyq1mzs3Ruk8sfNMQ1j4cEDln1d+aleLJoa
SRYA7O6F3MDPjbuB+F1cag0o6KnIDhmQWW0cAy5YWTI5LyGCOxmUPPmWUey8B9qiWrePpfNofOhq
zMh2UjHa7ZqzY6QDghIdP6c18wYW+0aJiL8yEQBnWKye0ZrlWQWQABiJhBB6XZDhQWQo64pXHB0U
o6spx/mcE8Pf3IRVY8EvD5hIZqhGBgzAISqjZ1W68hPCznhVltefOHmCn7npgI72dUgs33zPhQS0
bdWqcGRaLpZMikBpTKr8YguktJZV3iyX1wa5eYAJPP3wuOEyqICP6V4eYRXcmOeeIw4/oyBwI2N8
r0Mu/bERhQigc4JoRbOadcFnNdXapiYrnpUE64JcKko+/kGz4iH9yZTOMmNUgnvZOuO3ArA8q3MT
hLf5Mlalx+YCsEnK0OvKznKxn8rtSWVWs3EV0SoXq+WSEyzMmNaxhWd2NtAxFeoBJOqStcBh0ZXy
JIFO2gtWmvPSfvZtPVkuyvhykRvAvpan8JsfSjn7GsxFwENLSPhhe6a29Law8h7HKjGD7K75rOeH
ES5NtBjqkPgmiTGbe4CVW633ZYayYM6CmZ40ZR9kHbuYvQa1EUFbjD++Y4zNrRSGTo7HOl3Y1qPz
xDVf4L1JdQv9XE9quQ4HefjWXW+HYJTzGXz1RVilsXW1aNwYDeOfU7eU6ZMWoSteX1WdjbOc/VO+
YT5JNGnqAYZrV42kGjiARYMisadImSMecKl8jF37utEMa+CZ9Qf44wSRvy+6aNNHvxGNNZEyWTPP
KJk1xMgbyLQfc8xnJO3gSbI4iLfn1X1nUemkvoMGj0ZItjj3AFdvs/WsJYanm/3P8KCGHZFM/ayj
wndwRSOEi8tXy4r1QowdPn+opr9tx9F8lG6Xi0dz0FgFaW6Vfv7ce6I49BneWw/eM4+OnERG46dq
KJ5zFKWZPXq+DTuoIY3iUWK9JXFa6lA3EQEm2lvUayAC36KX7/+IFP7bhCfx/IVwZpGBNq93Jw3o
mHBDRrY2HgTdpq/3CNpC+XT659CUAB7qsScEXu0PgzTCDWQ59mKUr7pYwk4lmTV2RvHUr7nmDAuA
8C/wRqfgTjSeg/oncDHOgsFP3GKwzNswu18JYaCpTTRY1xJ7xrZ1qwfZUHSc/YtmwR5P6E+HS/2j
4E4H1l14wmP+nyFYfJJEggJmO3z7UZ3k857WoUkrgYSecsDPK+uJZ94zlZuEoOz2Q/SCoPCYwdCg
UVMSPZzLA0Ok0WnmU3IawOT8BL3rlCvXAr4w4yWudQNDqm7ZuVBTWTymwSskmNCkqVR7mV9Y/0s4
4i1X2cn9wHlEqn1x3Ewz/Po80+wYiCYCtpeuEkk59EaO12J3I+sseseuzEOF9Ea0dZGXvXOfHrgi
qwFEft7jsmgTZbh+9/ZlstCDeXZwbngy8zMcwPy5fcEXiZdcKAsnV/QNlB/ee5lWbfu6r0fjvyWt
8OQlCjm5khSLMjAw0vuTJMFZwJFh+W/vJjeEuaCLSUmQyRnsJxhAnTb1i3qNEAEob0jkTDbZvd6Q
PjLJv2BJOjRvj+i/Vt2NmnQLHvIZjL9OfveTLynGbI0cQ8L3FEL7hFsU96B1o6KV8n7B8ev5zpoT
gvKTmvpIwaAYx9z3DM7kXctbDNx8+QND5ggTGJ8jHHS5xVRJcEF/fRbMPXMlG0thwuK+gDRSBng8
D+Zf6gNfI+Nb24WJwLCA+9VJATk7OMPW7ycZj4zvJNAsH9xHdhzrzH+sgkIlG2xx2Jk3476HV0El
lwu7dgVcXg8w5vXnmroobjotKakhsXcmqojPZpAP/nocBP9/WSyfr9gIzyEakyz2JexLuPuckyey
c7a+1abbIDoFAX8/nTNLAVcXDo/B5H+HIO85wVoHNJh3hYYbxfypp/j75zsNoW5Gwt9XxPwVZZ9f
hJkhnEDQ5CmsGo9M9tZayT28+dSSVZDwvd9HnvbECW+FMDPZe/j9QodTIPc+Cs9E/2RMC1lkMbCW
JxxEmTFXSCjFA0zLp8Ps0FTL0+qnkPou5Pw++azbsy/31mPw+feFL+DuMv0dCwHtRiJXhDSYTn9C
e4/Npe/dnc6rAp0l6uIA0+NflP49APzyIaUm+Opih44rVCaz7ZsMZADl0bNCfEAVwGpts91bKol7
BG4Bq7//FbiLOmKfGCRNr6ruFtQkcKOAl1p5s4AKE/7vSQ1GtbVVboWd+BghuZYQC4KWmr7Tjtjb
geBB5Jy+VTOOg//Ul6H35M1BNbqluCZo2PjWCwCTYN9lc93SY6jp1B6DaIFnvh8tLbHLWkLkEz6F
rhDUhowaKzoUMGOzWLkloLgmzyBA7DP2UCAA1622BgZDLeayVQlwNLjKRiKr2agEH+EemJ50TOeK
sRVSG6aVpNiuhRtUoFfrCRKCiTeDMKgbKcD1bxAJRTcT3MI7yLPKm/ZQ8Z1co4QLQM2ff0gIL913
MBcBpmoVLrfoQPO1vwOEeEX/uKpMghnLAj7BKv+KHgjEBV6gtQtf1pwoExymwvKFrEn6R6OZQnTJ
vIUKyPKJi/m1AhrAgpegPnvosDCh5OQRHzd3v4fp7wLdG55iE438DWu9Whv8FpyyXSTwHI0LkFlz
Zw5Dxge5K3v5uU3LRk9l6n16V+VFTxIUoNGIFqiLqFcfYkoVDx3c1t9WA7IStKbqpG8VgR00YFPx
ZxevArqm4tEyq1qhyDJ17CLcdY/Sd6o/ZPFSx1+u1/uMYm9vzTatedc1owM7v6jbkkXFXKmL3zqE
zveb3j5m8YHn4wL3LKqmnzHdq9KKYP1/uZWykp9DiGX1sQ15XqRnxPgwd3pbbH03bLU85ySxrOHT
qFZncKvgrsmmW0znSb1a+ROE89olcRMFn/rnp26C2Rhg3MkRy/XhgMQN1fG8o3iEVT7HcNW8Z6mk
rX6wfqhmf7NN8TZIq+Iiy9/gpgmrCrZzF7btUPqL7Zuu02D6z0S9NuM/zkqvG1kpBznJBdvEc/qW
VBOyYufTFXGoaPDd6os6g1vIR+k4T1XqYnx6jA3TqsdI+8MOGiY7FoKwyWru5Gae7OJF+emuORW1
dImI+MvqIn1vlDM7xCy2i1VeXzbgRRijaMC/epWQX16VdVrOddlVNTOpKUCTIFzXTQKTxZgeb9CW
3oFhTQ5az+vxBt69nIPmtCWDz682fihL/uzLKyS6KMYIEF5wTD2862q+++1cNX6NPu2tbSTpxn03
g5YbIJ18wF8h3RYxLr6vwi3QAaXZY439Lrh/qfRMnO18gyGC3dZGxbIPHz9spPkAqFJamG6TK2Qv
/zBfyC1xk9j2lNxR5MWBiA8ti1mqwHzh2VdiULbbvRCE9xz4mbCW87vjwhdjf8Qh+G03HRG9VQSL
5QluExhZY3o+1/7yfiFsKcvYeJ4zVSF1KFff8/gnbkwKeP+n1yjmedkFsYgE5wlvkysMGqFmmbj0
U/7InwMB74evzb5z09v9UzrABOvKHbixPcDYGsBwO/HdlhRwJeFXGSxZD5zFtk8J/zaulEqAxJrP
PvDkTAtJS3roFW3P9P4NiMsfM6AJtE4YvaqMWbK4OlxrMaLHZycNh67FZOnA+ER7kXm1D7LaDwm3
a32VLWxm5zi3LRTlrXfbEvxJj31xxh/k86iD4NfFT9j7fcmdYmMyjXZGhPXQ6Hb0JijvSGtUEsHU
6lSsc8xvuIaiQ/LIn92zphIYrDJzBOBrnQs+Xhq6dB4r/3g4MoDrK6JQjTmBJoJJsypMVu+cUsni
FT+Vkn48D4mgAOpT2LsiedJHWTpYTdI3wAsyYt1u1NDSbIHrYVrpiL+7YfXDyyE6QwN4Q7SK/BLC
DT+VzYEX6SKF8TMLlVT8wi2i2mJhc9YREPQqfFZyL/KQq0od7tKAr07h5VcQ14OS8kZfs2zB4RFK
YlIWo0Pg4fS+0rsqifiU0oAcmtsCLvoCVyqkMjFIjZOaMd4R6/CxPjQNuwuH0t/jZM3tZ1snX0zg
Vvd0bLNt8HtJYtJzOzvhk1CAj/jhViNT/as0vzosoD+4e8wgfxulswU7C/UX1sWDtp6glxWS8E6O
/h9nBHaV+dzLoZa4UU1QZIH1mOS+FsSygaGBMASs4xDlxGCKJy1LZMjy1worqfHuYE2A0k+rt0fX
lHsJfLzVmitv6xKnAkWf+XVUiyje+thj6Xv/70RCE0/rGdU+Jefhm7SiVe/ST9d0V/RHEpE/cSvV
+rFMTUR8Gf66nGUttSTL9I58NHP7KoDbZyqwerWqluRXHm99rrJvi/N8+0tefOaAZhy9I0JtEbPr
AMYx0lo9vDsbedv8t/Y0+wpygnS3b5usvCeGMsqpg696apEq81rucLVMKANFRbLPz0j/6r3JWH3A
TeUWPCmhRV2w2cJ9YorQ7DyALESEIJjIRfvUQtwYW072O2JFHJN73Tf2EHphEadnozEyIVvh2+bq
0FiHOmXjRIwAtAt/889oAa/IdcIFIWgmxMnUM4hQX2MDB0MHnJlpsFgsf1HRX6dGsLZxPxIRZY2q
8O6M4VrJtLc+GI5itHfe47lelc5IQDxq/yBl3uzS3WqL89W62M9PsFSIofEh3+4GnYZpUW9RtXDO
q6Qt5OfzHmc3Fs6Jrj5T2RYXYQxltK1e+HT6/HXRNvyw7xjXzJ3AdjRQf/EkJ4YcatEJNkpBQ5ED
bm2dYIoCF1gauy/71cNVbSqrl1HqRQYeY3EANj+uobBo4dOT/2QdfMJpZX3WTUMBDK+3Nt7Bt/9V
vY6uToQgkSFpRCSKG3ahHyvrdd/ZcFcsYn7lxczU8+U7dEwBf77va0Db4Ya22YnUOCsb4nF3oego
mE8tL8EhHYj3narDPGmQQR1ESyFEva9mmT+2ye9Q6KHdSdEN0hWcEjGpakGPejl6LL5QAnnNeco9
v+NuMxk+z+cW7l/4M3wmK/1LPs2b1BHLq4fgMVON/dGeVF/mTV8iZNzOjmx0Q+VmrJjQt2iRSKp8
h7XAXjmcCpmn7VL1oLlVCbfrV76y/XdhYsaZLnQppakgfg+42GcA1TrNSKkbEV2/pnVtFQedkFf8
8bbjWy/GCDSea/c0gw3AKXpv3w2dksJBsqHxThagyGmId4Yet1lA/2H1PSG3suIjMSVybgUwRaFa
Vf80mH3GbsPbjHCmfc4xIIsr6xErGTqjTiWA4bs+grMLrxbdfwsyWYHPsqXB9QIE9VcALhEK1AFR
Zpls64oBkgtiQSS0FWpgwuemDK9Uow3Vh7KpQ3lu9MfOe9yBp4PnUhuoT+92dADNjNBgQQAixejX
njS4bFT2JBpiJJqYatoupopgaUEtsK5X0zvbEn/hPWMztcRtR0BSss3celukkT/Bfjb+X43z1ewO
qMI8N6hnJZM7jMk5vdXAIKFeo3/sYQtgmnSaErSCqjocXUXszQfpUzdDL4XyPeeyRCK9DJAJzZpo
8RVisJM/ZnQPXSSlfYprCVLKoZr8V+MLn4vvl0XjGZVuZ+CdOr/Z27bXmg1aT4obnMrbpL39bgDl
ZG4pyeUApVX2FioElPx6+nF28Iilb/6tCuDDBz/jUcjwKJY+0G3+VqUz28sc0M2itkAwgYK6/DII
plxjjB9Qbh7IQp5d4oqt4sz7MwNCK0IQfp1xj47nC45r8fEiFFove5B8jq6Bu8pMAAr2wBc51Rfr
fzRptmr/uuEbq8vbpvBX1+xHRJyhOY8nO0eImIXvo8HD6FQKKWXS4f4wi53RjvKI26WyBek9kF14
ha8f8OI6wbB4asKTPUs/jgtdh+V6fsywp/oeTN0Osh6gyqwZ+4LQpBLYIB9HieCCsrBBDyH86fhI
N6poOytbf2zuF5RdN/lgJWug+y4MrAeGTKsWxVvFAP1uCKng98ZLRhUSTjngEIXh0H+H1+H4eKKu
q5pGGKKEapgM/zQObl4I5iRW9Do92tbBN8eMyBCkL0kDVNoJmWXq1uEumzMrgpRTES7pgapzIGxJ
UBZUIjuhmD/0B3soQaG3JymWvyc6OAZMRrovp26JzWjmXYmVCy3w4LegMFQZtO/W7ubjnY0bUgsp
KFQByQY4ncNDPkXPlcwLWzn4+p+ni8ZcpOOjDRGsCokEbZe7GGW6zG/B1D9Z85FATq6bqv1F+n1D
RjJM2SeoS9pAW/A02ON1ZlbxNMDJ2z7XA2aVaOtcg8vS0ceott+hl7Nk9N7eEhLNT1v1+MOCyryJ
phFqyxNRtwM56XJGdpE5wtFZJpmv7fQdAZ/6NVfrCS+7TKw0BHN/EJIb/GDFiynGDrSo58w7yILQ
9uSQdNWhw1l0Hedwjz1eIinPY7mPRzFwayq2SCnZssmSEtU0h60J9au1QYtXFRg5Kq0H0FLvy7JX
qj/muthEXbY4XEqt+kIww21rVFx3jHOYWHxhBnAM4a0QFqfGn+IoW7o+yHDkbwlFjgcl1dyPh73S
OFIuSKZeT7OYb1R+D6rk0HrUMJwcLlnVaOn8XWfbLgRDjs5CQVShZDEBHsQbuVn7fXExWz4LVr0Z
CfwwQfCZ37EySNm1PJmshZqfaa8UmNLTI6BpbpuOW+eDspHp7UTPTqulPwyfaGjKlDoS6NAyGks3
wGVMGQME5fVXqQ5Wz31seRS9f/LIW353rrO7i9kGO8N3rqS4AGnftPaAMK/eeQmKst2PuqEL4jP+
GXPcaspqsO1RzdebopWs5YGcGOzDwRzSCmVP1ruGvZW5REFaNHW3gKgq/wMh58LHneRiJQiHQPE4
F2oOYQ0vaysGxmIjta/Pj4kj2dNNcveX5zsBvNYWA/R/RH9kZt6ymxR7PBJhspQrScPefpZxSHat
YXtWxWnn4ecTRMufqyLn19D6E0hj8Ju8bmpEiEGvx8K1NHogc3UwqPfT11f7JuQiLbKRVUJM5jre
BKXScrKVHDRoYmpn74tr57AZuQ+Ky5r5tZYc5rvcyU0VbSkNn0uZbo7Fp1YwqIiTG9RvpwOxAIyH
CF3JNpc5Ge8+T85LjmOLwe6b87FT7qers+jWBy/+eaH+ztXTVd8jGIjNgF8YnT+PNYbiPlwCrwSK
RWhw89JSd2vwiG+XA1A5ANhsen+2LWJQbTiEtRjNRyIXXj08bV6PvO9lVvuxrUqNVVsXzBCFKbyN
rPeFdaRlzbWJBhaSfmGB5El2Zxl8IYC0908GjyWg3v0USIvg9i/D1akuSx4lEnjDgDIT6TWjN8Dy
2B8FYfaQ8HvQDcHkQsQAxIk7Po8qdRca7lrI3SUe8RoMwwnhr/iwbJkZC5OW+G+EZ6HGdFJv4QFq
PwopJgI17v3zKoPS0mHfWyEeLBF8KWM/3s95TicbaJ5nsXBKsZ8JFTlX5PgFxlGejR7IZZZYpE9I
yVytUNw7fkx4TPrTJKB9vJ8c6Vwjbp/sUf+DGLvXSmHd3fBD754gQY6TiddivehOJ9212/4eBg0N
YZWm7zlmajWRODFWrQc8ZyvOg4SILuwDwNeU7AAfOyEqxaEEaqHKiwpcvNDcD66bLAxi8y9QGTcK
+iIZgIZNu3Mm8rTKw8DxITAhLSZyaAEW1czIktnH4koMAWWpdMK4CrkCkcTlzwM1k3vezewL5n+B
uVcfx/HsWvy4n55GuWOWcxJSJI91UnQEqdaaZgtIs1X6nwusm+mhaVjFK6Y1zMO1lgN0pFBXiYTN
Cq97lQLI9aviW13RnPMzbsWbs1EyqTUegkSJleo+ugKzVz8KqxcyxBy60grzmJJsXJR80mjZlv0p
22qhuQXH5U2ajBV6lX74YWagCT6wxIk3vqASp2+klrSC+kZQKmP5aU2gA5zgYHL+i1zQUrU3BWHO
NQHS0cXP4Gy4SyJdVYdSKlzcRV4KIkprwP0sU6JJfrO/2DuO/Mj3+JOCnz+14JW/K8zCOoV7JeTn
+W7OccaZZ5pA7gdngxCP0iXr7I0H9o6nS4/drY81rLh/ZeywAdVBEaRODp2BGiNfqSdq7S05ESkY
96vJ5fKUoTEw90AHki+uIihktNDx7gvr0004n++jfJNFIXouDmYnKyijAu4vUeuw5sQDKAC2yEMW
GNIEzMOokvxNIpFIy+2XceZmwRGmW/9xZ6p7jEX8CnqnIYj3mQrWYqg6oYqiJaeDbvQAVSbaS+k9
YcY220V8EWQZDNYK4Fyk7Y7DQ6s5Rg9g+SWAPxO9h0U1n6Fytun+rvHj7JwOHwwlyzNXKboB6Ozl
S0O1bOm46RlQV4SbDYYhB3wfe9XAiqubdwj6GkMqg+7Qkim7iXYI0XO6nZ5WWNsubBpVwWEgotMl
Ed3HOmi28GYDSl1Ud+Vq8ecxqswoINp1pywQ1ygUz08vlX1ufzE5n7fH+/7Gs65jYhnOl2jUE1Ei
+IEFPsKh8WDsFLTfZloP80wWR7i6aD5cGRfNFcpQgiF2VP+5TC0v+Qc/AU2prCurfT4bt51Zrfhr
4yozJUEfHZn4bnkiwpdwvSE/t3nN216Tg0uFzmNv0wjD46/2oQefeefjS3XmWfEqkqdXscXB5QSo
c6vRSzj8Xrbj2dtpHV17DCleT09s40/D3QVMcXfq9EOC4owbIAojGOpduRR16lSdRcQEQm2o4pzG
KEz81FOck/nB+KupEYlYxn+c/yB6mzscsyRGu9edNgPDwNW0LYK6fDr/d/yxjhve+nLqOHOlMDqR
+vdv8Ac0ue1BS3RewcJGNljG4TjaIS++QUeHPDgCAluX+tIbXjj0aZ5419+bn8BWQXlWhL4lUqGr
MYrwcIvmw+OGyiI1qErf5+tSPhfsF5Xp84YNedLHK9CMdYf6AhIMdlo3c1OJryQlvobp31IlxpqY
EktnuTuD4roqBgFUg7+I5gkOJKx4fS2m1ZZJmMatA94A+i8WUPlGTsOfiSzw1xS4Gl8hQ95OCoAy
AfAPUv7GNc6x5bR7E+PgxR27hU6MA32LUbyy0+L041jTirS+O8tIju0weqRuZFiUhAXdUeWG4pGu
ZzQuCMzgs49vH4YvXscp/nS0GnJuXoPt0PBF0OUsWOSej/3C47EzTYyUcQSMXmdhV9nylbjlZv/w
ex7SQAg1Rxs59fRBz0s4OpAAlR2RCjIiFqyukztLL4RU4bokYlbfum7+faltacNlhhTSEi8hpgQ6
r2Qpe7/At9gpQYeTlPmmtW9yx/q8lYxvsEq6gFCkCBn5pbqJUE+IwOQqMWAy2DVSwlqFDnaZhU4F
OyMfBujVU8E8MeEWQihsPWI4c6KVQvnwa+n6+7FEpW8yV0hgYSYkhlG+6y3LC/9zVsq6/4Y8mZqb
Kj6lZSyOBuwg+qWl+iRuIXS7V962YnTxyWy1u2bsG91e9c0KNVeNzo04QuG7KOS8zQpfaFFCwzLW
HYnp8wgQO+TV/aHYLwQZu2LXJ2FxrOuQ1P8S7Yas1b+bwDRz6ymsmgeQ6nXEXQEcnURWYUqrE1WR
UGbzE0pKaQDQQywQR6z8ZRqs2MVwn2+DV3oZi8F67Zg1S9++d5uc43CY65ujpUr6JFB5CKBx9zAA
ePeRLvNXoW3nL5TKZvXpGeEw9fjyHqTLS2Xa5hDxE4tXkoU/Xv/yxGhd2wbMSuwpQ512VKMF94mN
oKU6V/DYdYTwOyCDtlatYd9owRnW7NUcwYkCuDx9G3nsyohVehSKSqug3ISydf3j0HzhgJxch4ak
Fk0hKblpSNWxAXj0dIc89QBWIs/pUWTGcP5zzW6mR323zdcAP/yfETGHERFD6eL2oZwqZosqx1JS
8gMNc3J/PprT9XFbyQmSXHsRx08ziayt9t3luRM8mWEkVjUJuVvmyRc9gFVKnPCh+JHGHinxpL67
MuX7SCnrZz0j5REnCZnb1EwQGNwA+uiNEsPnd5d/JewY+75Nkbo8uKR3xTIGLxAiURtilyCR2LYI
wVpybeWNG0HlwdO77Mav+yfb538Z9N0tM3DkkOE59Vqcf6CpMB7o3tIoNQNQk4HKmnF1aw/AxwzI
ChSY07jwhs7ItHSZzUV7N6/LW2AsnuBHQGErrBxBjaVDbRiuLsU1Q9OHaICMcu8FmgGtp1jNeJeq
QE9AVQGRddm9VnGldgQ5TXbLtpbkUrSb9SbjWe9aUoIQA625s4HrpEr+yHnKY0cwMy40fTaapWjI
smQJm5K0gUqfP1SkOJRyWXVabk1s9nDMhWWoFBFWidSfCQVd60S1y0kmmpMovF24h1l9hCC7lOGi
RJ9sY1TY3xFp+PoPuqYNl90m6V59tFGlRhRFP2byFu7LATjKWi4xfavpAbHkXK3PsE/iFZrG84Uz
PODWriQLcuOxscd47Yx4Rd1qsPODWADT/mK8B27PaM/3BBoVcP/BbQW/QMZ2Bvu4xzWCQRw82pby
inRzMvFDwLitQgXggg5s15rtyQERlRFqwWKsYf5v94D1dM43J2Eer0SxqAchGryo0nOQlCqiXER1
pG6STvTnzBStxnADgrn0oK0P51nozljSRnwh8CMpIb3T5gJ1B1PWrrpkzTrmWeYe/0FGVm97pj/V
t5Qi2oLz/6gxBoiFId2qb6g4v3AhFaCKimPn6JkaZQXXnjyVD6YCbKElaNuUFnHK51CZhln/JZVg
7LR4P/aVARUWMlbM+2fuRirt91FCMl3zpatjHh9hJzBnqRkxVtAp6J0+jZ6FY7SrVJZznMvYxXyX
QsyR7Lf89cExgZ2peZQFh0nHHUwsIFmPv8t44gjhG9hFCzMtNb0+Zzylb4L1m5vsshAaw9SN91eI
DBcdrrlvuNF1p1T2RjMsiAu1rHxCC9fNm2Jen5bEV7GXM7vz7O8tD2O1pqIVOl9fYE/PSen8/ty7
fo0HWk9PhqsYPsMQqHfI4bfWwnWGwkRZzmKW4JdSpQseABnL1g0Z5tjleX6NUnBgV6uyVFqO382h
2SZCjJeBrixa4d+WQiNN0KqRI1XqIey54XXoiMB1o6Wykm68zyqinorOEQGSbWRLRFKEc3Oo2jZ3
DGmoAmRFhU9PR0FA5oSTJsPUwEDuzCbvHAom6eLMWW6dp4VqYy+udyEdH+gmURrmG8cmAqp/AvY8
xA5xpn5Jx5Fqob/GmBX4GoQiDsFECdShveBi3JDyl47ERmtIANwfLFQqaYknfZ35nN3cVxAXRjMu
SZCHVsKvbjxRgbxRbWPWES5kvbHnTYToPe3xr15bIrlnPQdfqgXzLU8yAXbDSdTe+BVvw5fzbnpp
AwR7xkj8no3nvuoiPUq8HeZtTDEAKCEfEJqRJOBOHTiEfX8qfEQShmASLSqlRGSMXB39z0GrXJIB
97A/8CY84y6FEYe8UNzW5pj8CNbjhNVuEyA5x3vZm4fZxCyQ528GTXaDIjxX8jwC6X4DEXhu6jiP
Y3mRquQPN/0wS8m4JGIGs7mv78NbEBamKGd71YGnBkgEGFdMFzI4X1CRTMaVjDCcwQiJKnn8A+FC
X3FLdzbAQ6MpK/o/xxRZbPoLz7H1lL5fQNRktheSK1TqOn6WS801wINhTz1Kzf8sGz9i6qwAR37v
3bA64Zk9lkent8rG25kmVankdSvq9woFdVXiZnC37ceUSoGmYUFGfTetAtGigUHxSRSsRkwHSwpL
Q9m+tTIh7KfU8puAYl9+eGqXZ2LOjUIt4Ro+Q7Zl4J+nw730iPLVvTxDHBPT5ErTS98j9z7VFwas
/1pEypplLn6eBPHGJ0vlUr/umQRN7E1sdTDgMImpc3RFzYqkPv7okOMgyxc4KIwiwDjlFi7rZBso
Oi54WgI2ZgNLhyEWI+OTVYt4oKWz6ElqEk/4+WqB7XMLdT3bWB9Ytapd/grEwJnqRD2dhSLk5K8Z
omWAcdoDRhasN+gMWYdGOd1rmDRx/GB6HgMfX/qx094b0aTD8oC93nTkFYSaO0HowCLCVlxoEWk6
5KjFv4UGYkcV5O/MckLb7GGjHNBsaOA4cd5la1TCsMb7GIEYFFLdbLxEIvXZvjkoFwNjC+z0MYRC
hNLA6qXeNnsNyjv088w1XPIMsWXNQZxNWv2c2ZT06b45x2DkTESJXIWtWIl8bxuHPq9Vs7w24QZD
IglSfCad/MQKlCdREMHPBGJ3t7Vw4xp4Iy/aggUAOwQbGcN1P4pWTB8lsUSk6qw6Fisf7k0tmJ6I
iZUGY+vsiOpDwlpjW5x8dTIT/LUsNHjh/73lXZIb201M0rZ1t9FQ4yr+B5TAB+0HyPmUmOtfHkmk
6mwy/1YdUAJi+y/6l1MIIXt5wbAYFZAVz4VB9ReG+UTVCIL0roZgdAOPDA36LvlPseRk8CFoSd96
100AVK5ATbbY4vkD9gE9KdHA8MtN2/qJGjz5SN86F9HrjWXCuF7srLcRe2Sh05Zycg1R+47dhxAA
qjvV7HiRdy3sKzcj/L40HZM/V3rgEicb0gFABIrZj9/1BAS4PzBvPgs0EhMWZpZf0ur4XlIJ4siH
xY+k+WCMAtEc2MaN4n6kgbw40GDG6poPGOgOv46Dhn2ZvOL4CgiKOwbO4ePs9TYS2w+CTik4NqXt
nIvQ6IxA2CUf15UUoOAyNhkWBwc9qoDOH6/UlRrfMgMmxSyIRPwbDLcSS1bAOoEjzfjvNiwmmTtE
xKf36vdm/LuuD5YFPzPxVqBewdd4R22ZCWqcqXYtLyZvREkff4kw1B0LJn7HymrrnJ9a87XbC9Vn
0IszbqrLvK/AW0QJaH1aHyvIr0EnTXOZ2gJOu8RReVfhPO4UxsKRaAB4rrmRBBhtC92fQnfpFtdp
PqZDb4fd+WWTgdE/POe1on3bz/08xToOXqFMoZWu+LHpgTwiWP3zd8ysdizscwGpT6tgjovVYlSA
sqPysocptENMs9XPucjKflyYRjAxPuQsL+0RLOKirGYmzUwKFYMeGHN8vg4/CUc7tQxp8zwhnval
qoHVpxXwxjkQhCvQ4InFhJ+la3LeJVbbvZSlmDi3L5DxSwvW4B258wMZj0DlVRNkuyySSb3dV3IL
YNdiXv/3pNYYXNUXQGWVBUBrO4LFeDFGqh6ZL6Flapq5mYTLh15UIiNC7gULgzAc/RGSQczgoq21
Z2silBHzm8+0T1ONWnT6kQXQ1shbum8QOshqsYAnuWW1jNCwnQ82vmN28BdP5795Zz6ezGKur8zI
waqcc14RCGLY6DzR+G2OPrDNGnocD+MiYxdwEGWXugRy/sprxVOReb6nmmD2B8LJ6HPV9weHjd5J
O+9cvxs+H/sxAgH+gnQxxnL37mw9GELHr3bM9ANEaroSElHI7TpUoQL6JvOH10j6FzC7b22Kn4xd
7tuOFi2obh3Y0i0Xp8fENDAavt2jVKwKQRup0bi7LVluywaaDsnL4541Re0VuPUgJJ/HCJDnVKA3
EW+ccUEDpneBvNnlCfppnHLYOMEjLpE36CyB8vUEEFDnLCpaFIyO/T/8Gglatj0/zGGmIUhm5jWE
gUYa/mhnQDpBX0UHTrzZ8ERrIxo90tQJwW559OLp9vt/a2WMRD97HPO/M5rsYhc+MD+/V05WPPxy
zaYIV9tiExyf1rGWYsguP5cluSA16Yde/hqUAbmVsoLAmbYF6qiS0rKjkMHgni/zhgTFjGCUxj9x
Vce0fgduNsPGGE9z55SQ2BCVHbJcViMUymiWolzvDQ+ZBPGnMn+gZvdE+WinkWCKsLNtOzz82yYK
s5670R7ev/HLj9LbH6iBwkMQV4KWfFWY0hnSlvbAEhmygfCUzXpQUNAlYpYsvsvVD0r0/OyXgF0C
KupMqLiazc8qVksnHlo2qe4mddr4vEUWk3W/+heT7/mZ2Iu17HoEx46YSxPfEjQ2Boy/I5hG9lzF
t56AUUpp4ekBcWJsWdMCwFIszYh3alZlF3mEplJ7LVEYoFe19ooCF5JJGFI9RLBM69UH8fK54mw2
P8E/mNtOWhmukVX1A7rVOWrDh8bBSX9QHHKeU9mbikn3979VXAf0pQD3QRAjXRv8YPe9bl11e2IB
n+sc6duBQUnpIvRgcjmqiVNPF6eKSV4VB3zzRVli4MiYpNtKuuYuWPUf7UQ8/pslZ87Lz+MI9OTy
ihfJWdlSrhK2KImZ04RrH1KqfPdrvH0R7/Mn+usxxBEOQoIFJaUSvth8f4AZ4LyUVscVFWsLZott
8kP3F08WasbFobdvSZU5dJoOsI4JbuIjdHbfGkKVNTkMtfAxOijqggc994Azj26NpxHVDmV2X2D9
lBVpk/Qrj5+r0XUDbzI40vdrWXGnL/uoZG0rNf1HYOJGQnE94KO19shEwoYaFdZyuzYig1LMbn/U
cfowLBik4nQtLjNMPNU+MCVat1r2ewCcNUS+/5SyqCRT/ZJcHHTiN/hBiDp6SldCv9lUxujSNJly
oYhP6FXHmRkHHp6KHfvaoqanV1xbOlCFlBny+IKFg4BdZX0WvIC9RfWGEXk9Hrmpn6vjh/MAhIpQ
s7L1LxUgHpza3aYHNDog62mpPHJeCP58iOadB/362xDUXAb6FzBK6WgEAsL88libgr+x6QtJdCJe
RIEBv8F5rr/EwE2UUWLgVKG7eTA3GkTBDQtAORMycqGO35oDuB7zSBv/3DzJdnDAj3yjM8ZhzxNi
u5DnSJqvYjFfqeh+mHRKz36hyzPCxcL2Ykao04Ikd489cgYBA8KO9YyxJ66yPsCrdVxrjpQW8UV1
y0Zfiha1TcfppoOb1K1jA5Hg2RAyKT0ChZctroHTCHaqyNhmSXNlpm7RZHye63SBjxfyAyNNX6AL
82dpYxwqeDJgNes8EGzuIcain8GAOWOmkXoVUU59S0dio6LhCKbDyFOl6c99Ew0Kk2nLNVzkz0bx
F96ikNSnXydSIhKb2im+Z2DJzgF1PEyCIunbiWqffGw4Q0juE7ozQUqq2EKU2lV8UtqdzRglbJPD
ZB/BfAz60CaSnElMxtZSlz0ZmMMFCjfim+9bpAK+VJRQnNG/XzkqLIIc3gvQBLHTJW2hwEl9uLB+
eXqsmVN1iN6DcrC5VZA6ArsOWdQS/ocitYdIE1KOsd8EGlo4BKvVCIBulYsyhYgAdU0G+ZBYFWRK
fJLmvH2vF2uiK6ZOhXXrh1ZjYru40PA6/wnnZlFMgMPzs+KIql0hEC6vkrHZ6BWe6SMDJ6X7+ykL
qcfZJrMSjGgtuKLSFNgl38caD2ZlHpskwUNjL1jAUND7VbtairGHdwVPoQlhm0nnWV5BtXD20aEj
N8dIfZ/TYGhxSfXljqnVWNmToqq3d1UpeA/MWhKaKhKeSnyjBEb9R//8d+ZC4egLlqsyNXSCX7Oi
Fj8E9mZPeOBah+6GuyXPfaR/qRSNba6hatIRaaoASL+ZQ4zNLY8LUL3PulX8Eb575oihUY2sWl8Q
1hZhO/aPyYFlxi422OzBtTdL4hD9/AbTWhtJFel8twDy8kdRlzxdiqRjwhxH7xUz5S02HHRQEm1U
Fk1I5c3lu/xe8pnj8foECguUPBNbZrthzbwG4yjW7tuydFLvq3spbkOsqYkDNZwJQOfBT1+S7d8d
fcuVZi7lZpm2u0/pM5MiYPP3NtnueEiKFqLCGqaS7sdj3QAjnsM3IvWCXeZDoDymE6lJsmVxg/vi
8TdysjyjVjhrF37hI1ZeLU5nEAMbns3s/I3lScxGcqDnxuOi4LHfL4bzRjcU5liSfBWzZGP5kpdu
A/M6jSmFPOs0XUAvJi+v9Vz9zrkl0XCeUVgczkbYhSjkPrcwT70Na8/DdHJRV4i2SwcfGzTBOuQx
1APxR0IP/AHS3jO/FQHUokLMKiLdhPX07XZRodWMgyUaj19ogvDKn7ZlHybBUjzfWAt1S4SRGGac
qrzKd8aGHfHEwviNj6wFyO5YQh9sqLYwxjVCtJfu9JVWSzyUYBtHroi1jryxh/gUND3b7T2sVjLg
dlwBij8fzvXmkwLS3UoJSTCOPyCA6Q4g4o86FEPSv9WY9je/QfvoeW2c4M7jQx4FaCbu4AHpyS7k
lA3d1Jt7vjnyn1c/vcDasdzhJ7NsUz3VGRyWIZyAsYAZwmkVym+6SeXR4gS8n1b++/dPKE9x8jk7
nchvHqjVqZYzRdy4X5E3X3DcPFR5Ys262ohIT+TM0Ix74f0fZ/Hbk5fBNYA0UTZlozwlHZj4Oebq
pdJ2UWBtKkqrLNx/Mx6omWGrTHVpd4Un3567us9z6DnzeZ30cRWwUAr6QXoWMPVpoqNhwI4OQOwj
3Zu708RMVxCwtaIuXRl3VgbJ2bXDV/HIdjHpZQ9CuyiDKDU/9nYnNFriUjbWY/vxzxFrtac9T9jo
BsXDjzazErfgQMl93jOlozVqTwmzYOsCJPqcvpShGjEoYj20HJZ8358luE8Rg8j1rwVR7kAOmnrU
U09357iQYjBn/gn17ozd3iZyYzBgbMrNYhM+DGexSgsmnJDRcH7Gj0nO86LW8pHNuYy8EsDL+99u
GWDihfmvK9qbZdSonD/GkmqOv3umNFn/pkFCYQyrpgnXJGsUNhloUMiGVkN4w3POrNGTQeUB62bi
1Az+8BXZGkOUydJRvqJ1jkZtjEcLN79TqmxZMS0sO6XFMtUGsmNMDTPw1PYdBgCO6zhfJhx0h3p2
r+8oqrOxyrkmWZCf6+88FWJhgjOlpzcQmsjn8cilXyKGRxDSWYlEbDvXgw2V6J5kqy1QvOus5+se
47BrDtqF05tDWv4UNhIHJLdDhxuvoGkl1GWcchi3D25CIquH4gcGxGYOSstA94B+bFRS0XrYUeG8
ju0nhsKLmiW5jqcUx+cZodeZ2+Ctu3OysBZQk6EH8vvCGnH0MsQIiKvqxujCEw6oP734DnuQzwGh
uB8gaGK0AsTYIRhRuETl9CY0Wrwz51PwXSDqorxWtNkLsIrakGRY3TT3EoXSVk6L5OgzEHuWDSTE
BXxGw3f20ricRMSuZwSUyNk2meWRyZw1lVgcTW09/yRhWdFSmuqLDAbse0rHi1JzMamTbtdyL0px
THEhv3w8JpHGXLpDZtCtpxCyKBnaKHZPTyWRvZvNqKMPsqH3M0ILq5lw0VJ3npDDCgTVos3za8+f
gPyuI/SzCpAImM8nM74ZWTGILxQxXwf3gUenYJRv0ClGBJgdgpNtj5oNaR26AC/b8w5KCa5tIm6r
6oHC4uI77qcRB1gZpO0uZCxqb/fc5S+fdxhLjMUrelq4S9EEQil9fRQuz7bXCmelMAw3BIDjN9kT
GkF3oRF74fLOB8BUs20nn2SJwqEoPeeKXB+gkYtECY53h9+aWWxJ5qNvg4vSXKX7OGtNpL6LW6Ab
lwmjPs0Dhz20jMAvH+sTUdsHL2DzHZCeJ6nBHOWNZswMQUOU4a4BnwbCHfj2oXtI2v/LRRQYmtJ1
Ag5fVXNIKxz09TCZ5hQ/l8HfSrA8qVrNU7OM+0IsPqm43mO6FejnDTKm3VX3eAAo6/KZPgt7SWjG
PNC3z2rO/HadKMIDvE2i+ZoJ9yXI+/qqDWLHcymH5zP0PeJyGzfIx9NxOcz+Fha+aVjNSeCI3kjK
CArYBmwhCqXQxwOiJW5AjLRqcectAy0yq7lBXVQ8V6kb7ewYJ8RSmJvf2K9AqMChWdhvPoforSZy
y96nHYITVNkV09CH6a/ziLo8487BkuE6NQ+rEXGs8+10ZkJmkPqHrwcPJQFzDAr4jXsFJUGISrmk
6DoV2w5rjMohgHI8cncIMPhwsMU18speo7z5A7kEZ+81Xusa9AZ32S0puxgUVyliBBHVwy/AW/4a
0lHTb35S//BfGBQtRBvzM8zpktvCsL3FZf7vhxt2op00KOeFzyI9K707TY1zJF6jVC1Jqzfm4Zsp
HEFHQgImh5PuYbW5w0dJhuax4RFUqLS3HKPE/uiJUqu5A79JYQ1DmAGSwFo0mDAYNSOiQJhNPtsh
KC5IepuFzJJ9yu4tkntiRj9PzxHymlbYkeluwA9kIyiGdQvBQLzpxpJZgFVWLNRa/j3cX4u5Yaae
7nzrGVaDLnbt0tfLgz8b4vwGgCAkoVaBRotS0BrS3NnirHRDbSuq3rBMgwqlLA4FpFGSnATRUAQX
yqJDbgEzLSJoXIw06mGmRNpXQ4zlObxfJKM8f/TV2y6moJq4OC+a8xn2M1BepVJ09twUcpO4TQuv
deN2cBmF7O5w61ESAPIHeqLIjy7WJNumRMw9wzhK9drJxAog+4q3Qq8UF6mTEec1FhagIaUSvO8P
PNrrn41HEDwVsvmgaOniy1HOfxJkB97gA45IWWbqqj9mm6lD7MGZMUaD+HvP/pO2maASDpHBJTPf
3y3XykudrYhJ5p4gJSXpTPDA/DE+Q7e1rI4kXbqOwL0UYztFB61fhdt4/SxGUot0ishBMU8fJiHr
mGYJsFZoSeR91E+JvxUn5so7OZ3n/riHhjnPPwKuKOaT+qHxSlbmFXWQ3gLvweXSbp5FpFeuS4YD
m4lKOeWONYvBRgoAYZq9qSv0NGTLhBIhsW8bH+r0eG7Xx7BWcdB1q/E+/I4dEtzEMsb9AzaVlcr5
aqDGN0ILLEMGKHe8rtISaTH4ciZYnvRardiFsRRJttAoAdCI30lVnHi6c4c7V4l/cb0cmbzC/nEf
cd882kFjqUm7pSYMixha47H9VkC7GrmDfZMJozGFU20g5v3JTmFIhksRgZAZ9M5z9aSldm/duT+0
QmcFzrLwIieGYuyIQ0p/5y1MKJeNT+T7sfmJHZE4ujj/ZUs8Y9zNUsUcmZ7acRg0TrL0FzcG7Vd8
4bwPgX3gdeOwfZDaKfK6x3nua74acspExzaCpZw0TeywytcOw7ukOyknLFYJ87y3iIIKiKjTEF2R
JUv4WaqmhQ2DW7m9kVwAB1A/JwnQlwF6WGY+0gO9DhjevLI65Nmy/Oapc+XDbdO4aN2asQlC8qMj
r5h/RpHvyofGxS7G3eprJ4VDuKmuC90LB3KqY+bJMv4nET3LEA86PeOcxEyTqfKFIQ/8Ykf9Da3m
w48xYrP+Q0CkehmTZdPSwY+WPoh6HhoyJvrwya6KYg8vlbEBlr4tm64qxCiLmJ2a92FaA8dExMuV
8oViAaog63yXKJ88LDsdrlqa4YK3H9GdRDt4oWrE8PTcdSJd/m/jALizHWNUgmuXBcMXc9kDKZSR
2NGYW+6zNaXykj+xdy5ZlIMtfTbcnIy2G0JWEUlyfZ/1bsJJksMM574aNw9F8a6ETPKPUmHmf9rA
RVhS5ly9kjsO6gPPDlVFz/nTmuU+m2RvSPls722FACYl1cK4T0alNyCXqpRUiQxiz4+tA2UttPW3
23FPSlHvELBSmOYTy0dCnI2rMO1eS/X0MWb6dIHJBwYfioG7Yemgz9E41TX3JFZXWCLJx7LIxjf1
zODxUGALSwgEfxtQBSp3EH2JqKepIg80bpneqr92snsmDwB8+4lhdIm9WpqPVjbjcMc6smLAQoWr
QencmLzKXs6RcoL5osR/Av+DAgD/nImIAYL7iHDW3PJVU9mwc4TtayA4yKlc7F7naFsVmR7YK4a2
90PGfFxZJyUsuLmirI6SCdXl/5IHETRTRo+DFAISS5Ns7So9PCSZUcp7jz8zFYchmZBfaQw1RvEC
0dIxZsN19ALm+NpxG/livpNJr8JviwlRtkakaNQPJdA9KVO7GGBGZB5egWF3EM2Spd1DDSU8iIay
m7zUHb3JwI69LQXMnni73eXXctTMJAlH6F8So++iLU+MBgaBZKPpoBcJyJXIxe82OXuizLY4x+XW
7Qf2RLqu1styamA7u7YeyTlaUGYMfv+SqzzIGcDeqCJUj/yPPoAJMeGIOI2S13ng/z6mAz0XGdgD
wWY1fDIUXP+x/uqF6jtycKUU9QGSDMjSSAidDkNyGcAzJiYL1QyDwIC6xWtXVjfazgimA5KHUQrv
pTky02sdtMwzwS8p4tcOQc690Q9ZeF65U/fPq6Ic4DkdcOt+R70YPoUMfgHpOJKQefbClL/DuspB
K2nnfhu6+5YF/138MJmpdWYcILfniTXuQZUDzG6/mZwku3zCvsJZnUhhF/rFEfURtUCWZsAwr36A
rZOmjE1FFp57ZxVn3O3K/yVP0lECCVRo2Q3NjeIAvexZKUIzbJScvpdUjyVKTrv3tSJIJJQkS1ib
YP1QCj5x9b0F8UVSWsRi1lFOhYMQ3FwP6LLaIaxSM/JIudFGQvg3pMbth6JgGcUsLJqvjEAh7aux
VYr4aEWVqVCt3AwiuRxTQIH+TONIc9VUYvgD+GJEfHwAYaxXQoiJag9Cv373zT5h93iwQHo92Tal
gnEnw68ZBHuBRE2fTGyIBaFdBcnP6TXbLAehSb/o3rH0KSR1WmFm8wxZVsQ2yyvwjVrN+YlZl2mr
yFSM5ExIMQmk9FSUDjatUvdHceDc9/0Xlw91e2LzN5XziZEK6tzUV7xjaR5b9YCBMqmwEViZ/EhK
f15ibbSxITZKiXvTkgknrBaDGBnJ7NCCQERfEVCaFquMQO4dV2X/+XJu0Ah4sRYYn5Sq/Q4x/yLL
OVcwLyzpc4O9IKxMe0CDBLxGLri0unAvso07zOphRp9OJkubwU8WRL5cXR6XLhIcUGO491a9fJD3
4wWoqT20P4LT2FJ8/bozwiZqWBAWAl/zLjyfwME/+b186DdUzEOP0QnnGbYKLkUfoUz41Kwob9th
7C8enBLzw8DTBG5V21VEt1fAuYjCh6Wmco7u5ieeKCF+iFkkK9NWgvDcWDUR1xqrJAoO8hlatpqS
5Pi/5+mt6QoVAclUBEhbXbCMv1y5LWuSaDnvCqZBtYLjfvAB0qGFaMtsPN4WFRnrvBUtJIJDQVHU
GD5oYpCqzeUXe+yNCUAA7gmrgJJEnqGiq1zT6/iBaLAAw4oLJ0dIadzuMYdi9UlqFwlNons3641p
Fle3IYhv/qhLCpUVsaxUI4EDkbNMV5RCuVnxA3q3oqsgkYI2xIEpdD+LcXCiBtLEROb2qc/786gJ
PFBLodjnTqe9Mp0CnyugczGNa5pUeUZ2ZxEz6nS9qPEfdWwNSwz/fGVVzbCFXU5eQSwKCbGzI8DB
+9KqM/WTvsekBjWaTIil5jYhTfvMFg9Yug9rMgDw6X4bJTOGntYr7aPmwOQJzA7J58Wc/LgQ9OK4
1A4KKjkcvZ6Y3zUMUnGIfQSq6awhR2Ffk9Q1y5B+5ziOVq6sdcebjs6c4jmBmAQTw0P7lC8S8EgK
4kzXefZ9+l/3ev5oMb9xsQe8H3SZ5mmhSVZnKXZCUSl2Rh63xc60NH3NCy9kfBMJuIU+WETo+Jhv
l2cSAVVxtYoANHMGmfOFpPys0As9jHEbBOf1e+IrZC4HfYBBcTBO3svXIgqjiBZLagRsb5lLJ9MI
fOqJA3aQ8Q9QdBH56dlNv/zCs1G41nic526rxs2Dx1xBQHBG5wqR5nqyEzy9UqSM91A94Mgj7rg9
bA1zwqrWdw91DcSGogchWi8N25gPSZ579c7+AH2Fiptkbi+1QzaleciWYY72fd3EJfi8Jd/amhiM
wk2s+VOiaWSQkzdXevXkwyRRUXdxfHkTyw87AnBtN5SdhjQtkCQiuUSPX/t7xpo7P54cyxcuOcZE
tyyLRQMk8WmIJJ2KmWA/qBBxqCt7R05qQqXYI3niXxgTh8ETFHXhhzd5pLmH0qwtF8f85p6FP5h8
8QJhORtr2Vv7Y/lt7rGeX89/e/wOBgICUAiU4q5085v6rATBI8FTjCaFBNuN9dLRUQKalNXViulX
i7RtwgLQmFeC1C5WryCMqNZe6Uumhyk6kEChQy3R4U+KuU4GVq8GbbWlkF0XpnKBeZMWLPwuwBsF
Ztbh+rZF6FzwYsiyjU6PfMXX5NDQ0ZVOEwDuog5idF9D/3L4KSNaqdoqZM/yhkfSg7l8opmr9n38
mjNXIG+tHqybpr0/9xRyFpEBrbGLB+/WUxx9kX0ATcFGAtZxtje2UYyDU0IzMy20CoVzNPAugJlZ
fdQOtluQegPH9VjrWjDRwni8PT6wemwCF6+K9o03pAzhLWmJ44whnh42j9z79UaMfsqTTB5QR/vB
KWOcCknQMx/AA9OEOqdfURdymov3eQT9+r7ESYeZrC8vupagyK2nHd6YU9ho77kUaapyCpVAJ9P+
DEN4gftBxJccWRXC4uNbotp1Bna1kyqdOjkV21avaBoqTVbuAlDjguK4J2Y/uNcndmWKaHUKgel3
OSOb0Xu9HIIDSqxdt5s/YRFGcuZNgNyQGaCl0CsUgVEVAr19kLm3dS23tLUXduD3Z8IPmAkIpUV1
5Oa0nBMP9LrsYoYy4CN4AgU88C5MljumH9wzQdiL/3d7joD9iPEggdpjNJoAPKxjwDLAjkHBsyT6
fmcjFxA44ZlEJNpBUfHAWj3YbQtYT+0DjBlcSTbi3SqzAzR6YP8pFmo4WJr/3Ik91jNGNapCj9HA
1HvDpS6Bb59IRg7vtpG6es5vemx/5hQYrjUjU1xe874ZH1H/3knctfl4q8/5T7wIVP3bgfIt8sWF
GeJTpoJxOXJ++VRq3INVH8c4KrDaud8y3phFtOPNzt6XXC7hpXmXqefQMMchE9+AQSh9Y9giSaum
GDl1w3jLro+5cN+oKA3ul0Re0YIutzDM8Q7KH9LbCd5dWXNpIE0hOi1K7Mx5PlP8k/5nk4zqQ1PY
tdZXZFM3flNkWvD2IX+fCJfUp5FF2NbRw65sxylWytFUxIE1S/Gy3IpQzf0OFhKOTUv6POyK4h/l
cTjA4H45cdmPzNJ+Sx+2yEh9WpWdoueAwFLgVIvDXQ/kKre6eJ6F94hHxDaf9LR9eCvL2vVyHWyJ
NVtG0KAUnK+Ns+pqfiBY6y3x+4/QRVtMhceijLoWhq8sspzY2NV9W1BKeyHSQCudUOldZjV0LMpg
5/FZlR8osEBDAeVD5SAtrpx+js6Q6T8AUzgBNFb67NDTjnPret0S079a53FeaQa7j3bqpRwiqU7a
VnDvFHxOMyqwNRhVmpVHPDekwJAGZ5oBSI+OtajtDjvy1jNk0jQx2hZputT3FKlGQNQsK6J2wPpC
Km21h2P6QdbSYeWnvxG8zQFXZWc0wYKeTppZjZ6cdCx6w1QrrpG+GUKVJFx+L8/00McRy5N1iOqA
G5Fjt+6YdivnDgb+/HR/fqjNvC8v6LItFQ03hg8GphC8CO/nxiGITPxogT5jOZRc7T107O5SrOWd
cjtfQQA83KKYr6VNUH8WPsOYh9RVTG8oMQtI9UjIvYfKPRjra9ejt1af73O6kznRGq90NlhULizb
XsJaNgMOh9jviCItXDKnw4jofGlr1Ag6m44OWg0MoJQxeizIWYA+Bndd6hdP/JPWLtzMHKnwfSRz
oaVanwtNpRExQ4MMdkGHwnX0Ueh4e0MXgRBF40dD+v5k+oONXTo6WLSM6A7KLtn1qJ6huJPezbnS
Eiy+PVAYCyOAeqBVNxuMB3lnIio8/mkwx7E5Zo68UV6qAqVDPrHtM+FISYBy4KDLXJazsSbtpEPn
k+Mzu7AmOvsOPahxsXBTh+hIg64CGKK6zXXB58sWw2NQvOXeoZHLVO/sbGU9SH4NuqzvE7spLHLa
/iown/1ijGLSEPoPRHQbHKaHvwMtzH0twQIY0jKizre33eeY5zc1w2TYlY/aOn4POunAf9sUz7Ct
+JsTMArtTzqyj66FhECf4t7N/LedO+jl1rrvLX4g0RJammyv8TfYWc0x3ixmPEAUM38MRmELvSyJ
X5iSHYlj7+KAPRKXQ4QUfVFIQT9Jq8iAxmG2kyGmQem86enmC8KMGQTyeQnj7MmhD8FfH15HGqgL
VqxAcYv3IlIaiYAr0oXicKpLrThxuAhk81dMENRTYUHq/ww+ciIQAjMpyh0oRoAH4hDwMqitmYui
4SXCTG6vH1fmiE1hc1ds3tIGym4MzoGOcyFd33Ie6wMJn6r55wpt3S3+/Ny35Hr0LH4LHy7mJjjF
mrDOrSMednl3RCQOHYkyvaRNgP6FjSXgE8Rqs1MM3/9pXQFKPgmJQn24N5yI6sYM7/EMEh1MBnMv
ebmUVb7UJbfXzMqDCk8Z5nxPddvdyi0UDfhB9MRDmX+Y2t2YS3qqwK+mxqlEbxCtjRn6neSGCReV
o/yHsb9sEbrKMrv+mZDvB0V9jVvJOBQJqcGEgAQKCaL53dtrrTeEkcQeiCh5subgro1JxrzmtLlD
Twih4DDHrslimLZrWfsVV87wsBZszuK2tNh58yh4hgvVtOPMjef451gJAkd+qQPlmm9Wbk4HI4ZL
PzfazioybGX+2WkGOLDJikudIDIhrL1kde7nRzrc4QUgmnaSbYMB/q/OpV3AC2qGKk0rSlVT57H1
5KsuUZ/mBOm2GR9iHOIhwHLlxbuA+BmEew4z25J0WLsEzyXsekUAKd4q3a9o272mzJYAyO9syGmx
NU84AkPfaa3o0C6d8348sE6Bd6GSXHkLbjcn/9QshpwlZCk2B9cDZjmemoclb6d/jRKUo63Yr2wJ
asK0YzJAfjv6g5LzZ4Q0VJmm73XgAiEmesbSTtgL1C+2DqqJJtpyRz5J1cM+FG+gJ/0RCbM51sQQ
GKZC18QCLazCndgTKoM+eIEHNEHe7F/9mQNQq6r23/u7LWZc7e14EjQck36Qmccx+e5h9nvYIm1a
dqa0l1DTWXnez/QFSipUZLnr7iSto6yUyFFlcVBFzF0ZDr2FC0WKQxIkPgGg/C2ofsUxCctC1oLV
14p7hutX5Xc5pwDrDhnhfHFso6xc6i/PQV9GB44Qh8f1D8aq9vsD9AYIPAs38zKbuPmHWTkS+yDI
xxgx1bDlFWdjn2R2AiWr4YXCbzhA/K697n6HhKmzdODk1ynWWgIam0CMkPzxk06M948kT8TZJaYf
rNWkNwX/hx6aevQZRGs9ZIfqNlb1Gmz/T7/f216kKs3+0bBXFiCPQXxEFczt1lQaPFy4huJ4+0cj
ofSuMpqZizHPLGbsacv43x8vrjLkejgFJtc3JmudQ4UfqXOh3/0YrsOzMLhTaQoXMXDQXIrzy6JN
9gxZdlcxomJ5Dh4xfxCBi97395bmv1VD0fuDCg5NvTn+gDCDg7PBjCq6cmXhrU9ylHkctxmKF7cK
TKAAqRnFSDsHpFfrJljyBRbca7twiVvLjSyLrghfY56zWkkhQt4FRD2QvmuC8fVJPIaxJ+/uxAxD
lo6ju+Jc2iwm7kVBtTZQASycKn7YKtRBsT+jr6j622qM35jxiPzWZY6A7RT4wTg+qIvP6+48Z0mZ
i1BkYEijbUA+N7V9fpDJe66Wa7SYzZasZjskJCb9b3tF0vwPbqxj9HrCO2vbCQfu97BhFku5eIYQ
ignsW5Vg/VBluucvxmwhFi8oQfswMCouqfrhffOHuzuhLh+TIkQYArTyEK+BwtQZfqaneFkRDMvn
j/Tp1c1jrZ8hmgioRavgx8QIgnr50pVhrtsmzvI7wkrpNqFUxSgY3KyHiurpSWj/D+258WDK7k6N
CpCCcM1shMNpsnQ7e2KAtZYh5jNzRvxvWLJR3KlkUmNEm1Ila9NdDehN+DNFt0lQq1EsVFbFd3kp
+sS+ZD+q/3PE9fIwSz6E1BEWf4noRjTqrLekSPzlnChZcnXQp9T7EN//Xto4sJfc68uOlAztlMg/
BY5RdyyiW9fYY5kKhCZEE/mcyy2SGmJMsUW/QkinvHFOoGT387oYsnv6rZw8jHp6oBLYU8IIjsIo
YVrvDmZAvb0K/ZteervRUNAEPx4BIcvJ10gx/t8sfsaUuVjFUbVZ1eONBW7GzFn4gVofL3u2cVKi
7ywXjAvfy3dP0yewR5b46EmyjOt8at5TNYeIrteyjKr1zD4etOv9v5D6TGdC80Y4UwXtwZszIFk7
e1dG73cihHN0ibrXT9zZIhFAZyBpd57o7oybkxyTZEIlCNwZStsx39bfplt8AzBtf3AzpyUxdbCn
DAF9gj7qLl6zGaGawdcOaBg9GgEZ1W9TNxMRTJQTJK5PfF5hstcaDN2wrSvro63MovQfkGppfpbm
AT3lIDbsEfMCj6PYndEy/60qmfntheTs//Le/rvCBtlT57W+EiOOJOJZPEsl4h5tRFvb0HYKTZF1
LMRX+hU4Yhmfxs0JEutOjr5eL/6tHKwU/DuWLykv8G1mYtvgzBmyaHwfrU1Ds5717CkvqXOvCDlu
PfYEB+QyWOVy1xrP/0EMcO9ZoIsSRzgkUoUsYbPRROFY0h2iYiBxPdMbYyONiWvqN3DaFx6/oBXR
W8JqSXZNoxRlqNpw+2HXTk4dJbBQwCbI865np3gYcLjyjB4AKescwgaK6gusJXLHDyHsvdX+dCVx
yzIYV/m/T0bP19WU1RgIx8zO1qCchiUhY9huzlKJCW7+1U7mfpdEKCfXTsDu0OCtab9qsq31WwKM
7OBDgixAdBPIQbHWxzIlW7UbbjhXiM651jHnxHCOHxwMJOtD+Zc0gkzh+Y7hvJIPCVy2DnVymLsw
Qsviz8ap0oKHjztb7qSRSE51BBye2PHazAc53k+m4DglCn60cBIjOOhxc7XQxa0q84R+VwEz/qsS
mcAR0gITWuGn5OSIOJrxLfRkVBc7Rqz2tJ0drKoXBV7ha1A0ObVh2OoBWyrqq9wfxrBzimFpkaBU
cpWGbmO+sS+O4+o1tESm6cR4W4s0+GX1IEMFx+GVMQCYZU33Q0LjRknS/+AnaCAZRD13yBktccdA
wEgoKolSr8BtAL9i8kd3hjTA8nlX9HtUY+BX531gBetXY9a6zYCUQtLpVlfo5zeZc+zzJyjM9DwY
OeYtb5+e2rszdwpxNLMh0l427mYtWYvcfO4Up27O2XIECr7s8XBGI9jTKWvgDHfak4fiBZJbkWmH
Pfg5fpHQA2OykgXjB8lMgihhMWWGrlmsgzoMwJwVcZ/xAAfd75YsFOanunl0k5n0vBoGEnxohCEg
JrfiQwx/LaPEq54ojVJnwK51mtKgo2qxVyiZdrxfoVb/z3O6KHvQUoI7tzLCMftwvK4YAyHtL6ri
gOwesYnssNzvLwyXKNJzgSMxl4Qa/zTNIA6TTB1WZ+jQhvVD0j+agfNeqcYJAGM1UNhX12Blg6a6
0rQfylft6z7rYi1t2OibN68XqmIRmMcZ0EAD58RPlaWUp7gqW6KxS1LSHEeoLML4fZmrHl0UoQCj
PnP/lR7e15gF+plX3CYmc/Har7ZeUhZqbp7bl7+XC5R4+8xXd9OJpex5HQ573g+xDt1aHUU21xqJ
l3LZqF4vHf0iCmf9Ij6lLzle0ulJdIV+E5T6KgK67gZhoZ/pf2e/KqIWdTv5YoS7X1M7Qvv8BpQk
VGM2lk5wRlThMvdLEBJRNVVpVqgPU7gCWlNm6RZN83397MfpvzzMB7H0cl5HsFmJxBjUnKCKXM7g
SetBt9uSnyz+8WHNipwpPBElAmP4VYi2l11OQJQs7ieh6sT87nbyeqenKhxwwkfHt0wZvg84IT6d
K00y+qeAI50ryEDWlumZHkP8F6VFIsF9iB+AE5ZSCGP73yv1/4ZGbREasKDwXOzsPd6eatkfElRR
iRtypl+YhkKv7lg7UbXjAOmyioqw8GP5y5IRK6b0wFK5bSUX6w4woutzEX/8hs5dCt7b69PqxvFD
80NEiCbzukfPJAlD1xdaN6zAcRCn0ePSV2Ezbb9jC9bzV4jIqlUo7sR9ZhOu5/4thirwlXB+izO8
wyMDVvSE3z5bB+ZmW41xv33hvWpsvDoSXVzx975Lb8kKZWQZKg6aa/T6Yc69gsRXmeqhmiCsCG8V
9SvLbVBcZkZK+JQuDilJa5vW6GPzcTgmZZHsANth47EkdueuIdSn1PoVG58/a+kHxLHkJRTLGxEP
L/a+6qG7aVQNzhjyobfGX1ki3OxYcgW5sJKzLKYTE56LMQQprEnGG9ktOjLz+Es/az7WT31N5UNd
x2LQjaYBfK86tl2sQEo7L4Czg/uU6QbRzERynSLlgTCbavihFXaBleLqNk8s/w5hocsMKurnZG4+
5U958GSIRl7+MYq+40Yk4js4o58XBqYjlXfvs5X9DYSz6t44UYWIISQnL4i9ZdzFRq8M2yJSgrvN
5m8gXzdQ/61d/xYSdEdwEZ9l95hI35vb+nN5wvOhcxNuLkv3r00m/dYN67DVwRRgv9UpdYWzQo/H
WosZpZtfvU+BpAPQZJxqLTNq8w5fdOTy4/4PIeVEccuX0KL3qLSl9SEQ+kNjMmAHK+/qAoA+EnLO
nESFpwGA02kJrsFm1jkArEWJQf2mAStNQELr6erCpmIOybhqM43gfe/QhHFWJ65ko7Wc6SDukPES
gvZt6prd6TYIZjbxn8cbEMfU1qRB6qyoXAms8lNZ3XPNkQN7EsyuZLOik61EoCanmAcvufAaZi3T
U0nQoRk3Fs8P/bbicQY0SQFnRB+TpWVQQfphy430/WiHodDzwpujLrXVgHWSdtSZdzVPg3SlWo1s
BKa/ltk3Ycj9SHrqyIDWzO/ikSVwcpg56LWeVlStIphPjq+0sKvVC8peTMEobnRmi4T+RhbQE8wn
S2KRxisWfLL4z4hNi0cTeF29QKk127UHFv/1YN3AOWK6CFyGBgzvTD4Q/EVSKNpPF+AM1w0l8wt0
4i7IxtV1dFZZd+N4sWeDWsOG4NXaSzDBmaT/fIP828zl66SiqxJbneUeZE+9cR7qYmEcamMC1UqI
xO8jNoYiLuIxQolzctZmuInGgi/BnIyXia2QTUXTugAY9SleQVSQH7tj/D/kJK8vG/5ff/JWcY3z
50TfMjtY4MWPyp1dPq+rEpKOuMho1ZFIl2NHgAuVGnu0I6PtkwUxuxvUSEPAukd6Z9MzdzoTHkR2
T9j13MaLvozHYjJG9aqKkmRCmu1DxDdIZ9JNkB1orcRMepyrpnpNP7fbPqX5QVa6zwJFYysAPgC/
y16SMFXbYWaWCacZ/Z1tS75T4hKOhqlfVpH75KOYXF10cgNz+a3r7NzloTna9Lw2V5x4RmbEGTs8
kuJQHYXSO4vrc8BRKaRGW7A8uTxwZYRxzYWYTpAuPGYINn3aTOjtEnTMGtgOvfitHm+viIML0l2Z
Lpe8D8t+zo3C4cNHB9OfQfvSbzvemZcipnOWqLHIIBCRmnE805tKGXIZWnAWj6Pf/FhWVN4zW2Bu
IBhBzzPxnbLO0NxDuEVLWRj1ad69FyMzBK/Xpg5qaQQL2PzweSAbAxpCErperTRpm9taILx5g2O6
yJ/aZYQUK5yXZwUMtRQuqr9f8cD73EGpZVexXBgnwe3P5TpPVE8Qh+60u6mwjHx+yFGpyH+6amVf
ykZr88w3m7Ei7NM4b/pYMOq8t3mnwag0/oRCojf2b9leBlPMOKsR0xHxVT75b3qK4nw16Zwr8W3b
dqpmZ1Bq0U0mU2p6lttCt4howp7oouCj9qG7kX5NHse2ywXXAhMfzQEjV5qbFr1KYWT08jjFIwmx
wESo0FIctQ18Hj5Y3LwoeG5VhRJJCopppfxQ+Soi6BTwwNKjmeZ6JUWaM/phorT4uwQTaefDSzou
X5kg7O5V11ISuAz2beszGC7wpNACfKXB6YTr0w7xXJGzxbx8S+o9Ir+zc3VEmKisuorL2ObWeRaJ
SOnyYgCU9tbaMQ5a7PU8AGIxv1bQnIsFxMOQdd9RwDoKUw+WW9leEPLPTSFjRxlqlsIW0qdzP8Ts
DTFTJhUa7EBvZOcU1Xy1prHUt3l2lJg1Zo5BTBbf0PR3/ItDWltIZRYWmFMiE4JEcfRNthXHz0jy
Q35wgQvuZVeP4f5MEy5kqDD3ooErC3BBIG8eJRPeIUulqEAFaPTAa724DBNxSOcLapaQCg/D6FhK
Y07V8Zwu9qrjt/H1Kko26ePcRPFVQIMp4FcrYd22n0+QgGd3tyBI6SM//rOttse5UaH4q281bRXZ
YHch1BFo5gSnVk5o6IH5yREjoKoZQ9MlaNvhWiD5Y0oWrrBuYMdiQLHh0py2WguvCO47l7BfmuXM
F6oP0vJsAlip4gI3khMCf1usdAkCWNeKQtdvS4hX4xGWaH0yQWuf4Ow4NIYJ8L/FY1UMp6AYGDF6
qqopOG/8vKAOO4msb6iii+H4CP+ituqHwoS01HpajCRSofmxKskHjY9i/NzjdidDgSdSfu36bBIT
NlZ/QhCO/NSl3Q7+pn6QQECSBj7TMjy0/W4ZdS+vpcHDjKeF7NrafezZe26zuda7+7LplvBfdAIf
BnbNOXv9+g7aeHmydYAGGPQsk4JqWznrosnkgT34im2IaSzEAUD9rBhWR0ciZGt0asrLVtrX7l55
aFIJIAwjlD96NDt7xv2hZSL5vWgY17YfXdc4y5XvM6JNrJtlmhiNfpv15rBBqB79+mnVaF828R3Q
TG/dHdc8uVv5XG8Hi+Mj4BVpg3ptGDWwHbzFHhptqCE69CJI9HOd7uT9eoY5A8YUemspQ+ElMD4d
0lfvgFlzIqDxJ8HZLqQ35kosrp54Y/vzEstvEau4CFwMsg3bUytSRgLpSWuP/kk4s11/wz344z64
evgP7CuvYWGfuThjneDLfpOUORO2V6B6x+i3V++PO5HeG7DiMXvLpqYwj66kofpcmxM5385xnsjv
nLz9TKhNCujPpiRAChCLK3GVrt04WUZLJDksjlM4a+Osz2F6rrvDJAIDgH0RRLSR3/jrFkS5sOFS
HchqqInYQFGesiQpszf0bXGTe5PQzYN8rx+RVm1hpMcotvJke6Ln5nijAanaesBNeV4S5KaNac1h
DAMQDl8MW4hcfnkNM2CsELjUNi3CcVL8rDyYVB6KW9CbZiY/PiXYh+PAgvAPl1bMhlFJVNrUbqMJ
l9fLAjzEiPyHEBgK8Mx7V7UMREawjDB4Ii8sUSL3bRK+ung7d8SHzEpQjnnX4sN9G6nFytHZwfss
ZRARydGzk/mAn/bMtBPfv329mLEmNujtj3+ENwaFlhesZxdd4lnRvAAfvynpW3PNFmuEYZMJbH+x
dLt+RhxQHzi9CWNMX4IFMFmevHc6zQSd9YlkBBxeJ5qxzqBdgLDblqmgI7LGHSXkCjoXJqMKoP0K
D1tA2yegyJ9NA7aIAONW7pVQX+pO0PSEsfWfjvZXUtAX7aIvLR/+lwcQW57UdRvBgC+lppWelU/H
HjIlXib9lSHHV8FNgVvWh7x4OUeHW6FcK0YVSagVIIYpSW30nlQsHGd6XL7RkJE3SF19W13n5asx
9eVmh1bfeynFWwQDArF1Z9pUXwUwNc0+ZYmRv8S2cfElYF/dr1Vp+XGohfNsdWLRph1PY8nHHPN1
IwgOsSPjCe2a5citxESBmCt2k04Q2v2ntL77NUbODWLls2TUmvpEOTwnenX3VVy+iPEnc8M55cC7
x64oO43F/Te0F7MGG+B1IJRX0nxqgznSZketMiwQVPV932vwP1auzcSm1dRdM5Z+zE8umP5scK+K
3AKiRn4Wec9nY+lxQwLyvXBvwsM3r9mpt/0BbVy9A28MfP3Adxy7aCgpX8r+dfcqaULo2C4fvpxH
e5MYJaFhdEgZBN/Xw/qImTFLWBRnVaD9N4ch3C6OwdFMgmAZSSlz2sdBVdn4CSqm7adQsg8jNgfP
1wdaGPSAfalBKJxYTAPsEHh6J+Vpgfe/vKOzvEWFg61sj7GAj2kKex2jVB5qHHcwygnXTTNEjJdm
RJKMhWp3J14p+r2aZYR2/+AeHkXcsWCrpv97bwkboKAaSAlZc7cneDLluRDsL4xeOAGpOfRTEjVb
0BdGc2rOpAAuVN7NSs/g1FmsN51fvoOHDYatCDFefK5iUHyVJlJERF6wUyqVsbHAyBhRQKl2pO2R
DimWJ6vjDRUr9ELKoqM/oDwYEIuZGo8v3ZOhTgsgjOuD5zp9vinHZJ/EDqX27+2x4E8kJo9nj9s6
JB2nS+EVzXduHPiCotF1XxIci6pNYP9G6PbR9Zf34l9vaYMrO84OZZORsmhPbwkRw6Fb37Cv+3oX
NRBgGqNE83n/1QGFq/CYQrcrFcmdYmL2ELf3ufLeYmWK2/TxDJ9ZwEENweHT3XeFgCSkVBriMwNv
ka05OD6f1GPt1saUaprkGbMFvmMrafttBAPIj62HZjs+b8ub8e28f+234Xa17PT2K47XQtKPIPg6
L9ejCQve3+030ttOOlL9iXs//A+qPxCB94RNGzIUfF2WU2354Uz5ivR1SADW8f1R5h4IENDeaTk4
WxYTSdJMxkxTjs1zr0ZECZczDrLsYY6HMVS2b6PXx1LjOIIp48wTHSwiH2YXS+Iefakt3K99GjEx
GyVUDJku2ldxKWuS+qMNfXaMZ9APtqHgNnK3IjpbLxegZRvv20lHwE1SdXx5AAs76/8/RN++XfYN
lbqmyOsOAhAdxCgNsDAXYbW6Ykv4a1vMoYAbFKPx7TmkJkSkez+i+UenafJLpIqGqmphM0o+ZllO
jkDju8E6yOJbb8z8MqGbw6uw5GERVilxHyBKqrPfjwu4JqPLHGB0V95KcXjlXZtxZJcBmLaVCE1g
0LUn5Yi9/wHXup5uAF1CNjuCjvYEGtFoEwtGq0C7oTtAk4K2xoiBWCQdZQHBpwKuVPwcSsrPRiRj
fUxs0OJuUrI7NvFNg+TNcFmhm1G22oMq/e0F1z55KOcrCw3DEkOxfsqEP53nauthW+n8uvKOWp7l
ATzQrpMZDTXIXlB1hDo8g0tsTXZgJmf1zwMX6puP8KJMgiWH1zRqiHrXbdI4OvIDcNHdZu3bhm2L
hy1L9EmOwcL+aFoEqIUVKbBbujRbJ0A2rOAlgDvU2PAWFco1NppqIpBFIYCZxsGfffZEo3Z1LD9P
ZoV33xZyRsvMiuc3ZMEuiE1SPspe0T52jFYah8ZwMqwaeoTWaRff4moBQoQW8vZyLPIRMx5w159q
JttyxPuN/dZGU+BkwyIr4hUQzKb+/p7KaE1SP/+6jXMeUhfgdQKtCdFfI7CZauAm5L7vS+D04Ao4
X1FxPZQSMUAVfIAYPtBH+lv+TIuDqQqgLgMC5F5Bb3VhIcOxIi1G9F27kX7Uq1sTKJpTZgYl3bP4
rnRaz7ifBydKqB5Cpr4FP8mFzaYfL8magg0ftuc3KDjs8xE0ezgfWsaeCPaMO3YVkHUlyKQgLnXJ
noiX1Ae4Ua6wVf0vTfDwcVLXvjuHeec4W/Yc0CZjm7urMYnL10js5aLQUuCBg/svwu8NDZi+AQ1C
3P+EjzIlvTpW1pjiQWVmpRPCh5HYlMRv9RiqOEgA0oJwb8oo8B0imByVXRdfFOcgZKQFQJa0BnJM
Lhe/4VL/p8GJPRgmIX0dnmo6J2ULSBH+0MjB+lPitoQLDb+vkiRJqmQNeCYLU2Q0X/tCcD7nvhcs
ztaYHQjZuKp97iNoaaXO84IQjFqNcYf9dxPTARHuk/gPERlyc+BYiLDKGDDWUYSj4NCrZVgsXaOX
dIRHSlgzo/8KPy7+xSjiVOx11cdLU7plTiwzwkH2MMifjiDFvy39kcpc055w8wOJNH/iTewtr+Ev
aEIxC3To8VAfzsrBy/vciHtVpeVidKUZVm6ggSXzaMvHdy64+VGCseieqJBMShnz9mGlHCf5Zljg
AksgHJkjU0U+OpVUVXYzR/zb5wXSUo6c197vK06yG5vU+E+OfAqyJ34uW2Yl2cpAsUyANLG1GxJC
xzFYq+MSoQiBZr7hKsiec5TSKbpyRPc80Yhrr9YCznsR+NmxGSoFB+W3vXXNy+tMjKYQn4lDiCbO
/KE/tybUFkPikcs731tCRthc3MjeO9IGCQqPFCS/FLfHU4hvDOUAFoJpLQACH1JRHb5zB/lWOCj5
p2iybNCzPI82+cdge1aIAyDRceID1JGXDelkUeN0zCBKnoAuTMr0IbNWeaooxxEKcPTn4Mg4LJje
TYma87pi8U4xxdJgzny5idGk2G9qp4FYzZ+3cHhUMSD14ijXA/nwxSQH/GLrg5FDi6TFe2OCCwgX
AN4sw6KUPliafbITIMpf8jTRhUkjZAX0DhQ3taxJnT9L7whLScNT7BIeCfraQDcIniTNOZM3rP5q
HJO96SpTLVkExu2c6dYH/a7m+SrOxdx1eqai/KaArQIet8Tp/lxH8D6pbqbJ84RcA7OdRvyIHOyf
n4pBLeX+IXbG+c+2Wokfh7OtqnSPG/MpC8JNIOeTryBcmn+o7QmBhWotInp7L+qoD0fpG7qspeVR
+EojTvFNzIjCmM8z2HvDmTd95ZRcDvbhVe2MxWR2jM9NpdGXi2Hz9bXAodJdqS9vImU903PGAubX
i61R2gQklG+KXl9DGbH0DJAJB8+R6j76jSVKDQ25+3/SaTSYoLIuAaDHVL7si3niBjhLevJzAKhU
I8DazXWG25wmlqBfCNVZwVwnzitM+NR2YTuPruYOo6MZUonKutJRDwQ1Ec9W5PE0DZADQO5/QfL+
qOwrlVKcIRsz5klikuBS+RDkccS3LAFpvZPgCXo3ErgKrjKKT7+pbQ8uZ3XzjnUExVzOS1Bm+9z9
HBTGE+zofepW6DJ8fvPLTt1vFHD4kDcoEeVe8n9wc6YsLKF0fufE7Z7sdPS1iC7tKO7MgTZWmAuZ
XwFjE++N2kmQ2bW0US2W8l0AaSZHc1oeqjSN6CsqA3baWwLAV6WHCBSpP7uqMHOtfqnar/HIuflJ
uXGjM33Df57Ux23HkKtEfZdBSuzQE6tlrnbqxeBfBwFnREVN+7dJVQwD46R/gQ0EpzYgVt0cOaqJ
7JHhruUmSWlPF7kQIdN3+7YGKlpmwPB9JfzdDyEbA6y/fsvcSUKD5dGWo6TGIeHMUWPW61pGWYNj
wx5CjvhfVyJSsg2J3/SWfbH02plWc9pGRUkShCIFMB41SdDA6TsMgBepdYfcmbzJMlY1G3iW3b6N
caOFZOneKgyDys9JcCY1m3HhPp28bJ2WhXBVAfGZul6orFXq9d0TjzP0P78OEqHGaC/DEeuEIFjI
1qiRmWsCJJ/ySJRQw3xvsV6tYp8fB5v+TfQ7iO8cCt10LoIgHwFcMOqmB5nZrRoYCQPbxMFSOHnR
pv8qnPC8TFXhcUbc6GjxEjVKGwGIntHqw5ZljChboRM+uzYYgt5wpT0AvgkgjOaaEvC6U9P9SGMQ
qjcMtksVmvNFKpHUw/QReplUK5lCOYr0YUGIqfa6WXzTWMFi/jf0D+rpHYJ5nGejf5I6mJeM7gAq
WzTLInSKlS+c3qk3lpTcEVu6O+8bxNzEO09aC29IZJGNINdxpiIe4lbi02jedpH82ajYYtAYeZxL
BdsWRJQBdpJ616/FGvEcjfIjJ39oxZN6MsZsgzM6myCTNWUEa8GCps0VNevqijzL1j0n51KORu+i
wf4DuDtd+c4Nw9CjWzaTDdBfvgaz6e6PgNY6KVFs4ywAzYpiHjkrWoa54xtG3NCWur1o/si4XlB/
nTL83g8jT1r99bG5yEsPpZyD+zuZV3nDY2JIzb52QKb1ryklwpX/bsz0UZE6H6YjxtfKrSWz+J/T
4GoIgT/YUGVfi+/NsS2IpjZMe0bN6aT6u2BKsLBj26KsA7tOn+gmrIZxsN9Q1FaGFtGgSHHnt6uf
9Oxs0qRq4shOnJtzjP+ExUG8+BTabGFxQvNUErgumidb1i71LuqIbDy9AqbTRyQ668u6ogGPQclA
4W6ArgCgWZCeyKaM913FEP7KZ6ZI/LGt2DJWHcy+3KKypJeoXRGh4A9JDmEo5SEk6OR2eS0qaque
QyeFnkaoKTn/kh9Zg5rrOr5ODKiair7PDIaSLKkh3MVlvIGY0/jpGgcoQ14U5aQgno5BAe7Be49P
dPV4pn2IINT4a7LgBXTVtCWi7ou93wSmwUomHTCq7VCwkyrPdhM1JX6E+Pu810EgwM2oU0kX+GY8
8iu0kcYNqxKSYH++e1ufy7z0AcvL/kHXZT06WLCoRxhh+HFTKruXMJev/xyrS30WcAL6aEMmHjIG
fOd1v9ZmtTy4hoMYfErSCxAFwM5T8NG7Ukz6IQ1va4mB64IipMNcIO32vM69lTaQieUVdufdyx41
nOP2W9EgTd7j004pV1MrF5uwIMimPSWge5Voe4bJa9JKXVPD29gyTKfNZ/LH+Mew9YnBlkE62hSg
H5uxYTN46XFGNh1JQBDU4Q1Wy6FjvCWTeEVDGBLTIxDhNBx7/SxusFW9DOUcM+62TwmRt5cW0qYj
ttQir6Z63VNkgZHsK/U0ZhiiqbB1XqXBqIBxxtokAMCfc3AxJ2TDD1RX3vPlopuruDBl/XABfK6H
06cEJVLYtP+XyOxm9tk8gpqulbrSy43qIxQUlhWrc7cFUekAU6TTu59kXAJd1sYzqIkHDESsdG4H
a8fjrfk/mIb8gnVrseQgowfUtySyBS524BXUc/VjGcMR2LiQhErCWpUsLi+HOS7qFVRze7fxTZzN
SwbsO4sB2f/PWYrEDf0eJ8aVwxTV81txOp6wfNgsPdb73jvcPt+YKYDPdaVe7hWgQafq0C7e4UNf
DbOg54wZgFygk2nxwnIhvGAw9jy8Tswk7buhZamKVzWq9GyZf6oJGd1Z5HbODPuLGDQsBL3AVeal
20+UsD5ape3AY8KJAiDVjZFZiS1XZC7icJCjjQfqOJOsjMZgO2vR5xn+Xd6KKsh0tZKKez668BeT
pIA2Z/MkXB+4tPIB37H3rEUiW/7w3KcX7cuu2tTmPEVnZgPQD6Y9PIn/OFA9iTDeh8jDVFyAY1va
hju3oVOrBBWIjYhXR/kDHHhQN3fatsXTpeC9oVGjoC9pL8++Q8M3+vnFq8DwZ7OyFJIuDN41p29j
T78Hckz1Kp52xeuBUKg2teyQuoPHaHrg0dDBzNG3B/Z+G7+uPH0EP0Ay25I8Zj1gtUcZTfXton4z
yWmxkU/Sm8SBsRwBiYATMgtbLsHyJWLT8gXro+gI6OU72LKOzoaazvAhuKLsunAEHcW4635EQL5M
HRCTCimhaO8kVuU6eNGLsS/+jGPbPW01c4T8dexvV3VO+hUuHgyCYtO+ovcQCUiGmYC7MDnb4l1L
CZb8i57Hf5eR9L47pnDLOdEwjBZ++kNhygs5haKkZxkSX4gpDBXL72olijtdiNXmd6tO4slnWj9S
yuQPMimBRS9f8Kzi4Lg0J9nl5C1yUq59Ko5U+YzsrxuuTxCqk4C20mZD1zdtDycGAyFpVMZ/LaM5
zKcvC1qfuG+QL/vf8GAW1HQZO61rczHlLUobBeOBO5km6ucFtFI1NhNSOad5+l82FnBAqbWh9VbY
5eN/MOM0PU44Pdad79hNa8PDzZOXgFO2Ff7mhQbQv1EdscKlU8zD7p0aeTh/7jFcK+S7ODR2AMRI
8j4+utb49i6v+jX/ZBp4msF28orZaJhnJeDdDbYJkDC5PAa9rqEhTM1W7xN/b3yQoy2zOaO0oY3y
C7QZxWV8cK6AAmHGzYpX1/AB3q8B2G+POYt3VFjLMLcyf0hP3N2gCNbkRLpWI2NrT5lqvo2ARZVy
BMLf9EESazOe/de+lX4VFKspVC90XQcwF0xqieHdqQq07AW0xW7w1tuD1flP63YsL3umf07dK93y
JoA3+6rdMBgBeuX8SyiVT6c88ntokOtgr4BP93jJFI3I1cRm7rl+tr84d4quOoXRcjeDO4tjphwN
8F5aNxscoigTROmRQ2SJxjsWkcuXlvU3KoZm2FD34QrWEVTZ4B2WEU0vlc+wpoK9FiNbqBJz6A0j
iHo33xjokrYgq3nkmeTSF7cGscwQeJ0aUTqI3HFGGmsdU/mfLFjMsoSA0Tqe7b+muUkC5N1OSuIa
0AYRtrgCsLAO/aR9bYPya7tbIdrJA03yebANViAFAJurR/f3vaHsKiOoAy7PglSVL/oPhLEknprl
RlA0NRnGyiVPUKkS2oka7AZx7MA305rSwLA7/39wbHKiV5pft7jodR9Vb7nytqAfQJvm6QfPCJ/C
vH5Jr/0PQmB8O3lUf6FXX85zpt92CEB+4nwPIV7TjulVVDfrDBSXUM1ySUrUCP99h9tp7i8Z4+zv
aVJjvZY3fel2HMfGpGDJhPAuRpv7mbIGY5YZTjcQbppBw6N3S37EaUycvKmukKrnqvCCDfmaZFKw
NUv9tFb7SMfIb7gP8RK5sXy7F+btjZiPVUd9mNtVd4Q6roOoI4YfJZxn915sfX5FI6aSYe9F6/NB
jr5mrxQe7bRaNQqpyWj2ZliSOZFWUdUBSVL3kxd9QgL171SSNXty0KEFmZc7b8etoOLMllCRFNru
xCG+vA+c8w8nIZTVjYySJnQNgLIXFM6QysQAeYySDvHnLGK8F7b/ooJFF1p2fW97hM/Tjcp+Fs8b
AmsJZnvDHixNShOPhlFnACpu4vlJpQKhZB0om/Z15AffyBk2YuFVQDxIKih7fRqE1C+o19M7kLWG
fSP61WokANdH/o3O+/A8iTqrJP8TLSTFbFAcegb1ksVCIF5LTBX3oQ9h7AlwQb8YV1bRTH/X4ULx
X+DQ7T8pdLOoctbxiK24iMsdJ90zcMT3Rc9WEQ1B4NCQXY0EEnWcF2Hj1iUQSoq65jP0ArkLgmOc
XfmPz4A9S3eXzdloe7yd7eb1UpRmfP3HOidVCaA+hVRzLIkQrqUg15xP86PvYVEnqBNyVMH1awFj
zDJWSo3RONv/0aeIrqijKJ9+72mxPIZ5221DSSSK0yvUphPbMYtGAB5UPf58/vNP+aEYRDz1JwZr
ewEY7R6lCKip0gtCSa/BzWKjGE57llJ2AZtErYgf2h3k2fIJjg+t8Q3UhkrX1rTUOT+Xp61o9DLa
OgxS+MG/l18Jd6ateM558fb8NRRDXFVIU4YfMnAoDJYCInFvzZl0vjlIAF5Gxiz7afSMPIPNdE9E
1P8vz5TV2+RcK79VQSqoC36aOYQXYwY7JolZ8MKTEYw5GD9y+PuYjkVlUsKQg3SQb3gcyDNxeLj4
4T1TgrVzaODnyD33c7DF6Lp6xZpqhGOdK0zpIKsQymZthjV72e6JOGE3APkGIHDh1jGcOBC+WUV6
0T+rhhHIukqkuccCOEm6MhFBf5GfOgEGp5vW+bmXo2/aMQacT3Y3REr1q8B06tTdZlnpq1XCf34s
ozdelWgkA6NwVC2ZZJLXVXS03D0YEG3Z/KuX1Df1tQsFSZBwJ8d5PXmSJn3aY6QZx8m086TYDoP0
Tj+7CcPEWt09Atjl1u5BjTtN3xue2Jx/NEmyHfkLatcxM38mZIIWIItJ+4YzQ2kLBNcLw1eZ7rt/
CDSc+77ksaJv/dlacLJ2NdF0870trqt5XvTbeU/4/lWP2APEw/qJLjuCPpwXI/PcJlRcWeRPJZSu
c30fglT0qf1toFgjNB7B966k321NagdMg+tJvpsEibY3UsclXCmyOwMg2VAHA5K3tcjTGSM2AiR3
k1+BrgkP9Be2pSg4vgdImUlsa1f8xpLJMjyoSNaurApdThssRQqGJYMvH40Jrnbhkw4w+WE752Xg
Vw0/PNpENop3usb8zifLpr24yRwSltGPT5FTOlDqCSnsN91TXaP+W3GERuYbzCJrNtLGxD7b4/xl
KUG5Cb1yzzQDxbS+xgkTnPtRezTFh+o7s81xUKJGJ4ONbQAv/MYJUIzyQjdRyC0P9F+E3bgbeYGA
Pe6akqLnRBTzBFCmb0Qups1/2SaFnDSf+yvUxM8ohE4BBfTUhmpRr+OWA0ZOgO1zSH/yfbvRFWnK
b18VPXoDviQxiPPFuJhVy9jjC49JTPquP0gA1Cv2ynitK1093TWlKMZ9sx0ao5fJDtFfmTpL+c1H
jEqfVCLghjY7AluZq9o7K1x5VrjcNB9RTss1xPeCeoJOAfGY7ip5w149eoyeX69O2EyrxREH8km1
CEarAc3JQ8JCwZbGE9OzxIdqDS1kteAzqFwXrUOeHC4vfCZFPOD8fqXy8LpplzdaQv63AwRQwxug
im2D+mN8K0b4DpoTBzP62uXKMdbNHs60TJ1P40fLYV3T9DglIYMUjM0GFxJMl/Bd8hPOUqfsioU6
tZVNiL4a+HhW3BMOvq4syUwyveSSxBDKA33c8AiXO4ZEABKykTsm8zYChZE/3HEnbwFUn+1LXa1t
tTAlXl8o/SSdZ8xMSOX9/ht3Kc/fBgbCVwlAfBFNct0MeBeg9Yc5AeGJf1GRLRpTdxKUzYz9opio
UEl+VtrmkvSzaZX+6lWO8gibgWHcFAzajnsU/4WZ0hMC5il+qD6/jifHMk6mVWsLuJgtJKBmk36P
F3tpIygek//XrjmbY5dSAK2oosX0eyCyAhVZLjixUYr2CpdVANf2VAPRKJMRCzslBBgMnyquyOr9
1DoKC5RTxQbdOOIk+5gr4ETE7Z+mmuYS9MAYSAcOBCxtl6gg4fYTTQHyBDfhxvaRghcsssUgmq3i
bZAsAijxySD5DOeFlgBsaYRBv0zHoyYYPUY5OHHDDiJwi4pcxNo7CGLvwssJt0iBkiFdkN9TTJko
HxnvSf9tn40PhpFvhATtm1wxyNllQRWw+Uc+miWi8QkPPJD3GYiMSAyJAyNk84i0hS3mN0I6fkKn
2aGTK0G1As056OIS2F4H8M/gDQbMaoLBA9CAndAew6UbNiqxbKbCdVKvA/QaJdII6KUSm1yigI74
LTGGjJf0ptcAlNK76trHdR1hWparKyxiugWZMXt1+g9mhX9s3ZusEIthlvWHSfqM4SXJgAEs+yFm
hUR04ttdVQGf2/nKqhAGGaf7feXt5Wf1xNxUc3Uq8NtHDtyEKOBa/xVF1gfg7XrpQ7KkggpO2O3Z
Sk1cjo3CoHgYhQ7gxachVECY2VDn9EsujAlHyujBbBkjyP/m0wPZj8CdJ91fBS0Kbhb9ioRWrLhl
7ORSwzER/fizTojA4ZrPVA7Ad6l4MY4FSAYNaE5tiRooOeliHL8G67Q5ZR+2pKLp8bbmAfQEHlZz
UBDSMQZg2HJjUY+w0asF58DY+3JkIdb6Zf8jsFq7PkO4XGOlVeWxDeNozLtMAc1y2mN4B2k0KBRO
UyolPMPhnFxdDZx8TXXGqfsiZUZ4DCzX1dCyOBrMoWktTpeXHdm0f01egt81V8Y47PASbzE76c4W
J2IMSJ3G/gi7mu5Yb1dp2RHBeBLPqKUQWchpkKDooW5bVXeGdq2G/E17XGUjXYOygLGYQquK4XCW
N9jjEbz3/KFj++R1BD0XmLK/MSGnB2C4b8NH5lgg7U+Hyw2OasUHAmJn2QzWibMalX/LeoCoe1ke
h3X4J0Nu20vCC3/MMGzRwdbLc34mguykQPX50U03yhj7PoBRhToHCD1xqthUX4mNoL2ByjJ0MaSi
M8PgHtH8jHziuCwI/v5sqMmT2sq6W2f2k5NZkFdN+ekyWmkmorfveH+iM6b0tJv4FAwbF/vnyYcN
JWsu5ANYqR31tlRZ1AmtSFnBAqoOVtGzl2cafPWyKWhy2e+7vEyZ5bSy5/VHIWeaVqIO4UanyUNb
5/TgVDqHfJC64s20/cNz6DfRNqvS/XtroMm1IJtVkbC6MBWHm01YG0CAnoCBcVzy/ppNJvp7Pp91
2mC1nW1k+fYjHvypYt3SjCjFxgTi+I0394FoaIW+VeV9oPjc9cepArTKEZW2SZMN8l6SRggwJc24
Ee2Nsy1zGR8xl6TqKsA7DGy95s7CvnWmhZbRfr64mkkbNELONQQyeapQePo9qVH1qYB6btafhBUp
YOXp8aeDMQLbP+I033SLtM47BYWHkmRJv5WuV/rDY140KvBCRy+aBXeFEFKbkc8ct4rloYXdy8Pq
fth/Ux8OoIAn99tgHQpQicXPO5szU8ioeQ4hiLZNQ5ioVk8tGLyTP9wgqNh+e56pQL3lO8g9kP89
wLlRlvN29k3sN4JStzaQ1LuUUeSuQZrIHs4FTGaGaUHQ6qDtgPtI4A1Xg7e326AGq7RrEk34o1XS
TCn76zAUAP/Ejrmvl8IiwU8hekhhf73c8OcDAMnTCtT/YcUcBHlzpDrXfrHccEdfLb4bbNyyC2Kc
EYGLoPh8wnprWl97RWvPelY7hK6P2Z1l7oDk3uMOr728yzwr5Kga5B78ROkwTRLodsEnL8EViIgn
1eVCu5OX3KeGwzQaSm9xljrpQt00Ropd0ziv9UucvhW8BOtr3+oaQtHzdfzn5+xsUuQSEob92eky
q1/CskAlrHJDGVPsgfltL8KT8vQOC+Fkweajdt/IipDJTOsslMdsqIjndXqpDTtFmqmW9/6wUMuH
gv3ZmU5Gjhb5fs0JVfVR1eC5SI7KnUCxfhAeq2lnXdghoM80Sto0MLo8SpL0+KM2GGvsxZ1YbECR
VkEhM7GQAGQVeYRL7Zs2kYpkuIp+7U4xgde8CedCmZ1BoT9rIQHNoV4A3JaUoCbL0y0j1ZQGEKdb
lhLcaP1biKP4x75UYsMMk86dMdV8FujThqDVSS467RICtnpWhNKaD+czrpESNNPtJ9dIH/zykrfR
IxdK3lA10cyyDN+3ELlltB4J/KsgNEB7Y4kfDBimX4ClqG9bPcHUR4LMId22abiooJIi7Ip8s68T
vYDFfkJW7Y5lh1eJ5ViJ/3IN3siBQGs9cJHeezF/IIqFyhETiCgo49URJIT+HNyFODtLcMD0LRgh
3yjsW3cuzccsXWNCUUubnAH1wjUkRAX4kvz/XWZvQX6qTYyEciNlE1fEQJJSgmWfl+Z5ZlF/9Xbf
5rc5EcP/vivA8vsYEkugvVuqVdrZfC8cLMQCCdf4s773qTmZp7bXXhZ/4SJfzr51hKey6H7MQoDd
jR/H1s+nL+x+5CNu6KeB9EXtUf9p7XtDJnUuus2EjUQ7f4BhL7BV4afQAp46lUdpSzffJoP1ZTDO
azcKGN/nyWe3QArpY6+yTTiwpa4Tksmv67HSjdCJzapMwpX8oY2dYuL9WZ7PsWXKNYJfUzjR2alE
ZAxP59YEeFfz4ch8QvmuxlRVd/sHCo8H1jnt2uIE2ciB6s2K2k5OJB4Sm7s1hXK1+Yv3rZSuzA13
l/3CtIbH/hTZmGcsAIYIMt+ggBhpeqbjHQrQXdEAuhJYJrPfTtJGa6dKb2VN91e99gA1rn0jl8qq
rIT6TQ+zgkevRiWMty8AX9vDfbVHdk8hEmF5YJ1F2kk9//G34bg2I1me7glbf2ty65G02/2b7tsE
gHC1cKDJO1n9AdRQUFsOiVQknC3gt1IbvbKCK+tYV2Ag3dkUH78Btd0YShj3D2UjkoIMtUEgAiTR
ICYINC5hmCmSUlk2iwi9Mjqk/Hv9vToGIM9TtQ7ZLAfqgkFBVJ0vveRlnVrj9NBtzUcbQMloHl/J
gkd6xrV3ZKObJpUWmSXHlbZCKKrh8u9fKbdahg1cUsvgY4YnaKIRaD85gZigqxRbzzbU0P32Q0Jz
+qerzfRm0QpSF/OEHEkFy7/KZFHf9dmVgklKFl9rQPaAxvwFtASvDAOgEeY7cx+Qe7DgCB3qzTHK
w03VDoXPcpykV29mza+gaGKE4Sf/2M6KNlMSO8sFNZzWf6kdbGEEAYV8gsdQ1GGJi846cvRVuqEg
EwFJjsUzAGiMn/z3OCJKv1WSgCAnNCrjNM8Ha9X5UpljsSnHKt92IRRVcxiYA5Zq8cHr0QWAudMu
f+NAmQJ8M/UFiKWTmS3Tk/OAJgtDCIVw6yH1FdwMHYe1kyHBNY+gIA8If6vnFAtYWCx5k7ZRMFkE
GR+uO12ST8ApxEqQqrBoke4a0T5l89vtN9S/7n25YvfUtNZ+IZBKW6S6JBW/6poCE2CL7BLjk18+
q5xzIZjyLoZJ7ALo432NGsIHPDKw1jXn5AfRrZNFs+UzGJt3h1Lo4Scm/Dc7JZDtVRPfz0xE3t4U
mt7tW2QgCghLmm4RNHjLn6UHCzulJmMIhRnTAoOEjTnvlIeXDVF5JdmppMGpTRhWo6qPV9t/lJVo
Vfn8wLCXDJ24Hnh77aKvpNh8yIUC5BlJJrezLW/UZPCoPmuxtBBIRv5k+GgBcs7Kqi2SQiEkgjr5
LtZKwTpF5vou0tssBR+GGjg9PHdcz+vgWy1UWyKnwho5ffZYnpEK4+kEES4mv6WUvlfHH6eWEjn6
z1vh1XdndoehDQ/4AskXd2cX9d9LpeIyMs3EcJr+TD5Cohp1cl3RmVyOjqmNGVSKd9wdm+d1bBRh
3DTP/9XwC6TuNA2P9cXaM6UtSh/+l75Fs4Doc3ZSo+EOqZaJsgRkEbhq4MlBbwv9NQmyHWg6KmnK
6x+u4AUdkFkdj94TZ3LW233wQqloguSndvWlmm3mYViqq/g4xRX8St+1Eja30eDjrESpAF+tFUrr
BueYpwaUVQFBiyGN3xZW25e4k2i8yFXpDZDubtEDJEtsEDqjgwle+Y/NeYp+iCSf0XmqQqs+ivp3
OI3ba7urlZWK3O7TOz2209XIKe317SvRZoL1SUhJRwtzD2dWeyTciF1oEg7wby5VIAUj7Dsvs0Hb
NxKaErRcdTXuW006+al2+Kf6F945IoBHt7Mz39ZNJJhgLhMVcz+aYher2GU/dSZQZgA/t8bIpREH
sAw6cGZDfP+W5X8EYLwPD1zN/VAJViMBKaEYDvCDepImpG42iGVFP6RLIic71Ds3uAMRXB8u0NnK
T274pUyO4mAxoEi+lUoaLFMMlQzM5dTdiyEg2NojsQSJNQOKkfywaVP7ldQSYUHmTaZ0qssLRBpM
VV+0sDZyvLOYyHmm5pi0qgWXLWmNTSN2N4M1N8ZFLYBzgcV99NB4amGSt5zuRiQp9HYgeVSMNjW0
WdEfvjavG3Ja1sXNAZLA8/dumZQ4X3FtXs/a5vrn43t3haVlHNlnZMc6cYysdm6RXSZOxSaHVvK7
c1fQq5bm72m870apCzM5eG3agIWUVT/MIVm0PnI1tXP6M/lzYbfgl7FNSqDmQWnKa91JkSeKbNUJ
quV0ilt15ZUjYO93p466++ZfzGsshmpjxFi8PYuDsOLHL2uboQqJz82VUzdwx06eHZVJHzYsJg+0
ILaOVfeIRpxpvT9GCERFmLWRa29rIWsj4ANXZHa1NMGLb9FryQysEqvM/ZQNy9N8VdcwZkZZMrH5
zkJMyrxWp55hFGRPksw0zvg/onkln44/hNu4sIj2qQJBceV/CPaQgAW7RpprKkKMiADlYi7bzVFi
BnKS2bxDfHQv8czKlL/e4ZIK4TicHI9vnWW1i5JExMBzBAWm4PYeSnNGpe9cph2b/UVCFUa7jpc9
zA1oFkSWh8l5KtzFc7wczotZGy6brGzeep7RqVhY+/qUn4zf03JQPXRxDcURZFppnRhZXEjGOnoB
Sr97Ow0aiuJF8X5X+9do7Gi8XPNms8hXzerHgeBgYcTZ35sedzM6slve73W1OXO4W16mKU+NA/2C
qc5wiIekcgZvnAllUXaIF6f3VNZXpXF7YhCpmZE8Vtmz0KwVX6HPe+Ot9oYktUhuW9viN4GqbdaL
ao/GJbfhi9eBRJ6zuUGQl/YFNl6XPvYYdI5udH1ZSRPvns93CxRPmFXDZGxEjLKyUSlv7eUbzQFf
oXM8Z1kh7qVFimMqV35AKBrCM6ZPqc4lQ+cfGjLWPmuFMxZbu3zKJvapyMYiHBLnK6B7c+7oSGt9
t73FZ5iKHvxFHCWL7bb3Cskp7hBNWvxWkLvhzPFX8BQPy39h/6xqgexLD5YJ71s18iM5iBV3MZhf
YjgXkCnhwR2R8xub/RUuhWpX3yOcmzKuS18shLAOpAM7jlB1ppW7iZ1fV6rBD6W4eiiTXlvJkKmq
dX8mk2tKs+GqTnvDDTpkG/GfhaCbMEk0uAKhmCKUDnRryELe/jBwSkGaiCN0LADt+M+0wvZbufwn
sFbw86Kmt4dE+XTEZvYis1ZgiWmhacFudXfKinE4fu6YJCyjpitjnELUFYjWv7YI4+TqM3mw9b71
Wldt2bw+ca59ZGN2QtjtNnCMq+2ACIPW9Aeae0xFi4mDpMB7I6Z5eU3R/xlKQpFiZrgZbFRJmDYh
zf5I4Hln6Y6WdsByYoq2cf7/V7QwHOUqwq3C4HxP2G98YEG2xFKS9r5mmE98ruro60rTgR8i16R3
kjWh6MOR0J+gqRtscvWIk06kW0URFIKFrHlFL7aGcKa/Qe0rJjSHHJ2m2z/v4PNq5zvM3n3oJgrd
29mZyiHaShl27nBikrfpjG0ckrMnMnWPevEIJswwRIqs27ZGzvcI5eVqSlvJtoBGI8uBFlUXXsSv
uX19Bo56YxVsvnf8kX2geMeu29eWW8wokkIsMN9R4wvsgMh2u0UbAi0YCoQpjh7HW5SjuaO/PARM
0SjR4CpsnlMEZN8tkij9Y4rW1P8o+b5zQHFeq4yKim0B0n2IlswkkfBewCh9KLVq45ovs5lAZRsL
v73YiaKcN5Adg4uNVKUH2YXTJrAstahVPjbG4HrAfIv7Wz7LKrBNyz4zhZLeznBK2mZcIvqPfs4e
KjigkPoXhmt72HRbG0Hg3MUgO0cUJOu3jgkF7yseQPRdZw7q9wwF9pBTGnP/n3x4Q+Nj35sFIJwE
t2eKSu0pJCkNuorKENF45Pi+AZi9D5c7FeLdN0bK3M3BXFdTPxsyZc48xNR2V5dhHKYgjJ5E2nVh
uz9H1+TKf6u/fDnnMs0Chz3izwFhnTg7AXgBMbZu8x+wvc2lCQ+S+5qa/4tqE1vVh32CPTllXcow
AEhP/zZREUed/8Bpi1pNolQPlAhKDtF8ULUPe/SoE0Am5rIRxjouVgQU3503GOGK2aKeKS0mltnT
AlWeIit+NRMn+sEcC2/3vWuk7pXXmR2QXfihpsokbcBGIzGVjJFKak/qdKONgdpRqH3+vvWFg/0p
7+MkFPwhULXZyOiUvD7dWm9lxD19MoEVzHYMCU5Kz+1+5LviIDLO7zbYoa6LDVCMIy3t8Cqn7Cfl
MHIuvorWUCBuI14XC3iNFhW03BBW82tzc6wgvhvBcOR2jSqFUtC1Pmwg34pp4iHS3EE2FU127mIu
ATICbKTyPZvM7pxzTWamYDC3JFpkCrLXZ29PowzjclNU3cY4/cWnanBRxbwuiGTU2G2vFHZ1K0yF
uIyl9T3QdDOfWprz5GCQIqmjwK8gXC54ygWwgyiK3GySNza5vhFwp5J7txMqdt+zMRLWwAroBXvw
vk10oYjxObGv8Kb+S6JLoH4L5sHObEFl58dKgHz1cUoqeqXOEvgbxX9pfPW26ihPaDoXvMyB8PTQ
X1uMa96iooTc+7fRsv5JvzQmVomHWenaf9RhJ1zv1W/lIirRo+Wm35WeHiJVA3O0k7tIw4mNe6Bd
QQ0TZlBoN04FAsymifR52gdHxupoQxREKaZHNqxsDy/WklljSX68BuTXez4n7FZ2CLV40uxshBkI
12W3rHNni2GTvWHohccwM5BoHSpbq7f3qQ7WQN5qkallEJF+xqMKZvP/v8owv9pu/EZvCVOayQ0t
kQcBGwdfW43HWPG4D+cInyWR7qQ/KZ/kWHO3FW3QvDUjUUxkHyOO//BuJwg6ATOTNDmHkt8D5o3J
hPFCDuuaooDgJUy3iLMOv/yXxwz7aD8tOVJ7zMsmryAxPr2gCnZfBeYSBFCk47/wvMWP30fa/p+F
erJb89o/PHV19MFUvzTjVBTwXBMohze5glQAreaxoL4xYzu0qu0ek9Ab3ab0BbkKIIr0lfMXZksZ
1yKVswQafCXiwxZNC/b5zYroIV0NeHhcx35FxMgnLWpLM6rK7JdGJmHSU3AI0Ip9yrlVsdnZFNEy
ADeiSYHu0QkD8MRO2UX0qaV+o8W8K2hR9sgZETm8HiljlksaVM1KWrmLCMPjX8GXUe+dnQbZDohe
4zJymqi1BN8hgnYH1bmT5mmdq29lG3u++AqgH5WNdBfrW4rV6+32iwwLJke1TfcdRKZhF4TEpr7v
RMWLC0SxSKbVNyy+/7gTnXVXZl+PJ2fLCFe7mCCr98pUs0VheweUHVM6Pk8hnzYKK4XmfYcRVrQ4
AwPpXVzlUMgf2xaGYc4S/0ZSGLQN2z6lYBub0gbMHLXtIZvqEu3qqcvQO8y5BM8of54Z95UvUCUW
If1YmJtFFyjTY3RaZ/F1LqGNgx+JWcJoVKiRhkOZO3X7tBz5VtNWwFKkuw89Q2uK5gfEGWOYL72H
fIqIxe915U+w/GvkwGm5oXod3QkYbGvpjRalb3ECYE433BRw++8BxC9A766EUb3Wxt/sH4az4GFH
ndl23dgDZ2qsXudlDJ7VseMQIu7hWg/cuyh604bdqxUt63K9pR86o7qOMyXy44IIEtuwxh5+bkG1
P/BIjc5b0a50iXI4TIpUSEECCMU0a8PsoFhE070cZ2oyV0ArPlxUqc2s+aS7ChFcOYD5YrwA+Ifq
B085FZPmx0+vBV2rlIdegwpU0xo/p2VfHDEDYHfxyjjontRQLk9Ts5us+/mVqkc6ViwcEnWgxzjQ
fd0B3oJopONSqTzFo6zUPpH7iUwPc8r4vlyfrpLxEE4wyr7od94xoS1KmwEExaEQO8rD4z9OfR1g
q7qwR83TJrOGyRSE19VqydRi8D3K+Suaq410gIx9ukh4Y4QDTw6HdhWKnck1KVhlyMq//QS5XA8y
2m5IChKN9ozzqqdeq2GCfqHQPBaEVrT9T28t31Z5FRyj/GX75ss4PHkTtIp0oSJ7wMUyed54CSYg
hbwCEJzdJ9CBppaBn9LJ8RkJFfUOAFNofW+hXnxS40xfy8iqvypd0eH7mnnbdjPvN/L61CAaRq7S
/5vTjz/H2sLXqb4xA8uXji+ZqQ9iWwiDoOamC3qHVpw5Jhpv5w2vcqZoHxWxgRH3dEu/OXmcipNl
w2Z9Xl2/qoz6UapDOH61aGa72wV0fmgw2q5uBK6EwFyAixGHxKI1wlR+yWTLaQWtRt0ZW/neRz5w
QkIPJA8l2xzuTcvHGpRv1M415ebPiocSLLtMncPpgABeUXkD31uFgG0c8PMA/Q7EccDtaEItTWYi
IvMrLEql1BejIg/ZdpgPp2LI+7qOyI/RLjkm3qcYskG5KNibdQUT1u+culyK4d9ySFOgax1/mNBt
EmSnG7L02A7sF8BG1PdlhM1iCGN0TBKf33EdKWrRpGxP2OILwp2JVeMTDGVyw0LGUWAdMoCoz/3N
w/Z/g3NgJSf2oFBUij+yJxSHhCnYthyPxl6hrXAmN15sX9ZF8bPGAjyPdxpvq1p+0EH12+wMmPiF
wEefmEYQELnu0ddmXrBPsEThJQbE1JjyfeKg8Zx0DjbVRfrx6+QLYbpHvE2MRmBmBwwgTb9p5mC2
jc/Cjyq7h+mfNWVLtCbKERyTMfT7bKDrMxuUs/SwWJAyz6Abp31rd9JZxv4gAZ/kfrX7v53u8Uvf
Zz6r5HWs/5tg4ybroPgMtrexMZnqwY5V6Pajd2er3YvyDa5EzGt5NpbnFbrtwsrnnZaMMzZ6ljNh
NicjsBowYaWrgo3qr7re7vZJn9p3ZZ/KxursitQac/qbE/msZdoO8wNHvvTCDE4OcpJtCuLiVKkE
tkJ9IEm6GUN6M0fdVgm8UvsOre3bSuX2Afol15ad3+3L8xsakgnK1Y4y74wifHC+PyDEVDhwzjPS
pyczGmkrPnWmK57VctNt0VlP0kXlhIAUb8X0AGENkxCTvaHSi5OO28hVSPhCLz7/bPwAAyGm8GMf
Cf/U4DIjOie5ak3UxxPmSf6m9jwOeIPe+SD47+M0RYHo33Gr5GQxVhrh2Ys2kCIBfYLwVQGVptwi
2KbwoqGXY1m/HuErph5L26zOyJGE++oLdGH/FOu+FvyxQhfzztmh5OzYk9GI4gH5Zx6YqHe2Gfsc
HLPQg/od7KmAeGuJx89cjpbNzeM4wNpav39FnrCWIoquUY2+s9kjVQ7SG5MdKwXghqOx+5+5TyjW
3ApiV65YZV6ucix1VQqJo+WTpAnmpMQYHf8ruhhdVuE7OseDGFmaFx+JQQG3Jg+o3HdD608ZLKo/
izbJADOCIiXSgWMdaoRPw63942qPOpKofrbutux5leN/AHR8Wu5xiNyfVCCWZn/h/VUuuxSAL2LK
gXGloABNKVFwKDXDx6DCOrGQqnzYe/2wGRgGwL3IAWjpkcdBR62WFmz7Fs2FCyjoa86q7OSeK98A
bVO/HRAuQU+7WHy3YqY13Z0fqpfysE1iUK01x53EAHjxvb16txyNtgaz1nFFnoUqmKDzZIi2SLQk
FdJBau7h9ooLas/vD0qm05EMnSrqtXv1oygst7Y8daD7C0T8/Xx6qUJFvNRlNoyPB8/i/PUWMmnX
vDpZdUtAZJMDJWXkgxFeHa3PsudQrDTn41DerC+0KO267kO4N9J70mTfnaX7JPnbgMhUlTDwW45/
KvGL0mqwu+ViNJTnaM8bpfRc8XomJgjt0d09Gi3Tr648vyCRiqpOTpXLK9OL0Am/7ijFEVu0626d
6ctHgr7+umhhvKQmRiFJn+lk4/5Z7he4cZhBDs52t4hQXrLMzQdRlINKMwFdMhPQpcbTxnXyWsAU
yaev53q/9HeuWwl3mjhkzumMn9p4tap4gdZ5EHBHGaQDEw5IpAPE+b6Y5zHK+9b8Siq32m+0De4d
l0SbfcUuNPvrumaYj26u6u+IHLiexeiLGdRhb/1IDZI87s2l7bwt0ISldiDKVEKp8yDRyjB2/QFV
3daUuzt6uVGzkLqAu6/1I4g9rJT1nRbWaTp8sTItuGtRSIvT7IuhuyMnK+LUdsNf6e/zOxmVfEZs
oJC6E9Y5FE5AZxGeWMt+7YUnqxApwSbCjyV2uZad1dULCAaBnY+lHjlCRhluriihNZ4RxdmzEclF
ZaATpRl1x74yKLhLqYmh6Uz71mhGmFoy6ZFTihVSfX3BX4qpo0iT3acmOgsFxfI94Yjnl9e4fDyB
FiDSLnBBePhWkqgfbEuO1LT7nHDrpkO5H2/xS9bJXNC41tdJzTkdKKDy8VbAg60TwtMr4cS3vlI0
sux5p4aOMjWcH9FksVn69SHpz3v8ZMUyho9kLtM4ry9WOeEcdxod2XoaVXh4ydnihMg5MFRL0jSE
7Rp/Df7bbVk7sQI76a7jrC+LZF2XcIRe/DeJuiv68LIDDDkRljXKelep3wloxwHd35ErofuU5Kgc
Cy0bt1hzDgj4B/wSQtXkR27f5y35iwNW+Plc8MeAVca5LvAEV4IlD8WMSwiSI1bSVacMTzrx5pRg
JGq4OZYI8QgL7Yo4L+EB549S07vHmMtkIFebOebBY59+A+l8WVn012z1yM1pf5i/t4wf1xf6RPH3
aYRHwOmLBTUB3rTVU4VoNKntOl6Hs6dHrYfJpcxtEHWdJMB+QWTHJ8Cg1fiQlGwQKXhjwnidjN/E
qZG5R+HLQ5sAQ+rmBIFl+lkUr4DqWDWAmgN4oNfvG5/MZ1KXHqd26YgDIV3VGEZQ/SLkYDQzoMXo
d6jW37YWYiOzTnGyP+EfnjBFE1PDua/i6r3brcla7Mg3Ioi8JFOugZKecPmSnGsMaqBcVBgBRZhh
BBx9WT29c7sw/NKDHX1CnhuTgZfMD2ffV+/fpGXc6zKgaQsOUdNko94wJ2VaqCF4vJxvWJKuuFpF
uezPUN+n6WkH80nsRliSiCxD5qCneBKsDnWdWEpMs5Bwco7mrv0vSmc7LrWwUJSSzIjCbBwJkG6G
7wh/UKVB23H4Nk2eOzhSOzRGfsukpEzSussUY4b7RHVZEdIrVeQW472hz6Bf0zH4CmJxIHTyxxq6
BR9BCF+jceMu3NSU45J5XbBdkGr4VZUMqMGcMav4yn9SvSxiYqDbMLIalJ9fFzek3DgNn4fz7TTY
6PTdUt8etp+qGStaZGcaBL2jc4kjN1iZrkJFpjOMl4n5JUXpkHpCoO/joc6mUrpy+4eZtKSD1wTW
TXkxa+AKIpyk/yIvvs5HhgXBvuNu8pTSFgPUztqIHS0/yiYBEzDsOPARijPQADhNo6O4qicZEgRI
i69YM7uZCDRdiwz+ia41FfDGj7NAg+fec0X/eOzc7CSGuu3s0LmBWi4LG+zpTxt+o6J1sUQWI1tO
rR7f09D1bQ+C4hEyZs5VfALo/NLhTcxue0r1vjOiGWHk8q3wwNJhcB1ImMC2J0YzVyCLT13JjxyF
F+IYbm3P+m6wEd8+cRQo5PDRGlL5j5ZGF0ANkJZ7DaJ8sgZ6EONLdTFv3DxjyJ0VCjD9kl8+uM0I
6oAn17CQty2HqtmZAuFV9giki+yBWmeGGgcvu5doVwYnIWFRVkYvvXctEsKTBYGE57WLEMNjLDhK
QYbtWWnDxVtluBbhWbM7uPYjCnXPGVkFJjjlyJT+ZItClzoNLkdWYnR4YPr8BqVx7PrSunpaGBwi
xsA3CzWTP62+6G38SYkFB6tFlCoGkOPQUS0oznuEZ7CagiG/6XMEd60Los2+KOMLaAPb3igrEV1S
saSo6V5hh8hwSCVrkZsqtc8XCFnNlH9Uh+f/DEeFfd6kAH/26XV6CwfpJ6W89DEzJXG0RHLixYge
YTkI7Kn4EUlybJsLFW2vYR+BX6RbbW6rkvIfaRfIYFSzaBTnjmHkksXP5JJTWcMWuMsz/3fSqH6c
CO21eYcfy9hz2jacCS7+FbfKrhQHLqbBdv/+pAP4d8QDpX+vcoWb5cadwUqsxqzl62lluUtigkzP
4Wj92pLsmug4VCdaixzhAnMAauiAIxvyHZIDmxnGMzT57Wb1HaCPXuf1fqEiwHW8AHORKLiB3CEA
E4mhKiFeW9clSC4BAOeK9/L5cximH0lk5NKq2mgYyMueEH4+3X0ZCv2M9Pahau3cf+YlqF82ajE5
kfQ4Xrder3I3IDHy09ML9tuNHq9ysNrLW452TbQCgAPhg014o7dFUJZHSYEzRuzUXint2lSFQgWs
aLhbv+N9qrTDwYenTM+qT1Yt/Bo8noXrxPyIEGT8Cq+jZQ/6FXYzT8AZQCJVCNwGFX5+ljIIXLrf
CjITas2sXv3gqRh8OBQZSMf2ZFkedtvOXwq0AjoEsW784yEX4D3u8equ8kldBwLiLXOVsYpuA9uo
kKOmzFe+0TJzTU7MjTqkcVh4dDCct1nLwlSkhEu/pAH9U3FJmCTenpTwcJ8ALhwDNw4eDljhjOny
h0xMqPIRkYw248fP7DiL2YLouQx8070gmgz6jtG8emDuQwYGT8ha4bRrgr+QlLodVWDYs4fCIYmI
YKRhWunAj6HoH/LXZ9fCCNs1wwGzatIHHfA+B6+HHwIR+wwPpQbWY4AfmQEOG4gSlfF9Vk3Rh1yB
GF7Bi7UWTZRx07LcmLrt6PTP3+uGcPPHPKyzrwQHNglqhlO7FdkmJWRkdvZ4CjESxFWtOW4rTMV2
/gE73ZQMXVvVD87UMO56GmZE5XY5hGG6iAdEY9TH1fIdRhog0P8vP+feU6mPWfgqqWJ6tlTlscRZ
B2guPXxGflmV7gCSIL0UCFLJodUv7Z7TIYMk8Flo16ir8jC5C9c73GszP1JgG+VWGrieVER3trFG
4G7nJxzSBWaX6pbx6nyPjwgM8mYcTissDPS5seWTWObeM1BWAOPMZB0vUDEKHr0GqHoz/r4nO4wp
EZ29RVB7sExnhoCVwyk1C8GYqtWt+Q+KNc32HS1MTxJ5PmzRnvrmnXeDg3Ag9rvBp2BnoeT6FHel
7ANQvHk6/jfYGEv6AR2jLcDVqqGNhqPsEFKoGoZgGirnILKawqRBV9p9JgP0hJPjooc/KzaZfXCx
ZcfoGEJTpi7T4XsajbQ/CBPkIRE4LiYdOn5budwcP4OJSVsLIHHQgV8oJ3x9kgJCH22eUs+qw1Ud
m5Eifobk0Z0qpNcAVvDx+h5x+U2UwFdIQq1htv2+HEkw4/9k6aTBbN34zVP7OqcEXBbuD1wPeXBl
LxSqR28DO0dhtP9ntfBBy2Zid98HvXJ3iTuw1Kzx8T3TYyefWSEViheDxEjteiDE6NwaHWMJF45L
wcYP/WCQBZL/SbsgdX0rec6nxv+9Kihbysh5jdAEetgnQiE/G7zCN05o5WyitZmr5J2nRtNWeReT
SS9QbEn2Akqr9qNkEeNjwFbOL1MVvEJu4x1hI+BuvrzSNahpBsJGKX8nYmO7XZp/kaLKrXPQu3B0
+W9CRPSXDRCFuej+BTIwWVht5te3rRv+E3bgLAZkwUvSRaEbzCSq9OjpP7kW2KMISM2WjN70bTDJ
RSW6b1UrSkOqq/kx5LJiULHUFCSeYRBfBy1Lqob0koe2a15SLNVZ/hnNahRGoLRf5hruWUAVXK7Z
B97ZkAks3XtvMw2AvOvYFNcVp5fefmRwsradS7l3AxMNUwgq7Ev0ekmQKNFD9QO7DNhLTPMyqcqa
FJiryydHTkfejvzn7vmO7ttRIkgl+eVziF543Q34QiOXACvJBwMoCZeZKf7HpE3oS2Oh22INyOJG
h2O9rAS9NByjykzzMXS9RZcPoS9AmJH7Fl3OvlOL1x0Ug81cORgJjKNgoBFaOXppg7PaGvFLkCU0
g57t0vjoeUAHPOO+IvexN0khS9fZhPGgl1pXClSCEMGiH9qAxdp4HSbqciBcUP9DEAypXqUA2HPH
NuKWBHDJhF53Ocdu81UyAD9EMIeMuVAhQqZg38X7iLrkczI1Fw2jhUgNADXrG1GwV4LD4BJkq5WS
+O14Obz6sBXGErJqjJrcuwLjt4mjYzdH1LP/1DTby+dRaEK1OUTMFLWJYw/Okmsl6SP/CfHIENUh
Fszr56FGoCLinRxN2QCUHiIw6U5EvTcq5BW6TUwpj1GI5WIR68KEVkhkd9Lz8ZDm4iHpna/H83k+
pIcji6a7MzjI4uMsiGPJ7gIwEtfwBTmlWbdy8Axl4f+WXL5YINKtBgoYQ+8Kt/jJIhu1RNBIg4Zi
BBPc5rssEfCPD8FKu9uiwzhDHKEThRVXUfmOCVABKu/HO1jzpWW3AbM8kjcHQY5zDLScWWZ17RDK
rBR1C+q5i8zuOsoMrCp2FT5motJAEd34vnFCYfOHxFG8KiDVYIo7IhsPq2Bk/yfAaa+Ev7Dq+oDi
WR7m6DLFPNOih84bpbyurvPP7H6rS8TsmTT6fgP8WhUfhVmHnM71tQJ0vr3ZrMTMu5i7dBABK2vK
/MGHQBUz+XlfUt2YPvymzc8ZoGYdFWvKPOBVqW5ADTef98iAd5l4ZJ6sCdwS80/P2s3zhlk+jovK
jvEmOODHJ6Ttb0CbfNhZMHo9UZ9/4hN4nTSexVrZIrrkgX7xc57lQoBZTwXwy0ImQx0dBXZ/mhEq
pHo7pB0uC5fxA7R+KWa7B4irzXvE+Z9+bos4mPEFHbFqFLRs3auE80Ia1+IRajr44eJYd+l2rITB
1lQAHG0FtZAjPecg1mXAwl3G5KewsgNFqJ1d48F4Z0T8qKDJ/KaNdKV/AB+GC7u/JMMnDadthnUL
gUY5KDONv2kGrgNBYY6YcW9TsbliNrTVqQda/wlNNxJHq/ame+lmt/+hyiNMCU/NVqITRPffLl1R
/NxMwE1Vd6qSu6U9S2ETCdvYJI8wdMvXi6dNop2jQvZrT2JzkjxMM2FejalUAyGRzYJn0PByHFde
7s+Rhp7vfEdzo7xPwhmvixJnbgEoydBL8ABiYScgpK0PnPIN0+q55JA3QZx6VMk+TLdnQXpacPhq
rwRo4VAJft/KvpCExAX8IBO3Subrk/8FufJiKXfpTEJKCZqtgbTTAlmlTuZ3KiHFIUnES1Qmct8R
lF5UyzLJgXC+kb/7dV57an+6ACmzKL3VNPN+NPMFLtnJ1SYtCthjFh6rHgOcXglDUwgSkRiUfHl3
7kZh2pITLDSnMnnJp+EeV3UVG4qZNwetmmTQabxRJU0ru8KrRF0vKvZYGy//Pkj97pAwMeeqIR+r
+UXvKdMDnXDXx8aDMwxWakgW3VVfZDkMl5pAK5kTZ64CfWJh3ZgdA5ucBVA527KKbbQj0Zg3XCqY
MgDbD3rZn0RfpBqsWWBhEPkBQVWUrCbFNMo5rEl+vEDiXEOYWuN8Vn2NciI4rrAdv/MIIQLIa8wd
bLUWTql9VCfU77uVSmFBHwcHT0PXaq3zBiMJGFgXc0EcVS6EAepEkDj17u0nFw6OrhdLJodKlP0s
DTUU13qBkxDazeLTIVYP5Y9bkXq0LSWe4AfjfxNs46mXY9NiTiKj41IJKHTQhu2DjTra7uE2Jlnz
2eOu8g5JS2u+cuZEbUtLqX4fIPQqOzIzweQE6LSkdv8NG8Ul6iTDzZCGO/8nLKth0Glmf1EYVkqK
oA3EGrCO1MZVa37SQNrOXKCA1xu5zMk5TrGbubmLgjsHK4hs966hJqksy/dwjUYvFM8SdMfi+1GF
HPJiovhAqRKAvTsXj913PyQjsY6/GgDqyhUeJLs7Cgmnl50GrlQHPCsD5AOB+sispJ33puwlt8f/
d37uMjSiBA19oAMg34YGZ3o+uea8yDWyFnQBx7OeV6ptQYD97mg+/hW+LS8uA+co8FVePKNIBZqE
ofmvQoR9BqmLU4BeAgM8FxwOUIkJyXX7LH9lsHO4griSUxbDI+MbyazTCRMoGgMzOWcnAQ9hEjaj
0KDZm3meHiI/EGk0jxbxSEndomqVB+YGhy6SYbyFDo1mjS9nMV+bDB0gikIDsRmODwTWFVdHZS47
AG5kd6/Yb9aG2a3do66594H1yl79yANuvQXECCpmcnon1gS+vKv+4og7uy4UofCqnZdhAOEZXwiT
9fEFy2v4ZmVhiGB4XZIIq9eqgFZwu3pFQo+SFqy8k9MYUIDA09Tu2FtM6ZBqRsstmg9GjQFelWbH
G9miinSacB9kSKM7jH8ycJdkG1+C3f/QMsHifagD9rZJn6FMnNhd2jOK7v30s4KabSPsYkeHN1lb
D6KDgCC4Isf9BiYTuklUajRaWa0Im/c9hfby35Mh8MD+uJT3lxxMf3ZgAmxhRC3WH8EjZZSI28E6
pY9uAn0Y9W8ZnyJyjEBNFwF7EIRfdOOORvof5vfIVVhZ6OXLFW0Ys9Qg6bnK7YfLAMqV/d6ULHL2
AaYlrXBgqzrsQNQmAK0MZCHOLqFsu1Z6Et8wa0WqtG/T3gC5EX3FoWUDlrSfYfD2dno3Qdltn/Nw
4+UnCOcZfEupjuDYj312Eq2UIju61PehADBlrenvRkjO2/foqeRe09PCPiK+57mGfCeyIY6VJmEl
2OnoVE62A1hSRUjOePqL13Hz+F2xkhjyDiZ/p9nbNeOiUVQl7aENf6Ye4zPkXxVJDY/WJZrmYbEK
OmEFenZJU3Ycvq9z+hqLv8YeUaO33WP+8dEHRPgSQUaSbWJgx5ImuyF1zd0Lu7tLpkF8g1TxvuSH
re6tWj0Mf+uetGUFJn1mGGnrZBQ8Cj31V9e1fPQAh1PkOo+XDHnW8EJlD1SUK/S3OdajNzkrbDSR
C1BWq6H1imzXzeS9T6DDZe6vSyQ4VNp0DkU22V9v9z+qEhYj93UNUh9KhznrVWT4pYwksN+W4ql/
06Eb8tM8E0OrVWaW76YPFhh/t7StaAY2Xd1uQR1oMpRpEJIbPmoCt8wubqr6HVGeoaPPyi4pUY5S
ovoVZ6t5XRSplLoPgM2aVfnSpzo2C2wsVYrizDcngCHbbytaw6hvczA21EwC7/7pfMTA3wEYzkaL
mraZRjJ6ppZrTJcB0nju8fLni8BE3HBgKUi1uRouAplBtEswEb0vWsxdycEQyVaNYyslvoGs4Ner
cTBv6FRxylDbHI/CWntOpGfiyEtBm0Z1SG+H7HgMSkuo+o89p4wjLYyaq+kunFK8b5K1lfh92rK4
11ihGJf3JMZy2WucIsQb035XOded6y9PtATa3mO+ImW8U1wbgJT3WB+kl2R0G3mMk0iSQF2WXS56
fDJ0YHiK7J7XjGVD3QyfZrkRWpyL5y8EQKW5xxRmMR5AWNgCSd6VIGm50/p88qtjHj/qNVO6ytQ1
4Ec0hlkzPXr2aZKVqG5O5BdxzyVcm9vu/8wwU3jkbxReOBPx4UBFN4/xfoGhh6a47XERPpX1GiEN
3IQfyxY/Npph/7yoe9KAr+eHGDzmNuhvw0RtTkdkj4sxNiEpeTfftEDlrfAwAiN6Zf3Hko3tjlH+
J2sMq3mb0aQZr53E6c68hzS2jrKcXOi6L5l6Q8o1+3/kz0YoBTy7bXOHOvEM746UBGc0O1Nv4M+8
CyL4ucs2H14aDeyxwFVjArKKjZt7P4pRyQmOrjvRWA+UygQYrLEUALHw3GpwgK7Vd1S/nLRxlixG
FygyOYBaQcsJVqHwLHxh2Qr/AP6Kn3QBH845TsxkrDYu6xaBpbWWSchJZLLru1csvSyZn/5kyfgB
HThZ7Iq+Ss0Wr/SvmyULiNALLbkPEbeii28dVkiO54Zb+sjPIC9pTb8SJ4/KyTKyWMUb4wW2eAFv
r9hxUKzxjgRYM4oJgsDqS0pCSD3jI1a6nGt6Rjfj0H14iIMhJD5uqIWNf+rtrQdmJfv6yOaYjbLd
a75iXv/hjwDUhXGWXvDDGzD3ndSoNURQ4LYYl+OR7yFS2IVF5FAh/9gfqR6rkm20JZI3eRmu4rPE
xsIP5/WbHhR7qJgXDlk483Luz80P6ZtRsRHRhbt1Y6WOnKSvzWLiRdv6QPmN7fcoeZAN2Y5eqKCp
JfBn0qWCUx6HyDcc/4ovmgJNSVm3pT8kHrtLrVvzTCbtYHj39Y+KJDCAuWU/0u3mYme4JCQkh9oK
KOLOZEU5/nNobAK1Cf6ez4NQXZ4wTY+yZ4c/UQm6hbdS3MijCNybVbFLUcdlHcaKDwsHMVVhZgPs
x13e9i3mL1fg6nJbFypJVMAkaug89/lCDfX1G1eo5uIqN/lSfwjdkwLfc9bfwn+l1DfdPd3mnOxj
vZdv6TZ+JducMUU+116K5DO5q9ROwKhvXb2EeHu8oZrfiaVxbNaIp+Si6wsXbtafkZKyaNXJHzFt
v8b+LjlUwBeyriW5iAlPHRCGLtu5oVdMB07jKUE1lJe1vDg2bWZy8AXgPjDHdACHgkfCyNxIdebo
SNYbPPBIl0LNbJYpsMmeFtK1Zbei9n0ZdFin0f0CaE+P80nZpYiEBDU+/FA3CIcJwacyV6a5Qts8
9/ehacs0RMpXyqrD4f6AegpKlYI8qGtNHaPPzMABCjbJCTj1YRjKym+ztZ8faLA7w7CQj/PL7b4j
qmDb6nlzceFVw/uZQfdKL0UzyA9u2NHwWcfI3c+OBLSMPtVnBPj1y/ZM+we9fDfAuQrr6USRGi1F
1TySSqWQpi1jUwp16wjwrFL5+7/w+V3wrgjjv35GpJQyRYAwD9E/o/lS34RktyI6+Ucs1YRgxcdP
8x2GVaXbKkF7N93SfKp5IyDkhMeo4N6hUHMdmfugU+7AbAq0hPSq6cO3x9/TSwZza5lIqrvOX6O6
BUHY/fsf2q3wPztc6vMcexMLZ4QI58GCj+x9ZcASr+Ht2/Psw4BrVJogFAzIeZAbdnhci9fyeDFf
zBgcD5K0TY0sw7t68SGFWAjQoSU7M9DxhYMAQhz50WE36RGuIPJy3XQEX6cWJeRJds8HRKT3iPXJ
rdM8R016/FDzQ6d7394Rj8Qr286RBpeve8zJxFoThbplB3lDFFEhkhwhACB0cixIwE3wlDA68sJO
qwF2BUBW6MqcXk49449wnt2QJAw7LgJRsbb+9vv0XZmgLXBlnCGcM/Xs2JuEibt9Uif3NC/OX6bC
H4yvGInFegdB31MCSoS+9IUxAjdhAerXonGOJtaSckz2j6XfjalX3s9i6ni1Hxv9YIuS44E8RvFN
jzk8r+KKYZsRCYscU8x7T6BrTFDQ7fmgy1X2+pJbbAFGV9Loi5LiLQKlIwcYwF0383vcvR/wNtAL
vmMjTJQyJahQYuGOD7kD1Y2oZPhFGqE6tJplWyNDBQCuIh9p2h64EU1S/sxyx4ob2ddXlitGFlNP
0/ifXGo+H5FAmmniOL+3qbPidyo0rQ+wpPB9Hd4+fmuEzN2Zj0IbVo9FBtXzQF1akrDYgra3Qt2G
7eS5TafvlNkMaJu85HBdulu+1yU8CrIFuMMsI029sB0G0W9Mvzu+tBMf5YVnNOmGzHYNs8drelaT
7Cwyx69GxQD57eJRrWxHO7eWuXGHq5Y+ztRdzdMEvArISs3o07Zpy2JnhLibZmqRzmVle+wUbCM2
S7l6LuX4EKHUERAz5YHxrAlhXBbZaru/+Z/DHc47F49L0lf38pFKxYQXjFIyTA5TcpAMuDB7fXzT
/h1O0W8mVPkmHyMFkOVQfirXNqjeunCq3Yz8NrsDDI2b9xiqV2D70oVR47bt93ItDhqmFOEWXGLn
04gb3B9fQHmv0tKZWRXki0yuYC6uPRruRwKGCz6wFGLA7nda81FDfQ3H6ZuzVeGd6g4hIfAtLMaH
5d3zo30l8SqZKEl+VFSt/JsLitqYcwMe2YggyZZrIEWm+a5/R/6S11xHlypa3D17ZQLbZRHq6sWx
OKhTfItyw/yRWY8HKRBp7eKNlBdeNPss+9eLzrkMoNQqt7E2Ch4hm9HQoNSeUVo7N7HqgXNWaSTa
SJMz1MFlCr4uGwU1s0gCJv+fHeVElosga0fbgySPbvG6q7JSEHBgIwY5Jc/NGOKKvl5i7bmAQMhR
hj2rfUS5wkIi2xKqH0s6D60bCt1ASfibxTQ2P6dglOU9OOB4kqSanX+PJY8khO3qOhRK94VBVpfF
j3+3pMefV0NOr8E7qogUicBZAlf+PkHRqCoZBe0cCgDtNkofTHtFNytnLL4OEn5EDsjPFdtXjQn6
KHFocnYNECoPK2zyf1vIV1fyYWdtvGfO2lI2eourdv9HYMkToOwvpH0qWOloJinTGEhxCybGpySX
CgCA2NbuABkD66lTfrKxL1d/9vd1AieN4B0TM/nYg0Bfg20yBE0kRpKg0s8DgDwtxwDIeV0qhs3e
4xqJfOWFmfQCOY+7JZP8uN6kBFnYt97NENGh2h5qktp4YyCZTtLgXeWTOLekjaQk58vd07R9vLCy
RBSvGpwDttS4u/ENapfPlKcL2/svrfRpJuxD7r/LNoF/k6seiCbt4RRB7duBoxkWwDNJ0W1iCSJI
NjVOWxjicsWpJMgIwtUbk13mZO3/dwzC83sOdYvldKMnCYp+D0RuonWFiD8oghhdFbu2PCh9jcNw
6wvh9OLTwKR2b0xMaFNLZT1EBAiS9TP32d/6XwFqhV0ybk8b6Ad1R8d7PxRKzoil4BLoFCfaNVnv
grhyC8nYNqa6mBxFX/4boMF1kJ8bSkCUnnb8E+4w2MxKiVi5raf7ry7HKEUQ9D8EkyMRk3Upsu/g
xbc4aornd4zGp/rljryG6h1TCPzKr1iIbmHncxTbpBBZlRljmQXR3M6IYcDekRvKW72f0SBc8cYO
bkXigGenODeXXGv0PvOm50BkbDisfeITbBpsYQ+3nF4vpnqC3Z3mLzY2XcXzL0I/3cwQRBbJYrAi
q23efdWcK4J+6JFAxM6pe2LNecNA9vuoOZCsrRIriE56vKyY03bpRPJU3bgy1IP0+PI5+adSJ/Vo
N6HBHnrJR9RLqqpQ8G46XeC5JlCg18+mLCPtJDqGH1qGQe92jdA95wPeoCP+N60+xLjWGBihSf3z
yEkKqsW/mHS45p7a7G1jYNEfsh6+HLQTPtywKH6qDui31wyHJb0zZgmA73/milpBuqy8oKY3S+GY
LLhsyOa92nWsAHRSsPtSmcIlknuLWFvhFuODR+h6s9c4mmGVnutc11dR+bz0fl5F0QRGr3ofXwa9
f372/j7q+TDpDJhJ5iElo5+MgipkNiXhhX6h30Yo/kKlyBtAe63KpMgF0e5D4drLJCGNArsxHl1u
TCqBG6SP8gnxpTceTZqoc1YsRDEo6lCCpVXurJdUvVg/vO+5BOa6S41FUYrRXnNHJqMYEtvrEN2O
Fm3xdXEuCKMxOYYeUZzVsKmczs40DqIrR9l+xzOnKennK80h7cRQ7f5PNIzFeZZIEfvSVtyjITQv
NNMWwI89OoI6OhO5I8UFsSxKI8mNEGkbgx6ZaW9IaryaO4uswExDHBqiQFyx6B9k52O2qI+7zyVr
OLhuwueVn7LD9XsyrFrJn8r3FSwbb2i/+Usbol8N3nli6D44gd45BMRLqozOsL4I1dirDzvlr06t
/1WD60qelhcpNogmpP8OMyE+DSWqajnedc4edbywGhucoaFMqQPABR1XZkVpNFTxH0rNPMsnQtsr
9oKIFTamVH86hBMkNKvKfNQb7m87dbdywkFJ0kEgBEcfKzVmVsjaseAN6oYuqJb5noiJwqgJksTX
Gfcyd4onhKTiHtwUG5uDs4a/1OiZT9QD8XmCpfTjwnEb7iwUN992WLjXWDeKd7ddLhyRRHe6Yp/0
tt4QYfTlSm7qQlRKher14rBGDVLalWE3172B1E9b9eEWZSVEQRr/HNPQQnM/wluHIm7MALiYPnvi
J8foYGYSnDDsqiabRU4vVPR2Opx6cBta1fJIvxOlM8YuiTinWBN7jB1thfatoauK9YQPeP37uALg
su6qE8KvQy3LN7vRNQXMHc+PTE3VZt2TB7WGjaGBgrfPoSwk7ggefX5GSUxgGB74mtRsGLnw+kGz
ugctRFL+mNGtew5N5pVDw7d9qCotQGFG3JkLzB0SZE2llYCBSbE7M/u7UfAWSt+TyySD1b5BgCKO
REkIGnRYuh0VTeVn7WXO8qC4mrN12p0PwaUfcVW+JstiHDxwahQTObMbGeSqwozmPYZakBrZaP3j
OKBB26IQDJq/j6nesjHtqXczkAk7OBWNeVyLG02ORMFF7BYqw+ZGlydWmCT7Jid9wLLrb1ke3yYx
/mfnrNPbLNXnAKVDm58KpSC1sdLpcl83fvN6zJHJf1/YpKHlEdlPgpUDYJkCXBRrfVwRBhUABh2u
8A+4FCQSUvJ4Jj3mnI4anVWLRkgYfLG8HKbDC31xsfqBN93bWlSf6363ToXYma5OLU/Qc3ZNYwUI
4TgRNw2pz8GWS+EI1zJkyWuYD1CyYyrmJESyLPk79x6obBJoUQ7typbZS8grnb7b3pVhveXsaout
6MvzuPoZiVtqi0CDXVokF91lbZbPkFC/HNQVv54CjzLE1BAf/GRmXcUWhOuc/N+e9PdcKd8pQLq7
qhyZ6F3WCvq/mZ9jIJVo/56bLSwcZxvY2qaR+m7tLaj2Z/usDLD4XC+DjNmsx+/MkLB3eR8F7xlS
6Ay2AIzex+eKZvQw+9ewoE1EbdELbfGX6Kjh03oXYXUscr7mdjWays3A19pCxW21XmIPCrMYL2cj
UNUq1dO32KeM14lMiUX9KVv65BVqzz/3Dm+vZHvKl8+E4z+yAxx/ArZX1wPqzAjFtxYiwb6UDf7p
empLow2hASYOoXDf27wlALMt5OX6GMNhBdXiCzvm6kiQ6MhUCU2gsBLsZVWvebzR02y4YhndOYG0
l4nKRXiV7m0UtOrYogLxSIzxojKMRoVLs7olJ1W1wqs0DxyOS8hj19UmdDvV5HAFTb+ArdyXdepw
n1T1Cj0JKcMK8Mnir4YcVGqwV89xIEB036A8GXfpjKSOX39CUL08GA+dSbRQs1oMk2RtzTa7qY8s
DvnQ9tf8TozFM0PiVxfweXkN2t6OEA2dZZ61MvERxMsn9HOEU4K5kkNm/mmb5FEd0DxOnzFUPqnD
Jv1smajKsUL81+7i/ciAnHAaffoW1sE894TsyIFluw4WZ5F9+eGctFv1F01gLgN1uO1qSzIPvgU/
P2XNWWZWiv+Fcu/FFr6x+0EPsqqeWjP1fckLvC3rZqNgBPQkuzxXUWq2+8jdyWaPWKiVka3hnPE7
SC4TUH1hYW/Wg78rqrydbEz+pFsqDNAAdr8HUMmJqCMuCbNcKaz0LPxDM9f6+R4CO70NkfEdlIrf
O56ErkE9uqx5/N7A1YLbDLi8fByj/hb2xqf1Meul7FQ8FOu3E+31gySj2BdEAjToFVTu9/n8Za9m
+i+QXkziV1t8LC7aEgLzjX0wE20a5p2p0NGbGnbeqzUVWI13Jw5lrXhKxSJe3pZ8wwTgVw+G3ZRb
P7KdMrmrZX1bH9tRDB04FN7noum+QvGYoc+iYjmDH0nAsvIXIl9G4F6PKj8q0nOgjhun9Ti99HJ/
cUuVydPURj/gBjS12vL+Wx3Fo04so6G6C8nZ3iIyzeR+h/KxRkyJdQt1qgDRuNrsWlBV35MQuaQ2
JnMXlW8ApUXkhZ9fUM/r0nyWhVdd/wG6yGw/c/ejrAbDOcPbv5MEjuSYSLFpnfmiMO5p6oTs3Q+C
mPlZWJ9cVqlPcEeweqsYSMfPlhbdsjc3p7fPXoS1uERgUz4dsWeZPjy4urPWqPqj9CwY60JOXIkP
76VqItHRg/J+xCNfCppWCfBasRPSZtaqIEe98X67KAC/FB1/w1T7IEnQMK8tTNvipbW7MLxHJRy+
tiZ+ZbUC8WopcnAjM/0c5F7rEErrBeiaZHsEXmt7E3zV7EOvGATlc4hlUbSvLnwqTkKvwisocqwr
mHXCr1AqGpFydoUiSL4eV8KAq2HO8/FONFinCHkCtipQsrpRM4vmeL7s+41rU3R2pbx+U3XhedD5
YrZ0q+XP04Fm7cFePnA4HLiUamNlSV8bCjIiUxulydr69HGZ7I/e8o95xKYmP1kcM0L8q+wpX9pP
cLnFYMu9eaZ5IvzgecxbXtSOaO6p9/wH0ME3GMqVYI0B2GO7T/qOQPrjvWsL+/KeQzG0GkHVqU94
KFEXyowy35+iaGPnjeJEfHkQcQFM5DhOUU//z0MQ1iIy+pSYkC9/e3XbeTFpJBkW3oBZ1ojFE9kr
BxXtjzA1mWCCPfz3AV/jWbqhwsxoVRL0L0dlZSLemKd5/fMUuzRMi8GZFycASZ1/KM6QHzIGuYln
qUKtcpK6KVgHQrNlVKe/KeLmJviUIvIES4xSAEpc53hQAb+OW5MLF426+dAS99F3WpBYcFxJ/oQi
7mTnF9wUVfLnutUEw0P8an1rqeWOw9Es+wcXnE6JXbBB8cMqT7L4lyd3qI4X7cGZe7FoFFImERvX
jVZmwHuIQ1s83H806xwjLo0396UkiqmNsm272gOptbGa5ooGbJcyFVJ3N3uHxO0X8dBtChMZMzEn
Y4oxiYmVaocA/3jTu8IHHGCaPwbFsS04rhO4miGhd32UBBsFzJ2N8ooYbEd1jhPYUjwah+uG9NmT
lIDNNBzyhHymTfSLxYOfJwV1Ht+2q1eGkVhKyRtVq18ZmmwfUmtpZorhuFte6VWZ59PeibsvbQ9+
UR6trCMrhYOyXwarJz+gBG5jQBnbj5m3o/oAICbCW5W42rRbICdrMVLBqyoAC9WfmBGwil7eQRvj
aNFbtoxywcEDEds/J0a+yKtFzpvl7dacVlZR+bssoSaiJdjabAvXuwaLhUHHw4o+EET5cwFTl6fI
Rvv8mWgFdYJrZ6MScv7enjdQTxouORC9lRWO9Ax4/u27ETKaMY8V/UI0SaZqxBwcR1qn5zgFPj4L
1dxB0j6uH8K68WtmmUb2U94wNHh6xj3IJkf4drZy5diygW048gY7a2KLXQd3c4OhIfbyuCidW4TG
z64ju/56wuVCj7efi5Usk2ekCKyu2HERAJ7eazjCi83TDkvxR7aq1hYNGXSCJT8kwYZmdDa0exf7
pg6kr8HosiiTSyOpm5qpNWqBYe+F150i8h33pWnYvEeVk7affYldrhON3+2xrRK329gH0/i9aZX4
Asw9oCxAW7r/1uoAudEZkyGRssnved+cj1K9rdvZdw2hWCSJvpIWkYqpGi6JQN9TVYNGtV1VI47e
+TaejkrC4HNOqB8O+IyWLAgq89WwbhFYPMsmVJq/B7odqjUbw38q8/ARI/NoQeWbhO0IlM33WvzJ
ej1B0LwYhMarRxP3oMp8AL+1Y+EJ39L1On1orKnPdxnQFU+kUlupOwanW64KBCgUg7N7GSIJfQCi
8jiu1rL3ZsNelUhpQFT5NL+v4DIR/PTbWjlKC+K8ur8Ha8G4RWiaYA0MPbi2azBf1e39SK0lhXC4
zhbKHLKNM4g2jwstyXG+iv7pvzPnXT8VOlbZmRysQn6Zf7jNy6T9pD71/+uj3xYyLYR3y02dvLxR
CjdZGD6rg85TjwCInZ1eF3aKBX6BAHMc4LTPZcL76EsgK7Beg4aVh65h6AkSd255ck1hI1rkVIpF
SGRG0LfMXLUska/EFS3FEQvk9/AE9wIWpygTrdtv1cY4cFqbZv4FDGP8RWViROeCBOyKB0F85h+M
aK0SnphmZKlAhOMoJoCttv0338Je5viJoTMZulchHXXvNVG1z+RtHx6TeMwgyR75S/SzeWlJdllW
/IV5f/zk8MewlRkSMq8GDmAUJta1oarpUGuE2qoulhoWJuUTDmw2d752DvyQv5Eu/ReTVlbUCHnE
xwpKe9lmjwY2rKn+TVo/repktI2Yy4G8q4vWeHPgwmu9s2zE+YEBUhdCQNrwQPwPBd2aFzTK0L6A
0hksCSdM5nVEKPgpVKOd54p/Tft1pYGhi9cb6WbnVkBc2eoGXJSwmKubFuARjxTBRyST3gAAlJTh
5Skr8/CVFY+vF4yovKolhTFltWyzX9OQ32sFvG5xq4h+RsshNSjGeniDAuB6T1+6zEtuQXpYFlly
fG/0fE50dQDvVodn4zPcGxkbxKOKsuwBfAhLdPvHRs+IW0zWzqd4FVJVw3bKCY7ABqj2cFGX46JP
8ufZ/ownql/4tq/1tbRZLwlsNljUTzqRX9IlUDL3KaID8l061moLwBT0wQ8szuuqOy6enAljHLDa
AQtqh1WfKUP9acv/3TOeCAMJKj/VfiYSF2tFp/ygIf2SFv7YiAHu0DuIPylI0848zVpYkqnvyt1g
fKlp+XiQoRezX5ITlz1LAaM1jKoiIwdrd4LD5hq9ZvWMjyYyzcLsa3mcfu0qkzs89sUwV9J4E8Yr
TSZVQaWpB6Kp002mtwIoXhlWUcvp3l7ns6kTf534evNyEiZKBEvrzfIqowMRlCYetJPzpBKUcKkA
BP+muFSiF6p4iT3HmOcbDoFjQtKx6LRbjAwJHktnQvAyEMDVbG6MMRc/Y4eeajH3TdfXaC3kQSvS
HQ5IO8yvX/qjOsuthu2LlB1jKEAg2MVyAkeraanKg3Y+i5lJer/07ZZxnzD2OrOHlkdWPJTrFoC8
L5Z7CDvvm5lrBRnlGa97irXJpd1HuAogaRA/SXRyvs1qc2m/U0SP1hPiitOYt9LVWE8uoOkHsSrj
8AKbLvD/8HjZHq7TAu2yJGKFLTaGSa1dFkcFzQGfX/SFJsZ+EGwaI8VU7ArQk2V31hDn5BZluiya
f7zXSfmNrzliHUA9jciD3RTO9wR2Al7NcA7H+gqOgAScz2HTR+eibD/Ti12+JrJmoCyzPKgK9n0L
MB8i+vAkVlScfG7Vmm2MnzjuKBD7okVvGWjmA0y0hcOYs4fLMkgPTnmQG+NG3JsypPmVBMJkf7hW
TxhdgEAUELBNpC26X2wM0Jip250LaeKRWaTTed8/BnJXGomEeXanogwxPbIaxtzbGLIkks13Wn2h
EqLDRZMBLCZ9rL07g6+Jy99BdAF3WjnAr+1+ObSD/7l5K2TBfqHf8eEhNedQYw40wFI9f4//UCS+
nH6BkuEEOpvtWoOPShkZ3o6Cm8/wUzoEz8ZBpA6xgcR+PVevU5Vmnz+vT9yjJsoTSYvTvEI6+wuX
rl65+3kK2T6DH8992ilzKSFSOyH1CrASuKNxPJ6pN0gBZ9glkRKPNlbd+SA3/rEOH4piPijkrYeq
/xtQA6Twpda9R62oC8B6hsXgooAtztL8X8RvKe/xIHu1Ho4SLV7eUn6nDe7h9YQLbEmRgYVhBOjP
RP8TgbRviASlLnzv4lYpeyKAfuzN406Sw15rE47jy8zBtd0v7ICEmRP9+an4zS844MGLM66D8LIO
7fXuyEdb0UIY3qNx+h+b8ML+6ZCy6+DEIBAufh7QTC3LEajh7OC4iGKZl9Nd4lqTBdLHrK14VWiz
OfNSsqITWgXvGnFgbW97fjj47xNeUbNKdHKDfh18y3E/d9y+7FUrv+hZW1oHw1s9KOC4zH7gxQz8
rm8yY33v3+B1vbWbyrixg6BXfF1cbtm9oJBQU5b/9X24EnGBCYeEgbGitfg51mjEMhzIdqJDVGpy
s7ZlEShsySarrnZ2k0379tM6JWN04BbeLjfLNlVfQbQNng3ZuEyASzFQhLW+D7uiyUPwmzSfbSGc
ItJ7WOO+SpgDYax5Sdsm0HBH2aQLMcRe7OnoOjLr9+ZLB5aED1BaxlSF7xdRfog9rAyGyvssucMB
5a9RVaSSiHcOvR6zIUC4xy2PJ7Dax9QD0vrvdiWJOTIRGpTK8ZT7FAt0zSeH8IcNx0FjYIb7IBTi
ff8VNSOfX9xhQuU/gfKfX9XaM5vFtmLmSs1tNcZqyF4c1Qf+kNZuFTWYhbVhbacjaiaODRmVbUhU
VUxpfGx6PDYsDNLhEWRMfH8C2G6ekhmPiFNf5ByHA8cb9oKMGgEZvEU89fDzRr7v1uf/pYUDNXLf
gjuyIa3xGLPK1MVfjZ7b6nQ37Caftbe1Lv+N4fnyErtzUGedRWz8jTETfUgaYA9Kkbn+HsFpFnvU
Vu+VjVAjDDiI/shWST7QvSoJfouSBxQBW5RdKQoMppogOHfKNuT6Ut5/d4KdA/cjMGdNjfDKQjzd
yj5QUneKUFluT8wy80IAP7iPMdw7Zw8yduyXxTkiy1w3haUL2cR9jpnwznR4hSMcsvwRKnpV++nJ
cOUbO9jp1MkCQ7Kh2ydCdvmv4onyaUw2htYlf77ScdMbYvPrFJAWyZF/SuYqoVwRQ9dwyzah4mc1
jRCyqCoxcjHQTKvzal9YVXcX6AL5Oxi2Q2FW7hoMnuBvdCr4LHCfn7punh5qkHJUyXE5XyxndTUj
iJkvhauTSXeYep/7mHmyHaWjrq8xqRlCPDZwhuFTQpdSjUJptHcnTxQuCTkFAwpjPysSImp5EOJ8
1iwNilQVrXk7he57/8NlFdRTkVycY+sHAkdO2n+CC0iN7K9AaBP4QtuHs7bJNLyMF1VvdvKOyf7u
U23cDQa9i9Wc5HkhosN3zsdKMS07UIkGm5O0FdcZAQWKJYVqre8940F0q5GAA07m79OuBC48UgOy
XzRqoHj3EP/1cDaGZ6wO2sSx1RBYBnl3Fvakaoiuov0t+vUoIMb8hx7Yc8LKFhLbBCo6B40s+EHn
/ZH459FogvauheAa3V/FpZHNDfc8m01fmvYDDDyfzW1jjxlpsT2d5qIkvOB0faRLQJS7mq/WUcvZ
RFDfrCQGntvaQPFLgt14EBNoF9TL9dPggzxKW7Ng7di8iH7xde/GZtrG90NADt0p2gBd5QKTiYbN
ZkAvpkbRaeYeI+2FwZYxsaxrXYXKrIHATOCJO15AjqrFFq8liOAkEleWqU+dvXxmonndrB6dfnzN
QIAM9wYKlquxYinnVHKS6oQtXzuc5rweB1v6Q3Hvnp1OTB9eVY7kuRj4pPkW7qFI8S8eihN4741S
tXCJnt5okHGYvmR1ruXnVyjqsKYBPNzD/TLZgBjnklpsJRn2lxC/217ERPwS23gvd0POkWDFdfII
hS86CbDikxt+VPFtU54LGlau4ay+UzdEj0sssnaeO7e6zvHgrpNF6N+z4Kq+Rb6xJb/3T1ebDOa/
FI6t7DXgNrN+T0KVi/i7S3XVZzoZm696nxEM9bX+/XHwl7czgyucjHVsxFCK6P6LcbXfpO+GKN5x
4KCytvpTQgSJOlzJv1jMgOECMjmoGurnJ2k/aVrnEbMtrkUbiD6okaFp7YpxyCMUZ3QfN2lPSsmu
hU1hlarenUVjFwvDh2xZSUPO6OLdfEoUFwx8RlyfPjnFnnWBL8zYNP9dajIBmH+jEwso/FVpkGxw
T2TxBVuLQOBDPNzFhrxSWrb8qxHpBUUrA4rTZabxExXKMI0d//88H/xhJBvmwVC7cchDR9Ua8Rdd
g/QDhaFe+/lYJRYQ3MxDuxDlCZDbvdWM+vRsqj5N9P94iN+dEQzuDfPpspwWwFurRbVifuXB8HCW
j8XxMhur7MEFMtv2kMqLr9Ahwg11CZehX9uF9IvD17KmRuahjj2uKG7GaXfS3bRX/EMjBGfV2jkF
x7IlkPaxr+uUxOwFBoMxCDyxITQldzNHMnjsiTFzVuhOHlM/JXbDDsmJES+z6qnFGgLYDHU+eD/j
Xju+9G4/ZH8AarxBV6KRuxA6ztQfgH8FJx+jGJfiTa348lM1skOQTFAhW43OYhHvkT6wrW1eqtIh
uNtesxeoEzwfAS8t17xE9IluWLWAJ2Vn5o58sNKFbZ0ewD0gBYAyRdJtDHeiwg4d1jM21xdpE31G
BVyVTYNTHclUcoOWOBQjSe45UJXfGY52cVkfTmA6ZBSHH5PeYxXFk2TEvyyIThdhjBucnYcQnMXT
no6OS9T6t7xWxvY/ANsI6LtWgyOLU5QlmnSX07X/CFqj1pjTd1qOKEb0JlP8Rgo5cUJuk+jnOjDm
88D7jnTTc+EuzesLA2OpoBhqj0QKNcZPC+2JAwxgr+EWqyeldVL/a3bDGUW8ZHl3G8dsaRPV4vzy
4bqamhpiQViVhF3YCDwiFFHWANGufAQQRPYQp4RkR8SlxV7mmMePNlwx5OrWoVcDcXD7mkolc0Bu
M+TxYae+ZK2/gLw5cy/KtnYsfo7NlYjPNrEQ+RuiuyUoGZ60cn1AUB2Y72hnyrL4WKm24VAuB5yz
1sRoIjtKwg9Yj7Dv3mMm6Wl7n1X8Qsn+iUVKIU/AQdNx6abTqaduyp7jUXzN53FmJ9df8wqbFoT6
b9yQQFWZarGvUNxLJA/mrpCXoZoe2W2l+ydCNJ8Sp7voPUxJAaWWWjVXYXOr95/Ww3JenZc+lDxh
GSG0+aSA990ga3iULAM4tW1p32prDWJkE5Vmv08fI2gajiP1sHKeMwgIME2hYzjTSToJvmkq3ylm
tJLKzSlXi7mpSeyjgjYUya64cjBNFKXWCdBsVliLc3J8H+ZSactF/vn7kQV6e5vi4kSfoh93836+
HlDNZyhXu3cJlg/0gWec5rdPcTsnWjoOy5TwiFaUf2UHpeyy2XgUrM3BTfp1S7eQ+YFUqdIx1zvl
snMgyFoHK3ukQc2A8VdGu/JRb8bH7oTQsqrCpHGvjNgTNYj1TFpx4Xg6wqio4bnxOrjGNhcldaGZ
jd1nakrWjDZnqWRthQkd0VHyZYXsuifDr0ABwwo2BGwnpjpS7ECoZEeqHeMbFv7UcFkZxr7HRvJC
YjBmP6FjD7voEcUohhulpnDATMqVUbxoc7R9Ejs/qZc2t0Q8onWr+RZs96VF8YWzlL7QcfjRy8sN
daRoPfAU9+HXW822pHIu1jcMprSd4Pb/8P26XvMFhE9bDNrNpoixWx5gV82T3A8hUNjRlopGWatd
mItHIZfWB7CvNiIRW2hws2eUOUvHagzMsIluEot8hQLLsHBG7j2V2DuGDZjAEv/J1yX0dyOBo1/8
Aq1yjYRr/wyyvDApIIerOC9OARBYFNqcf+LrjGSDQI+sd56jz1V8NztwDG0rPAMXRoaYCljxYhac
V7XT5MOGUWtK0k/pEDQVemRL5LKYhIbxEmRp8KDKMmkTrUEQHfSWKKN8DsK3M7MW6mVkKU1Sz9qg
kPzVCnfUIrse3qH55xGSh0jd2Yw2H/tnAseIMgoHSVGaIn0mF+JijIjuU60LN6gg/juIjIADCyWz
gi2ytwo0GzurAn4qT7b6Pbw4PsPFYMJiEJrGlPt1rH5iQ0nk40E5C+WAukzPE1W+ol8JzzvvdCAs
IbMF0iWHGDnfbSnqFUhWO3iLfDU/Re3OQc4vxwWUlFKXR/2TR0CWt6RsZnT/9ZPp4tk7AgQITWsT
rsSxkYTByGLISvUMgWHwZfS6rEhbbMtx19TUK6UQ3gjulQCQmcm6bL5RtbCGXkIdyRbwvYGTlJnG
Z6/HY2fwXrb0NMqnmD8r951VASZbUfNlOVtDjE2ALfCYX/8wLINsS/9kZPrpbhxkXnLAh6KODUhq
EmMj6P9Wa34gxLP2MxfMgaiskvVzxPj9EdXxSguICdOVa9x/F2JB6b02NvmBO08JqkDTQlYxZP/M
GS1NBwcfYr7HGYtXIoc9okCu6jq19kRaz9J3m7wWktR9oTxjZX7TcRXgdVUnJGfVZ73eteEF4val
svVzx6ooZEwCgqJm4RdgieRhctKXud7MxmEHfsQpS4Mo61sQKQxGV6lqH/4t+FnZAyLXiY3zS3gC
ts4IuqyvQGtY+t793cvhhFww9bEPDPpcD6Ph1nfFKLzCZMHss+2Jo465QwV0UTH9tJpGRTq5F6YA
E1eDcCXB2hlfr9cYoRzEUjTC/lNiLk5Mcjtoy6bgfzc6iqv75YQOAMdnMbKsRrO3xUZx8iW4SyGV
l3Ul0DnAcAXhNxRsHXiYX9C6ukO/KrhvRhaNClHLu7iVbftFERbZxUA7Yivcfv6Eltuw5TeWAZas
Tunrkti0mhCQP3hSG3q64PB/bphhpcO9tagIY0psubdx8XqtghyZuemg/it6hecHtqzCe4LYOB2e
sO9NhXFVYEOKIBwKbu4dw7rx3ococM4k1O7bzXLnIMuzTCaC0K3EloMRyvl2ZKfQEFISk2wBMLSL
UDcKR91GUQyqhSBHPb9K3cXyuKJdbfxbdirAbR1wuK1zIfgFRypCPCdhftp3839zFsY8f9ge+rPg
xUmPeJWfL2rCIDoJV8uHQ/xKzmgxrsSV1ALi4JzIN3iN0ngnIRtLXEBNNHx/VK47aw3zQkj3UQcH
HlKYiJulLTPmeLylrCbbHfEIVPoar9LQT9wHdw/GwyZ7NaLcYbd5HPm5fp/nUstAeac/TNwVUPex
5ZoV/8JqZfHg3qYKbqaViOoCN5b3vN8G0jMg3hbEHXfN0N1HnQhybWHhMe+dTpofSijfFnzNQOnu
asDCZgKw/GnIulw67piA4MxHmwJoKazhAth90DHlhBlOARwohnMe6qOCEribrfLlJxoymvPYDrrQ
gyVGFDzEOzt24HEhR0Akirz8BDxKDrddT6nA7xq3sNa4Wi1SBKSxOd8C0sgmiGcc6FdgDkMMum7d
++O6WaPEmZak9J8mgqlWxWc1YSZhWI1aUCb/QxaQcpz311cZ1cnvOHH/F2ERdfeei5mEmtvNK5c6
B4i7Fbsh2Bxl5jhHkSbzX8m4LFvzmGFgI0C3+JvlA19TOhRHlxAvoncR1xJxaSxm0WokSTo4VJkZ
OPVd883U2aVZkTCIng8v/+lGLOox6TVkM6x7u0BmSQrOgaIhdYPZMe3ByCcf2stp9KKau8szpI9v
EIE3PbiShr9IoBDr/zvpOms7/pxnEvYVHGzys0lcyE4TLnHX+LVf9LFZ0gFMmN0DUet6I4uJTW3P
Q9z275bYJ9yyiJ6nQhdTuAW9n/vLbJWFkpGTdBMzhB0z9Bfms7XPyd6SfTsLaNWX+Ih4/oIbSucG
WUJj5HjluJAdzk3OC+EVQkYEqdQx4TW4Od+wxl1VU/UlulXYDirh4CfCCEkV3S5uQEVyBC0cVKPD
PidnD30VxRPOt7kgY7+nlXlM4h2DIWIXQguNfClqaF4a4POjaG/uyJajSyIy9iS838img0SFnW/O
dnOGUYQKanVWsNX8L9xdtABHPfY4YpZGEBZcxsrl5x7lA1Yl1e1oiiEafQc33Ja5VK2sIGPGnOAp
m/tFfeAArEXd/EkwzfhNIV+59/L+7LxjIUs8g9VEwfqDdMTCmPbCTm/p931L7nNhy+MDSQA8s4hO
MmMZQ+benQzIFUvrMNoga2EjGxUvrCs/pkf11/iZtZi2sbwmacKulbg6iJexGAlrHIIS1BQ3V5Kv
w4l+Lc5VwO79LuUcvDKPztml6ZthiYLNGYnBea+stFCM6fRQMG8srV9SKZ/Y/tjN/ODC9ZGrKtst
fh0lpZmyPk5VOm4GIqD3k/Z1jT5/C9dZG2BqStNp+OdMRElIGcxnz06l26LC7DtfC/MoaYfEbE1f
3OBbMza3TNx/l4Af7XXxFKx1wtoYu7vclQItZNYEoh6pzocgoXlYeSfpvIr1Pw6UQ28Onbs4FcmD
3TQNa6Fk6ohTE+RdSklsw9McSeiPNQ4nKcSFsa+Pg1gWf9tEjRizlvd47KzvNqnKe75scEUdNjni
q+Hwvf2tK8Asz64Dn8kdOUEJu63DPz58Hfuiz+2zcQ4/KP2eBTEaECdiVRXglRPM22CGL9UjcGUU
AUUJzVAJUgwiC+clq3/2FpWf0aSAWwKTLqhH6jda06BAywxhh4nue3dQQyxywB98w0zViYDTWV+S
o72QBLwG9AEUHOReGfiAe4+Py4YUE9KgqBSFvCkFCiQIZq+AYHoFjYTgLf38VRqKqaRaDu0yvJRV
q4xjhvv7BXwjbyDLvot9n6BzAPNBoVtdfBhD3kbSEbA8wz3QkniN0fE3ys8n+80NMGphscFdwEba
UpnqXTyutndzf/WVZPttJ/z3jRjY5ExKXMm+GGLLjOPXBRC9cIlVZ+723BuD3JwYyrNPCG8lSV+F
biSvChaHcbRLJZYjjXvggtjGrbI7qkOEuska6SYEIKrbyO9VpNV7rFxICMZJLTW4Sr11+ASQkWej
PajBt1JjcJ8YrA5dZkkFnpqSOid9lEpJYqdqoh6MSTQRy+++InpdDROjrRXHk4Dx6xarQokeFjkV
s8vG43mYBzjLkFwhePVAcE+Y4dOQZmjs+Ji2sgZ27Jd3/ex8AxZaax9oYVR11K8ObMIYJuXPflYx
84qUOTGTRAAGKLx4S9vgbEwxrYYh8JPoaeA7jq/fWmI5W/XyWGT2I6UJ5ozRJpR3pTY6dAXtxxJ+
CC7WdaXv/xrz30r2ATZI0i6c53xQr2mGxbRpcbtUiwchVRPtvawcUrmIOl//Ao/G1EoXWXXLUGhg
zlj5cEzXf6v7V7dksr3VNml2svvaVbgOJy+2RQp+swGyFmOd9KwgFKiQeNNfI6zCnaWU2xtY83m5
xU5er+BbSf1Llhbkf8LcJmgFXxyFZwzArS79NkzXML+9ihM4m74KbsKbmCXWrdX9ARwkPyvnc25C
ZJT6msC2liBsE7hFdE4nSt43NjQ6ay5XbOU+KnlQlXHk75vwgfai3hRAMx+S8/x8dyyVUN/FpzQw
r8BztE9ei2zUV8d8Qd1VOq4eXdyb+9thWLBh7qbs3h8gwqZ+TKDnC7E0SNps6MA4R9F3Vss9N8km
XqaiTi9NxGBF1BrEpsyzoc23zysPKN5TVUG94dPFOgbQrO9TMu2o/0nDmuqCq1U8UkeLKBe5ocy0
qQPCmFHtzIbvprrIosGFh+yXBKb2TmlI1tnkeA8Ajdcs/2wkxAIwMesN8JFh+9JpaOH4RLCkHT2A
TMf8ZTHvoLJ9nsExebeJPpdUpQX0UOPqRe58qs3Fj1XC61fcrTZa/LETcFZ9rUMTnNxBWwD1AFnU
Bizs1Cg+PMIUxe+8Adt+l6Sl0nQJgvHiiKWn3uRVo+TvXT8e3ndGYLtweQSyLVDCt4I3wBSB27c9
5HTyKPnzwR5xO2iNeXHs+Gju9JUKdqP75uk7IOzkENrlRIFIjYunGxBs92lMmIfKjmMQkdGmK3KO
MbZN0HLuie/6LkqtegqrJeVZVnQBVzITTr/0YadushuEyWv43ggX/Jp5f8spyclKbTHAdmmWEI+4
su28dh0QRyKSFdRKceiyqGbT+PnEDPUkpeYybNEjlMY+vHdLs2UXgfip+gFjE0244nY+CaP+M2KG
9xpxwije0a/AAocS++HGWFxppfG3xs6QErgV+aOVQAJNfYZlNRq1fOXYnu14xEf2rQ+/ar4GwqFt
9H/qMFazHnmGKi+R13VKLH52YZlLIH8bEaKhBFUglNpr5L/DCV93xclPOkT8q2FIKM81eK+Kt3wD
8D8W4jAdj8SsWd4hS+rpaEd8jlHnuYxvE5ldmPTiAt29HHEhhfOa5e7HedYDr0ZEKLUH52a80xwa
k+MfL0N0lnJRClL5+NZcEgw+fX/XRqT5D3chz/0xV0BTg6GpXhYa1HQDD6oZkOKY4vvX1OVxhu2e
MOjkJkGojSmTwaEm8u155NMIU+DrZBt3YbaeIo5sgpCcHm4NSVe7Q4qr0gc70X5MmFN+UMHrJ8VY
mknTe8GZT0z4coGHDB65Gm798bxe9L3sTI0nNfdQqkAdn0q23nMnzYL2Hvja+/YPwedMn4Um5jH8
hC709N9wIYCQi5+qSdtAgb5Lr7AJTzKXHIPV7uDYGxZEgbT7YC5fHQ067p8nzSvf2iWkl2aHmR+0
GPJuZDqfawY78SkVXzQGPh7K3Ht6v1abooSLtba+89mdS/3hTKZuoUOLf99Dq5xaRgh8eoP+eWPe
6OYcw9ThmPFupgrvSRzv/435BTvPrixfxwfsY7kA0sfe8JdI5/YVghcQ6KOMRgX5ssywxCKztBqH
heDYCu0dTTn+raFY7fmtsFcf2CMy6iOiICXxFL9sK/aAvxB0q7ZQHnzv6GZHYml7/fC23oeu2fDB
LlrnSHgWrws0Xx6y8J4xLn4t6gvZR13kdi7tnzjCaikK3l02Hp2gELqmTgMh4Sd0CBtBpRrWEKw9
E3fTgcaFuuy88YRdtg9tYgiQhuRzCeCOIBDFfn4jrbQEJj1qdQqgYYLR982PgHMtJoZ03AMUo/sz
HPWYd5dRgDej5JO2JpAqcOuDbI3UoiyQ3+RML0nomk9mYnYkm3EhLY2WcRlgcswvNiuP/0w+o+xz
CXSQxlHCBaFyMirdHgHbUQ5UV3DFEXDy+LOJ7d8RpugawS5weSLn0teExw4HYQW3OcMIjbLLXMlr
Fgk2N8+rXvVqL8hq2BWvCB+C6cByTt+j6+QzhIzijAJOepCjG01am5J405mHzlAQa7pVEctGuJ2N
hFa4SxmAs96tmAs/l40raiNo6cfqp0IbOyephkmJcS/uz88mm9Smwdr/ZklQ0AuUS1lmtCTzIOh/
RY5iWjJyNvUVcCG8k3xmIvPwGJcz6btGD+YjhN69nlJLXw2Qfl39UczRdC8gBTYW9y3xHhLALTVV
7jWCepNSlObY0+xAIJwx2mibMfsSLPy1nVKo9h94a0diN+tLgl0SiGhtOtbhZxRhnxViNdWrw7kc
iz6ibkH3iQJJ//iZkHm0TZuuXcwOepDNPmgg9GYJKqHe0PkRDhlNKuJHPJgnUbXmOSj7a+CyGYsg
IhQtPgNN1UOXTK35A68JsaiJtpl9WX2jMgzXEHOzFtM2wvzhVjBCAcL69XM3ZeE9DiHhKMA5d9KA
hB/TWKYz/3EkqK54KGwSwVEGmkg+bJ3GM5rWdY6B4wFMoF1zX9ZxNgsKNRvtH8QHow7PTYZG5vX5
ImthQSBPLGNaKpsxqCMr2Ax0TGC+yRgIY1lXhYeGdeD0LL992hE04PQiOM0gWOOwbygCRFDZRPGH
xNzOsOFmPdQr86Hla8j7AlzjED0HdCdKhll6RWceBOZkkQroPEeqLSOz1DpWnR2cp5PZOccH5S2j
GEp+PwWCuyAOxPVF/w1upylSheOZ3vfl3n0drdqsxU8uhVgsRJQ4QN5zQO929qxD8vlRlG3NN+F4
RPgx2EvJZlP6cYpqeH3dmvXYE961g+iTPLaleq0R5CAqU0M6DTKV/z8CFgjcUoLA14bb9H0gjHAc
WWjJx6g4MuhEgQlboRZAOQKUDv1rqY8Z5hizHUxXYQg8cedQ6eNm1ZGI2YyWbqyLpR9sWkS/pBYC
CDkAZ5ViLij/1ZiNtfobV3amp44icu8aVyp5/G6tTfDUdNpKDqdphklCQGL2GFyGa0sqaXuqbKmR
sBWiZg4/cle/yZV9jREDXElJZ8SPVMTasF0mmQI5etpxHfc0JUYPwHWJuvIqb8+sU+SCmnNVNkQ/
ZLXvZSbdDHdWSav7hE12zoEUQBl60EryoIdsV84FvyjSPKNKTnxREAYGxNd3lqpNpkIwRHMR3tF0
4LSidZUOn3Di7ez583tgxXPZSUUY5ZHXIQnd6ij61LnB6wSCImcG6mMbbMGB1UbHQQ0SBz0Dv3Bx
pCJEcvVxpRXInJmW73OMYcuz+h3fdxc8jrqr7whJNMTtdVdHUn+YlfrS16idz/zpLHL8mHsE5FCJ
0jIkxNpemakiAJuEgDe6Wsbx1XEM+9etwhEnAhHR8e14cCu+lIqI8VD/+YlvLIocE6hXKt6tv4FO
+4y+JeNGhIrbxHZ6zGxNAK3Yk7zIIYPy2UbwHXyyOE+TFXazDT6Ghyh2ALEQitCq+GjgxgRouepJ
4WjbXkh9FkLUzbZ/LVtSGQ0zLQa+NE43AidbEkX6l26qWnkXZj+9C8LAYR4Oq7L1BVkRWdwsbxgP
Bf6Q/mw17n7lpUpGeL4KrZzhxJQdQj91GWUwOmBbYc8WW8u+Hv4ghw9Rc/m5i0ltYg118PLTi81H
6qwBn4qQuUPOIEc146H4iEZynrGbdXff36f5KCmMMTHJrq+9WOhJfIrXVOzgT2sH790O6LAU82uK
erqvAnUfE9TelZQPFygOZhCBk8hnecD4/vrYAGD78hBdveA9442EcMqt8LHWoav5+IWOmj1xyLZb
MEe34WEIvEc+1/qmq+s9zFtDinsbj3DJKVIQ7+M2t3sIgjjJiaI/WdqvINNzuZ0RFCnijb650Sem
+IzSCsgdBa07j2K5K4st2cM+rJYwkHF1Uk7ucH8D9hA7rS5V6CgdYrI1x8rEOqfEC6YEM8zipodd
tGh1HYoiz6zdNVkFy3MB/dkLX0IhbPU1+SNmYqr4OfadGO2GTfyFAousTq7h9KuR1Co+swDmDHBX
aZiTxpyuQAyL6Q9liQu25abAUoKg6yqezg0IFCr4On1qy6rtOyoEXMAXEWbWjiWHZMjpLbD11dmG
xGwR9X0SYkVy+09vZbUDCLe8oOYAby3f0LnSyn/arbHGWN2v2Sve7dHk9zDm4NMo1kKqP+J1qCS3
iyhplURl7UGnRkTE5UezAxHIkCU3siKBmsGQLCSGrIdGoRGtlMgqGYfhjKxRZ+VXI2QyHVRxcZIP
1BtADj2OLp14hArF7KTY8kakKtzH9TRQbEvubjirYPVMkOVNFZy88zEhR3vaFAy4d9ehG+R2VabD
8GsYToNkY2dF5t1rO1M38qKabDNOAWAqUcUNF2OlcnUpB7rbRkJytQSyX2ryACUnoArMXV4zEnh5
X0nL9HDVVoEAMfu3eHsj0TI4z7s+LChXKZGE9zGvb4dGPtiJ5iqF9iUIsVISiW0/izY4kqqUXNBk
xtCj/xQFdGuxPSk3p6gLoilN4kSJZDwclU/V3TmZKzoVgmC6dI1viMN526P60VfS2w/P2BWntZX+
HJFQcBRyn8x1KCy/drkQYbz8YMJAWhQeB38qr+tXIqaIanZgg5bPFAoLyFiAfRZ/DKJi7ymSyLHG
2DyYLsnt4yFYtfJOGZHceZ2+qsbehFlFuDFkWfUgMQgBzebACn1++5pZN+aFyBqTk+B9mR/2vFFW
BsdTJNjb24apKfjnceYvSp/wSU1wFkl0b/Jp7uSZjdRlsz5yI7Ru0TdCRmDzhBtGixPrq6qOQpf+
hqEYdjkTD33hoh/KTzQW6bXKdX7umbkU/6nbGS0lcCU677xe8V/MkOYHREwrQpwqoLrI9OIZCnZU
AYqVXPZEfGA/mKGPSCYM6HysDCwwT7V2Qmj+SiZWYMMd5jHLW3MLS/ojPcoDGckxDnWBlTk6SL09
LMU9Ix+rF3y8nbPq+gutcWayT3C25N8YUAJSQJjTQgydR49CQy7c9sn/JOuai7oRwVCn2H6zJvVy
AuL/FFlCq5qplmKb0Krwf/DnvCJ6RobOWoFyZNGD9shdYt7pLvcALIaOtLXDvgEDMQkU7Yme/kC8
ujWWFUo5qTHKP9TYqjWuhNA+qUAvHLSIrtCSq0C5185pilwN8A5EyPvXNpv8E1c9ojrKvyX3XYGM
n005XD1RxU+RK6lWSYRE6o9y1Kp3DVp9I4ENETGcI9peC1qF8zWDU/UE5bxSGrP/TkXV8BCRlLbV
YXvZLlDd0rIwwrgDKPKhJ+j7IwwiDl4RpnovCMH39igSwR/8GVg+S2PR2Msp/PzINEU02CYx93OB
HLR5pdR/ppVLlznAkCHAXgAVvx7Mofw1U46m7LOTXLaZ5J99ykwlIXRSMBMnl9yeM7EZPI3jcQMI
WlUpyPVtSYBz8Mv7UC8TCR4aIN4BOwIYHtUSy1rNphDI6ZgDFXodV0pBzzrYQOCFNLYNP9CCcAgG
lchvxEFR6Pz8BidInKBv8hToCZqqh288mLZYQK6ccf3pK1TgJYh/ov8jVORDovaYe0mpcfwSLdmK
vBBFdR/bmZ6WDhduSmn81nUJazgiZ+FU/Hqx1L6QMYvpC4gdHOAYTMyV7whxzs5V1yWDLYOi5WrR
YsTeB/0J+bl96m0Kn9FB1b2Hw9Z3xipruI3Ycc48Z3/4VvA9wgudhpgHOIuivanufxzkoElmeNON
yijBTtneETkuCRdpEE+IOqQ07x4gOznrGWV/wECRs2jMMB20q9D1lqHpSfHAN/rINPoD1G7D/c27
nIuF6VkltPjwQ/ipjRQldw7ecMFIYA/sWS3g5wLZ1DB1IHJRFd1PLStRvh+dIoT5ZkxqHJzicREN
QBh/aXaY8N6GdqT0u5X/JlqrSJv+ZzhAcm6OWD88el6gtZsXzJdNF3YSiJXcpdp7y8f2Jy2x6NFL
SYaNl8n0k2kM+26oYjlBx027MR9YH7THBfWd8sSj8nIM6TS0gI5sabdayQrOgaoOZT7bLyh3d8TF
94KRaVpqGS5JzM0kX6yAzEUHlylNUZp2XveargfUU19sbnjsBlUD0Q2BHBSTXAZnNHi+QO3C8vP0
8UbGIvY73UULM91gYlqLVcvxxdZC/dCCRSgJKPbqMJ12cbPBRuL1GG7aHrvA7NZ2pD5ZKbfU+eN5
j2dvKAVI8Z6HqfiVHj5b8Vv303HzLS87mg/2Mvq69UvDlyKIDRAUMyTQwEQO00vxrRO7u4EofXX7
JiHUibJkF7czUWSxdR9GxsqRfj1FmMzQ6lQRdMy3sg0e6veojAM34uGBH0/U4Tzq2DBEW6cCg6ar
cXtomEZGWni9rAjClGWqnXPawkenWq1Oviakaf55o3lhSXOP0r54parXn4yXz1DlICMdqUFl0OYU
hlP9bV5snP8ZQnUqcP/xEGvWBbEexPblOkWEt9XWBAoxGSFHt6r9KTalu5LeVMFhXqKtSNtU7mS6
CAr0K+gFEhEq1BvkAIekz768qd183kdoYtrX52jqm8BYkheAMnfYgrkFAIFmJOrazVpBHgyujVrT
x1BB29Rx8D2Ff3MIau08jKfK2EgcIq6vkd+Ji0aVbfIOrI9FFBPk/1yQj5NDZryVv+/Vi4Zf4Ewf
5tvIKLls34sjJiXkAC7+WemaORS/ieWMnaV05k6YyoMiLRn6q8BoXsr7vSXi0PA4GhkRZgrXQTmG
xmZPgM4TONP842Tum/1A/0pqqDEWErwh2hGxcUVZazJkHj6hbowfyFcHy7qjEaP0L+dYfzsrPVVN
loLSlMrHw4W2fMExlVjHIYt/RQhabMPvkJRPegtFqTujHujAwrabVlO/8gF+4GaFwwdr6zwVUZwy
VgSg/aN7HylqvcWhjweIF/Io65xfYigiHgTX0E7Fe0BSE6QusvoAR7xcnbONQpD1f9t9Tjwh8yfx
0jTYFsYBzMpRzTst5U6cnulDGl6GKn/XLtxYlDdICrUp9XjUWGyYAYFWtTNC04PQUDN3j+u00/Gs
zBrObJ89MuR8oRT15/1HY8k8eBGQa49J8SrzxSdkybNiOqV05VHBWC6dq5bLkHS09YXTOohf0Nur
Krh9Pace+QFv/pYi4106vqcXoSt9OVBnPtoJNB6haiZOR2Ku4E222LdNAlbZRI1wptXvtiHbWcBG
Syfs/SdZuv3WtKdGqU9p26ErUtpYPxVii62Q7cg+57rZXBy1A4LsNMXk67wYziZJIepbuOKMemyd
w9uh8PezhXRasSzQfrnT/n+tjKkG7VDN9MKQQT4XrUenTeT9NjnjGAbBPMjfsFmzZy+cURpaDI4Z
QuGFtfKnAcwNKJYliQj4vs93Q89Va7OOAydy7HBWgFOrhXYIdTFO2Jy1vDQgbl0dBAkdp3NklC5I
ertu+4fO+NZQBWqLCO4uFEegcFJX2abtOdR1idm1Kvtwglqiic4GkL8Fs9HI9M166i93sV3wX9of
lI30moPz2pKjIcjGO2X0cjENKhQQL9qoh0GGif214yEiUzsGxkqElOQ+X0RuotCx5+efb4qhD4Kx
jxaY05/QFV3IkwhTRG0nAC0os5K1dqzG+Ulqw+XYbPZkMwRZn9LhwhSh/WzqatEhkKGZCuwDwNug
teagNqIx0210ifwv4Mk3sVqgIlPlyoCaYIVIUtLZHs/xFQyMGbN8aPC9YDeFe7lTuWRrOU/1ZR7I
7pSmqyBQGKxu/KxZ6jQZbg2QPmrYCPbL3RgdougoqoZgNlEl00q1KMHcOV2QAOsWBF3ejX0pE3Cf
FRhCC5kEXurtBOm28RprD+JcSW6t4a+5P1Wb5Vi/MFcChhyLoXaihd/6BgD4I0R7cipJnXByl0a/
/WvZodCExQwu57NcOrZK/6O9npLRtrs9gl/qwQ67hoVsxv5CAkoazs/jAkHFE+S14no01YLeGDhW
TdsRUMguRiLHq5OglqjmJQ/rXQ5PZB+iJp/7g7MD2yGjj8S7o+4A2H46Db8ZDf91Rj63qTyTGuGb
CTkLH2PelIFAz0mx886JJSBJgQ3n2U2gctAvpUW2X7Tou+ioRfnNLex61FLq5iNyQ3LH6n8CGOYy
cR+CRvhSPaE1ulwQYYUcwZTscADt89x79fdm66byjeqQo8tAdWcy3eeUuNYBYJsgyL0NjLYOAiZd
GLaZ0ZqT63wEDanb53rp4Rr1QfNMXO2KtBgJJbcgEErcE3W3VoDEw8NNassXVnhjpGjaRhUxzkSp
2GRD1pT+nsNchbYDAyNihReDe4Bv3Be6yCS7/IKL5xRO/ap3XDj6Ppm1/+z30tkJ12XD0geLmTIi
AeNPhnKxCCmhRbLTn2PZ59+5Ta+sLbeKHUaB3Y3AmtaoGAcDaVLvdtpjDqENs9wQuTB7+89P6pBl
KRffnLmEkqYQL1XSkf45dZS6sI6PUGKRBkyxe+rft4SXtZEjL1aoYW9NQj1lJu5PR/Vt15+yR646
dWyA/hmNbLxF3XlEA96uu/7LQ/bMWCIqe1OC5nKa1j4msHaQkw5ZE1kW1IXDP7Xw14DI2VIwzbks
fGi67C/s5aDMzfvpy7o0Kaes/MZ7hAF9LDpvn96EJSxqZAdVmHPhlHCCVU520GBP6Ud1ORUd4Jxs
YIm2KaQH/tjDKdggH2cjNdpFn5KbJesFDLiaB/7w8K71xFuTN2ZqATyMNStoeA9Gyo/leoPdYCnG
ejloowUtV6avTxKw8wziDJFqX0n94nGtaIrF8lgermRgjRHW1oQE66KfIwtfqkydkzFolxZjHJ1m
etb57N5LoPz8sJ76Tp/38ubQKlTtRr0UZoUfcjVb5MlS0btgAvzvB9xEjDI/LEtycJeE+GhMz3ka
tsE47oyTP7Cn0kcHeHZCogjrYxKxJzUH2IhF5pcOGeBZel+3GDkZeq1x/m6/aJVAW4bGx76D5TeP
IWbnWJnyPJt5yo1gZ31qko03wbBi4JYKTQwA95d2NaCThONwUn66TbsjiAVLrKJp+Vm8AwZef9Fe
nydXsYSCzvAID1erZYu/n088rCCnsdA4yZ9DKM1c7s1LarZjQFExRh3156MsdK3YvrzQJds85L5Y
DcQqUnde9elvoSMIbqWrhBSnbkPprJEcu0GoXxTVWVJT1bqtFJIxL/K2ywWqMe5ntJUeCGi3XbDW
qqZ5qbiSf5+XWvleFonXxSEgY3C5yrfNM1Z4MmLtvcQnYeNwYnFfaI90CbdF2ktwI48njv8zPiZ2
wAUeDuj5gZ38IeM8NMu4HCto8Pva7FuQIMmHMk8nA8gLjE03qWIJLgR3I+/ApZkD0aUhji1l8QrO
14rQefXBS+kOMDxGuIKJrR+QcuicRx6W6TwlcssvB+ap+THIlDUTfCm9Q9NhMXpNu0s3vgFpOiZ4
YMDBbR3CAV8EPwEec/sszlHaO6DWJ+4N7XBpHVZCqzxpiNyFNzvaQobcQuA+Y5ApFSpP1uYxQth5
iL0XdK07bSSIhz4m/LSF0KVGzYmb1CPp3xvChtuEM9foboqd1F1fAuLl4ToucTNJ2NlYB7A1SH5Q
QJ6UYd8chX208sDLxywnyJP/hEtz5ULfFbRGFwTdO9Wzhx3GBNYE+BM/fBl88bK8gij1PrJD8w3z
0OMbzFYS0Oiu7j9qpKoGtEr4H4GVV8uZfcg5j/Rr5JRaG95s+ttv7+GZRkjW1fULCyD00IG6A3xc
/IMo11KdMdYB0YQnkGQfq4TU54s60J35t5oSyUkRbWWiWnpMcepsnNGw6BA3bet4+WfFfpNEYtLi
XNg3qcvibwYoO15T1yoWYW+F6GYp+vW1afMQVp9Ewonuw89Mppts/2iCr7gBYS+QBCcHHtxB+Zaf
/72t7PbirlAl4pDjwYEd/dFWHxTNLdoMNYEpg5GDtpiD9PHjAWrzlk/+4zNGeIAxYlVeyL/Mbtf/
xN4MmFsg65u7uMeXMI6U/5Cm2rcMi+Re23rJyXIfIfl6zO6wa7g5AJ7gl0Ye06BrfelVv4D9cwAE
UO2FE0c01AtZBpyplkyRm1kc6jChNy9mXzl2UpIiyvmI11AfQgXuLj8pgUxEuE67eDPyPBwlaxLr
pSW/yAt9IphISakZ6op8Wuk9zl4sXF6s+ZfTbxQG48EzQcXrSZeWgsdN6McHy/4uzY8jhcwpZFvD
23j8j9jDHDMH3RHZIzR+NmhmvmPW0NQ35d6Ta/nqojmvI4XiZ3NvBA+8ZRVcJ5WaoDAExC3aMrGK
/Upc4huDIC5WdmltTfJ6NM0x8JzVBXa9rsRTWyBmm3GU5kZb2042QGtFPGlJw7PATG+7jGVyFnEf
9DjFRBUSR8TGAulJgvFovAB2NqLQfgKuLn3tLcPtVA896hcdyn24Q73njiHv3LRQxBJT0H44aAAW
v55ayFc8g/xfaBAo1ZRojwP2xiDLtPbMRELkcBXtfbHRbL/VXObRbwVHGJZszGIXbyWqrPAnR63Q
d2JbmGiXnJcUpM9QWj3r3aRJPpuMCRBgIEp2SuDf3eEoFGKeYmLcDdAhd5VSvXx/YOk6ZvsAc2Zg
T+Ls40FkQZP8wP1s8UJFkqAv403C7wKk4gFtySOLn90o6AefTUzHUvo18zN4fYPfh0Ah62HwoLVW
rk7Y3LPEcGgnojHbcSlBiADiEfGNuSoWzUNyfggAjRFzfMzejBT5HT2ukJlDmjvIgCY0dGwjGarI
kXFu0OZ03YXjzYZuHaPg3rsYXPWg9TXE1F5R63E7iJdL25OmvNPxvrwxhWWvMZHmtui/qE9j9ZdU
Rt5FVWhCoHTXEWtnaqZRRUmvDgDZ6h3MqayDZZgQD5UmJHo1ldpA7fvoJ0iIYdYbKO9mGAlC/C8L
Gnps3ovZRfmcw2pb6m698HR7qasxpmcywd7Wr++anGRbvYP8hNHVtB9dOM9bmwTUk7SmUZMFlBJA
xq0fVHgzFkqeIGrmSaRYaWfq701k0DpTxiBCo6r+THOkyXGY0wxAmb4eu6ftsXxEqGeWdR83twQc
OZ/GohkuNkQlJqHvUyPLNRA4Bxauan7ggLCB3bIxWO5dubWFW9s2sScGCVvqw1wxAJGoEUra/nxq
sgS88quC4IDZGUi/C6/jTh2NO30G46AHYi7feEdOsIOle0mD2FQLzOLXIfv3wZlZC3wnnUBtDcGV
d5SK1ESV5SQ/DvZ6WulOTKgUe4hgR/eEsI21kw8vxYKmfPfo7MKrKsw1Z66tQhw0+5nQZzrZHSYc
LZN20iGQRBHBu+C8jdCD6mU+B4FZ0VoWRZaWKfcRR2OiqZ0lrzCBUT6C6Qv3Ka7AAU/eVj6YQo/J
VgXztNF0zmIF9Lo29ISHlw4y41KQGFnVPr8rHBxlGK7kjIgyb8Y6JOpSE1d88o2o9o6q7i+2GbP3
j1mIZCKZtBY7J8wFJ956n4ZBCXLTzK5LIRPTUGyiJSMDBYoalaNaZhAiasRAp8JzgL5pZ+Ij1xVp
IQBcJ2GvjUNS5goxfBbco7jKF1kBZnkpXq/c3tdzNi8OK0+Dck2+tDAVtnkNM6k3knDCcB355qQQ
e8/fRZnqvcKjk0TtDlqXp8OfqZEhWAOcIXc40KIvUhPC5l6JFDyAdpcw3xMYj5pzrtjLKeGgUGhn
TVDmKLdpRdgPpHHcTf8P5J/HS4VoRzXm6HZZKbG1EE7QRuEjPbeXmS5jD0Z3Y5Y+7z32HF3vPhMW
hpN+XqviebTpqYm+Yfx7rDPgEm3DBgMiVyCtRLT0Np52/m60r2uiq6+uYXGxbCpIsanZPS7vwZlm
pT5U+7UhJljmFTFZEH0AqnagtXj1EdTwP+0xvFc2QYWzixQxQiUiICeqb36WZELrThYD+fXOzTR0
0mcU9LcGaaquqe8obPQ50k8Zg+1uLXmzEuXxsjke1yHPXlmNhBxEQ2Y8/rUjpbufBAy5hdnIOd5z
J3suZwHMolehGqsNtRND1nIvD/230WzrZKS/17zb6IfXwUpWEvg/d9UAhC2LV1hPPTpIoctIfkKp
hcOg8QABGbXa99PmiXA/Ekv5tywwdeo0XqTw5UU4cTPOI5eeUu2F22hHP7PMlf2uP0vP9K4I+8tz
OUvRCiIwiHAwjXVjgBWhBw07ZwlVuvKszn7uh/qpAsf8oa9BWyUstQAAeWoURnNbX4eRAa777Kj1
7OIHvXFZVlr3H0B1VRicJFFsMVyP8L/U5eAgVdhCGtMbe/k/PR0DgYFWaURyjHvlQESr4+zse9oO
QC54Br6Hfd4CeHegiz0TyegbOovWOh89NNgi+IKwdLZJIf2iWyLdDJV9b+lMw+YmPF71QsMuUusq
gFKWC4Q6czs+YBNkoIjrlRS+X/8o2uzsHugHmZXBl7Xib5OP4vAKUxtvt0jUjsj4ofvGHUzXx+Mf
N94zPFfWP1DMcZd25LEJOkNxFVF0tcciMl7BU951n6+QVpjnrkzGJz9PLw8WjJ3W7TBJUy0wIcl7
LXyRN407fxJxfOHIRHN/YkikYWN1MkiV1eFLcGI8QRqCe5w+qopvHm+wjyu9Fm9fp7jz4+zkvkon
CGkpZp23iIUmk2Np8w9TH2v84svH3VgEr8xLJAqRMogCL0wKUzH5TsQ6bMZRLwJcx4/A5JT0U2FF
k90YhCC8d99slbo+97pudh9qDpHSgX6BUEntHL+Q/r5uYzLFZezBdZEuX/OQm2HrbOUXPTuWv1fC
2ySWPf9p9JWPy6Et1de5XV11a6kqys6ACRt5Q/rVQvh+rCnIz3JmhDp28Wu3IXprLP5mu9K3J31J
UcIZC0N3qYjDBIe7JNmYdcdNucsJcgC4D7etKnvxszvtU1BkCXnlfvrjYA3mhUnAL/xuBAerHg5H
bVxpZh+ZaI0kuRi+HToP9L96qEMCuwqyLtJYjvPZVnnnF79kMP6sLWikX6OcHf/Wkq4KPem4dWC9
LKM8BNWRpAr2rA5GgyMvLvntAQkV0EOtr+FLZFdsBVAd2M+UogNZujU8lQjMVeMco+F/s2UBs138
k+bU+HptpWZXQcEOzekhH0OMll0HHHry6kxt1pQ31VrPKE0WIXxs87+72U3CGP0xfWv7FI1t0fGH
mfDx0eIiyMJJ0P5zFvTUbJ6mbiZ3J/oEc6JGHQE3EVog+bQa1fnW05/K2PXHVc2JbRp/HuIhhIN3
tuCaWpV7vTyO7wZDpsHFlCcktKTCFtYk/3foHY429h/N4sDzpVzohXEIAprTPWU/iQJri2EDcN7E
uh6hQx/+R49ukeB5lENRGi84hD2t6HQfkhpo3cNl+ZylvFj2BqsS/9/dHU8/mdTED7ucO2Kfr7xd
u06EvjRsirm5ufZl6UwJGQfmFE4vpZ8+oG4/+GNEFUz3W4c5oLhBHiMgJOdlZeLFofM+axJEke3k
RTjiBGK0yOzoRjo0WEcTDW10ItQ2A/wQ/Ipw5F/KYDeZaG3vA9SCwW7YbavxFr5XY+JXRw6HGPUl
anJ38fbh/iTbwV0eVYLCEIKk/Wm++4YK0PNpCT3CMs5L8LRL+2ARo58uAxEqdnHzKeGrj+kIVyBZ
4GE8d+0mtEvx15kX/juJCgSD0MI1fxFRxdgiZRkxVKLF3yNSqQzfFNhrdKg+NmygaqcQIpLulGbt
o1g1KbP9KIdaAfXL48rOphmdt6EGCUsWf+ipMEeXK7ewnRsUKRXn3hUeLq3RxUe6x3B4tmFu4wUQ
jQxGC6FuxqYFLW1UNnJao+BUxQkx/Q9YcsxuRmoJlZD4q2R8ZF91pwb5y0D96mbNyq3eHdRvYg03
atw+A0fmT8oxkz0F+B16as1w3brQUcBEik4roi3y7Ljiob82NpcZaSFyUefj8TOkoT23put2rRzV
v+f4GgtM+dECqg3/iVD5FTzzuABoAXAcA6Zk/UfxEhxX4TQV67cEQ2XoO2BtDLjk2Fcj8u9r6hu8
OPQKzN1+1ISB2Q1rbWdKxK7GsFtfRjXOWdfXy2YcbpB4qbzhcSxu7y2NSxGq+x0UVFKwjohaDZzL
LluLD75PlDvCVNhpmd5t94y+yCFn9LYEJ3D376GOeWJbJWI5fs0shvgdKvW2Z0ht7rwDtDuJqkF7
Bxl1NP+SfQcEiSJXbM5wQWNjq0CQ7dds9hJfk63LsAeUOQOh/YjIw0HIkiTcs/l56FdHOcYSqEMG
xaNhr6p8LjFk83xJZGaZmyHYrq3Rvz7/U3XI5XC97o1fST2WLg5i65WqHI4Tbek5T5XIEOKbESWC
5OMMQbLuUJWG7PLJDhK8fcf8n9Ypzd3y3sPn4J7xYV9IwUgfciISHZXPmcdFz6+K0kfLd12Er16a
fmAfS8p81eDF0C3idEW33zFpouiHSDtIS0XXCd3iB0d/6hx3sOqJGBMrOpQv7KS71pYL4Vs8w4P8
/cgm2l4Py9igWe6911CSJlYbfcbZox3Qm3cnBBeFN4Jz+8n/fCRzgLRGEooITT1+ytLbBwCOIyRO
OwsT+6PH/rpzrOWYHEJCQYkuwBrAgX5dLl+BCITVZJIVPyXKSksprocJFoWylWF9a98/KKlwPDXu
IWM7cpGlNlb0ER7CIXX/3QAPuRulJBawY6FAQeFfE6OrL8X91ioWKv86O3R5Z7DkK8bgV9f1ZyBV
mqM8nbZp5Q2ZMK+hKoErbDoax3WcO5HLtHWU5hjYEuTDpcLFhllt0/5JCyzEIF7u5ksHElVnmBBC
H4hWAyObA4GlWp7YpDMY1pI83nQY+mgbeb5YSrEh7pz1PU7Q9kpwp5ZS9aZqPMZRYpeN3+yIENct
aQSKbxUKKYBx+Io/woyEz7IJyqxn55MRw6zpboN77VgD+kw4BuNTOaxWzB2+29fsPE9gAvh5Z8wQ
JSS9jL4ulKNkBT/dnzKMEFOn8L6IoXHdSELAwpNsfLsdqKrW+Eg3g1uDtVykg8Qyoqd6MJ5OMV4K
40LodqCW02QIVRt6cqY/T/hjZ4u+O7h/2qJBlrAiVVQpZ4xDZGC6EQfIW+l70jWTcRaoWlt3I3kF
DowuLzNn+rh3R3khujUz4cn41B3ZnHjwvm6aTXiNZl6EXY9rqHYjnZ1zIO6ZlSlC1ddZ67kzRH4p
MNvmGgNYBslG2G5bDOPq1NuvJUVHyq8koHHHKAQIebgqAHFMPVAq03D5kuIPffrR/3QWs1xaoPVr
bG0O8F32hFP3wLgmjcUv6QiEIvJCZj0bQSIgtHkkon2CPKwNJ5FQ0kz8U9FMTR3a3QXGtBg4f9w8
KXqvBvKKvps7f2fnZwmthxalmOGbyoW8JV9EGTmPSijj7yLXQb0+tEjEdjcMBdz3p8e0FdlpJT8q
X9phsII/ZMV1txuqwTCFvA+Swn/mrzfS3uQ8rgHdXjlAD8w4hkuXk2hwe0Eo6k19t4Hr31Zbra88
1znNJ/WHIh/nSXSmy3o1ZqMW9HIaRcB8XDSEURt/tnbOAStlcKlVFc6zfGniyQw7qrKvLk0vzkaK
1s1vURx+mJJFXpcIUddFdvgV6PDwYpTJWvXhxILRF3dyO3No4nzgAoxKJVu3v7WAAiof9tNXbvHQ
HXBCqr5KhXFRfsQ6GNM6WhbJsINSL+k6BM9OX6w45ft5mLK7M4Vi/Ccuxa1yCduZEQOdAlz2XCCQ
HSgxIigPRwUYp2wB5j5cxWqjEf6Xk4Ocpo3aZADheL7JdU3MhO8Ya2dIOWireIInWeJmcALuOuYn
BrFuTpcyopodCNQVWIhYCiMTJyXHeEYercxq3W4jh235yzQtK5oLB7lxgRDx/X/FzEvZDgnlvFqG
iVFGrYn1gowXRg81qcWdvKW/vbWLyxdKKEoDRqH+Z8aCoxuaH4qa9HeiLjTpnS8454e+q2k1ZAzG
nJ58Og+1A6DYA8vN6kxqXr1YroAmg+ADm3a0zKGs6vqdQt4Hhxui/mo15ZZJahR1ZHIDkNjE1O3S
a91a8Z6J51zs0tWcpXA4YevGyOUgJOy4j0KOdlC6sq7HZMqCN11U7ixA48gQbcjd5rJv5JCpSfYs
NIN6YdMRcrrC0n+TH2qOHQocJPeJRGv4+DajkaeJxYutF3DFJa8osZxbeDO/HHnsPRKr3+pUo5IE
orDBDK/AJ5+QWobdjRG5eCnz9OVxPHhH+DXSoWKAiL6PAL9GQ1j2wsslmqEl44S24XYDF0BvZ8cN
itbVp1Q4TEFDpti+CXdm+CETbaVv0Qi6JevDqLqKhXMyRovrdrxVu7qCV6O2QtY3CRMvzJqRmqmL
snLrCeMENpmdBJzKk4f5m1TGYHau4NIX6TQS3f+mw477XWy8mbUEkLsgw6O03t7eAUIWOgAyk+tB
6YF2uLNHa9Bc6UuakA3UO6IU3t5IujtK95/Os4QF/eMXYCqfcfcisdPHVTCmw5Dqqz9RY2+YuIYA
j59V8hDqypNn2gB7Qoydx/02UHTaTK6/mn9YxPeDw+qYwQ6nBbcADZl9O5GYw8Vpcq2IIlaJfsTZ
dLOYiMwk3XOK4wRaY7tCXQ9yf9T5Mrx7ZnAM0JwBWk1MbOEDt/Xf3LEyGpblXSUuaLSY6zEkO3h/
ODP+8QX1cNxBe0j1G0enCJPH6BqJg39joTaAU//bG2sAJB0sYsb1vZpxgev75r0kfEM8b1qWpbQp
t53K+vSb1FvKzS3FFIIG6lTBXzAp7wcPYoQ/2ypdUnFmsCS0bNiAdvCYTq1IkqteM7IBpNV7PkR5
ZAjhak2Ya8HyqnvGEqLK+FbBwVPw1X6b8tJPFkfr/KM/lSJxRVPPS+aXZt1X2rDz3VpMr+946Qta
i6fP2DweHPWE5YpF4540+NtcPg4ThFbH9wNvpIlB+cdaj2Nw7/J7FQ8k1GYsRAf7Eu7yYkaMENGc
u3O9A49OTeQZN4wWMdyt3g3IpLGaPU+pV/glc56grXsHLrA+eKSCcgM95/ShVDZrKY+vayZELvlo
FMZr+tyN7jsFGk6c25rxUczvzwiCuMtaPpHkoupH77lgRjDpFSblxQcS01fieQGpb2+x1z2318Mb
Wt2xc9P5LsDGbQ3xVImayW7EMoUjdeUKonYmBoC7dO/+J8BtwvcapwvTwcQLgNOWfCD2Aw3GVSz/
gh2ltWr5bRoW5/+YWJHfNil8oi7wPrxLD8/9K9W/DTBk33Ey9rWux57tqU4ucwt8eFnESy/BGKf0
r0Tdj9WMtM1IWXpNpQ24+6QGDjcEJlrGmZKMptfigxsrXls3/gAJSv3OABxM1Uf9sOKKRjHvvV/+
dnsgfUh+mqRX3Ntw+hN6geP2qtkwwu43/f0ZpyiI/IgtcB3uTW252bifktLIJoHV/Uxm60IxWHQa
eWLEUA3hLTmI73KM0QIFFuI3v1oTYfkFeYCzeEnLkUEirLbyQhfqsQnEycTc/09WIg+1+Q/w+7HX
uXfbzxQtOhRdVSxsHW7B1plvaWiR1uPI+mgqvEKK8oDbP2yuPnERo9lG59FphenTwuUJ9DBVllS4
AoxP6egK8bV6DThb+0iqJ3VKiSbKgGE6r5ZYDj7IfpUTy+uKJHFIAqd7C3t+maOQ/pb+yHO30KrI
ItGf58LBYn06MaFbHBeq3y7BsltzmN2kqL3c5R8aQYmVkHaF3TFXxZpUjmriOFMuNeKe7GAdP3aP
0JPmQ1DfcIym6oz+D8bA9ktwDxsB09r+4TwgtlbLp+XYEiq1sMeQRYwTSicb0J3NoLewkgaVxin7
xl7JxEG2G66sZILn0/6juvs0szv4WPKL2BD5Msx2LZhfsO2BqLE6E5YEswUaJRM+w5GZo+exEM/1
tovqdgwFmVSEpsuWs1zJs2uQRW2KkX2qM/ysExUV9yOMu9yuu8IRCE0Okvp2iSOPaTwhbGWuT9Az
1zHwgZlAj6/bbXU3D8zkxIn0Hv/uG4mdo4ssUNPK+5yTJIFafV4crnMmxjP/gLlBSliuHnNd52H5
6tc6ckvrOLxzOt1DpIHpplA4vHXd3NdmNHSBpjjckrZ1hfsfH0BU9DaSx6cdeqK9+JB4IWa8gJlq
lzcKPGWJHYLB1YQ0AT3eXpQX9zKi4w4bp9uAo5VduUyjqpL30XHxLOjfMSdJJ65+Jh50f6UqNYn6
Y3JVcbzGiMY1hMhYXo7cxFTIQRoRSYSpZ1IaFxILd3fLJEZU/9rwhNM0sKTp+pKruzQP632ibS9F
JDeup18jaoM3ZiT5IIHhseE2SBlF/Dlkqw6RixJ5oCny1vx7KGnLDdY2u/lpcT6MiN5STJ4kkn/v
030y41sqchsKd28XiioPEUnTFbHWX5K9CRcTYB8O3ucQrWOPIij9pYE9SbhFNhKD89QZF/Nb9urE
Q5Gf3NSPu32P0q+Y47Os9JpDZJL5RpTg35U6wQlVbSErLfgt75k+tq3dJIx2RSzlIQwntPEVnnQa
ouYwVqjxeYRPotCZjmanSFGUA/VuXe1TsjEg74CWym/KgTUdHfQZ7/QvPWchjhqFfNrurljnHMXp
gkURi8vM+7CrNdZmho0xUim7scWerxvzRjE/isQGQ7SzGZjvjETziC6TsImNY1svqnq3djpFGSnu
MTBgGQObdnirnKQYkZ+IVOOya8Z2ue5qGciTomPSkXyWFMZVjT04ab+cmjDI8z6I+6eAjuX4iJ+L
+nT4Cq/moKzfnmFgaUqjdKyuApGR9GQa7rej07qXp0mbznw2pcKUoZIbR/4BSdynu+qx71NjSndS
bRfpnu1pvgkjkGWvwJv/CnM8pXY+gjRKIcqUfJRjH0/txpYNUTo6aqDMVGeMTcZ5qQ9mBRqWZXE1
2BebX4Bu6kfPeYExo7uoFRrUSv47AFpLDDj8/r/BtD+X6qAfBvytlm+gZG4RWaRGNAA12Nbxz7ZD
ubZIWjOE9wmZN8x8AlTutoDCsy/i9onFkSmNh8y/39GrsH2RlZCFsZ+GtrBce/KJhxV1Z7LwvRaJ
BnZInuM0rtme6mTxMZ7j/K+kh3T8XYg5Bem71HCHuwBQIdRvFJ8nyYOte2xwqziIS5UQVWsRJ4zE
dShMzbs1DO4v0HhkVDYth6oSMBaMav/G19tHjSiw/MH9WSppkZcwSl2X6wpthkHcHM95gSeSVlD2
Rnk0oEu+i0TDLvWYqw6BEQ9cJunVARj3itMfTlKUJwaHiMYK81pwWdrxUsYPldIsPe5DAKxEYDRa
vP49zRuNl2xjDm5gndqanzQ00sESiRbs393s6I1i/q5O9n0iPD2uF1jGsem4yL934+CbCNlvzmv0
v0u/JzbfPBLqHukKrKGgxT8ryGpXohCmMajmF/kEBzeBm5uvHwHg0EeKexejqxlcDaX50X26Gdrg
Qnkibabz8pAi7zOVKu6z2oBh0vt380wbEmPa68Ln5XmddhGV3uwBksz6bDV4EgbqrXUWuaAvtJeJ
Ec9lo8zBdtItgVI6Qz+o+UZiI2m+QsWE9UdlsLg0Lhhkplz/IGiBMWEz5MIXS1aavBMYSaXLvYpq
JyLGHHqer0WBHWn6mJT1EJNSJDUYWWMNS5PzjvBia9wl6n6/DF1+TxCxHm+Weh5kkcl5QQBIyZYE
hU3VtEGNYkYvSNaQb5PmzrJmgQd8trgWby2ntnOHJTXR4s9HLa4AEKEz/UiKapl2vY5B6hGohZJ6
lEbL7DXnivoM+eszgNIDX6+kxTl6sERLoGUVmETCDapJMYlysgbvGzIJypmE9leMkOjpWAjyGBqg
g3YczchnYpViuyMLXM/3j7PNd+Wx8p1gnIDe68YGqU2AYdoOaa+1ISQuQLyETq7qd5YGkqNUWgmy
w9WYiEMFk6zsk+VRkSR58rzSQnlFuTvc4pu6KiqcnFwLrOsiqyJk1iq5vgTxAK6JUnVUL+eNAz2u
33Va60uqvGJBKRdEWJtSwyL8PkWzd1kyFPjN4zgPmXSUE4hrCGr++2PRPNLQavzqGH0Z1qHMRYfC
/c4kNAjHnlpnAQJvm77pgALBP5QTCNgt0TDJBVGlCmsuFqOlQ9xUcW4jVvpysuh8YSNOI//EcnCe
GAuRtI0OCtl1Ko/bJSuMksk7Wc3MS603Q8GGbj30WMKUeVcRkwHB8dYX6FmuLj/vGNN/wJrWMshP
rc7vHpxkkfU6cN676BuWQjbTEVn+Rw403w3KSGD8jGq5sjg61RBL2rhoxzEeVkVuC7wXcY+CP/+y
/oLKJlrwTxCurYfv3hLQm+iQs+Z/RKWEPsEwkbJjlhbaD1eAlD2X8XzfccyzJk/C6B8Ib5yRA8K8
YPCuFjYCiIXw+rCT0kKBwiGOCyZGCQ2QOS7VgQTVZn0RKUXmWvZcQEu9IhoF5i39H3UAB843nVSU
g0xJzRdnDoZRNMTY8TwEnUibWHvJ2YDp2oXEIKvFFUdxl5U/iA/kpy6plXlRdOcAiGiwmeiLl+m+
23sfHxf1NNj7+oTSN4oOyc6DIxdqYfQyCzFBYwRwaEAN0LfOPNcvgGgKCTR9IuYFrOZOkaPtz3Z0
3qxPDh3iyimbwGE4XgTlZ3e+4uzUl7un6Q4Gw0+oI/TGppT8iq+Tzi1Vt03pqlz+WiNlGHgMNOWn
Fe6y9+x+gggKVLO+7yOdohx49n+HoaJiy6EolN7O9DHcVDw4jH4da0Mt3NIkdkfxtn0+x9B/+1l1
Y9WkvUzIqmmW9m7FZWiJLdHMJmXYePlLVemR+GwGNvjiSrZicfC32FvJcE0sbB71Qc9zIW5DZGdG
cExjcEg/7LkaWQQGKO+yjdmchSSL4r/cICrgfwquwvAIvQEnnYLYP8xPPc5N8UXSoJ8ALNcGS5UJ
f7jWdw0U8rmLs5xbtd4xTWYURyUXM6gcVbOhrDQMAfD92jsA+Aexwl2zL6u7Jq4Aa56WHypsd4Iz
z08KfMKJXyL6ga9mXm19gerMmz2LvEH1RYfo+aRbIs8tPPZkOoCUJNtCUulVa5YmJBCSdYchoJM1
bYz/YtMR5EbhrLwq2VsAtmGUrHoW1ETF+WKp44khi8iSyNuMwBc55AuDzvwBIEMj4UVK1CZ5l/8W
R8arUmpszD90ltm/Tn9SnKPbHEmogdQ7AT0GsvMU3C+/SFzn6b7DwyxjudI7DzBjN5/C3mzgMOC8
2Mds7ZxUqK2xJowR/nYSqHp5z4rsBwOMSUk4Jhmc7o9fR0ZulR4jyeHvIUICec5OYjLxeQZUKwaB
iKoqZx80u82YhdXCvQRtjor5jonb+WU6rS62Yo0mZWQXSVOVcmBFxm4WWbN6J9q64yxyAFwrFZc3
Vo7JXy3qallcOjVXs44CgUFZzMSrVHSWmUr9eZrreT+mrYxG5IfgV/TH+5/qJiWCozCjL/2EsQ0o
LyzitPeoy/XWpnSEQqaRxiu12x0JwDTrqwBwm0NBbA2kSIlPj5zThethV6lcRu3IubT+PPslqyha
qQ+Ba1lEVY/ihItiZAOm7QVurw5OIu5aztc3K2jJFsy98fnxUuwm0o4bxgFezghiCCNg5sIXlXVB
0pzLl/BvUrewl+1/9fiUlTzrxoFoP78TAxZyaIzsZEPwF2byJi6+yz4TveeE09w0Cv5P0PLvdDAC
EhU9Jqd90TLw6GARWh13ADjzvcHv7XtJ9I6faaGGRqo54CAJ6RAWmEQOKDqWQ0W4YULpfQ3vM9nk
x+VXVkLrfiDl85vvZco9DtyPqR8WAYCwKLBTOTB7X1CPbHxXIW+mxvCmad9+4sn5ZqhTUYF89d3G
bve+jJ9PF63VeWPqoG01AdWtCFNqSO18ZA69rgOhPz6+uxICIRIYaqeJOeD2C/JaroEYqqxM9mr6
D3CFWUnmDsTyuwJ5i0BoJxdnjDEAlGQOmDVuAnfurYTlmybdWqjbpzkpPB/Olj0hKjmQhSc7w00Y
ljFxObbHNwgfkIMiXEBcRJN54/1HvjhEPMV3Oeun2Q0NP5JBiTHRAUdqer9iBoQvBdHElgFgmAE0
J3nNStcZ4xw6293VVU6AeHe6Cf0OsSc3MrULl+FjZf15T35GA5misL26jIILYPZEBSzhcnqg3JGx
O1MG64kj1Sn7fUe0n/37/nNsZToe0xBJxb3E2pz3lgCPEw6B28zDfeCaEKDVDmXvSnhM8+43gqzX
RQDXRWWNdQGPyxb0NFdXc864KJz4cpPJ1JNCRaabdKfDmFzbN6hwf392sopdmqWLtk9SF/P9E59t
nYuve/KqVOyehuTzR98tE4PauSeaiwiJU10tTOxorTrJYGr6ux+neslTPBHUE1+JclKmY6OBOTpt
H7ubm202aiIpOSAVaRTRFK8H1dnUmrLgKIWBbdTqvzEnFevEpL8O1v9D82ij9DgWiSBu+OBIjeUn
sHUz93HqicplDbrINrzlIF8eklYUqfxa9rQSF+TxZT7NSNthEzzIx/WtP5wzSLniZp1N5pp5nfMV
h5GMMpGrgUz5DUVRu8RP4COsb3PixATEOIJ2D9I7JP3qRJmnWzecpearAtheazUTimBXLVWr9XNk
G6I+WWNQlMlI5y4etaDQfdWFhITOM7wsiejUUmfUS8WmNgZyn7r76L/jrITJgFNt8h8ZPBdvYQGM
v438eR2lnhB58/QwCaf1paYEQwaI5ghBmeV2KyDwhfoTHdVspCRi9XFOc3iEKzDsbMJcFEsgmog2
n/dMIRoTtmp5piD3LhWZNqxX69O6ieIkvSe2R+iAMOqGHyivLkmFapWg32zCX42V7kiZQIznVXe3
MQuA91BPIM803PwJR00Ke1RtaMfBFugDPDDbQLu1/vBSedQZIaM/yVy8m5bEJ/gkeobY2Sid/17R
4g9Ksec9pRj1kgQu6SRFkyAmN7r2cezFfmjDDtG6LH0eMsP9jSrO8aImm3PPYFTl7VbEOm/e/dUj
t3g7U+CIKmrXgfW69cJRKCzft5mqzAcoyTpptuJ0eU/F1C7BtvbXSycs1AjIwZLDe3f78/Owxwsb
oamTTKrqeQ1Zxwf8zGfxstYorVy8miDZ7WhFos5VGbxgHJXr5T5j2g0/ZRoX/rLOj6BXGxl0rjMX
9R0OJ2panL7gOvjmifhTjJVKoCCVd2apmuO1KJ4gFCniIA/UoQSxUZldwyvhLaDkqZJLh5Yhuptq
bu5WaHAX1FxWM+LzZRDOle89d/vHEA8KSmQlr77lA4mjPAHj/R8fXUAj+Whbz0Flz8pYGQ2PfljP
DPhGONiu8tnP6XjoG3mciLrExZqzY3M3favXNGNvzWjasWuKyixQHpYW5YykRgY2yPia/lqiQGWJ
SORhircJ395jpqMN33Jw6QtqujZIcSWGgTVclfXy0sl0AmJagrDXfAuhqgmpf9YTcI32IF78XzrA
8oynXi2qJXObzTtGlwMO5mGildRWVYOMRmGQwnkTNW6xMEGigUWUR4O5GRzOLos0lq8Ji8W+c6V1
eQSEyizDq30pQyo9iPUVGpelS9wqRA2kzrtUHOJUQV+Eolxl8WPR3BRVnNT1d4YuScjg7YCZu3M0
fO/DRndyJITpXJJV52y1241ClanqZWto7PMxOfo3UF4DT8v7qOIbn/nGJc+pd7ooUolrR7SX1a8n
Ksrm5Ov1Ebs22E4XbIbBw6MjEGrP7oI06EB1FLwcVwNBHz9hy+RpE443Nx3ChFVmG18uALypISak
uB2bDfxWn4HNNJ0SFqpasNJjlFSdKJcAwq5ifSkRS2IRfNpHnJXffVQ0JhuwsnuYEEbvPdexNoud
m/mDWX32Sbuuw0Kk992CdqRQwHEL2K/Zbmb6J46GwzuiytEYGVvOAXxcL3ZzmmgKKbyo61+P2sgS
JVlm/JjXtGCCwEfFnEeGJY7cQp10gu7w27GwCbQgfIHAoxM9MQQ9/7rO/PsuFL/McTVYLRy2v/BI
2PFB8dZvMqRXEsYPZ6DWZZfWqvcBN2xD/wjWqiOnonDKhdx3WLNjO8KoZsWyQelm6mErCXqY1wjg
RS1Kg8kjKErSwIoPeuVWwyWq7YmoBd0mLVvNKpKAqbt3F5mmA6h/LArMS/oxZeNi8GEkPEqh5odh
cuFF4hvoj96tr6xfOg5EHNlsj3A7h2xT3cFrY7nHe1/IopLBW6kMLJd8o9S2XDfItuzXqi1fQv3f
1eGMRB1Gqsp9D6u+TgQdiGqhQfkGlBFvbdEIEq+w8biHc5QkOLb9xNT44uuczbhgvxKrvLA3ebyg
nXd3EsZWv0NK7+q2zkM+8imxv7Y/OYQS7pWyLXwoLm3XM/XYIdq1ZZI+o0bA0tCtHtDwpMkfyFby
UKuhrknKDfzAWzzs6ZfQiFWzDQNSlulp5S5w/jUQP9PH8CfoaEjrRpjXVKKS1S2zbwj2zAzXBySr
QweLS6+O+vUED82Pldv3YCFJsUCh6n/e0G+St0YHx7DQ/2KPnzOYLFOuG6TCtYQW4onDY810pJKm
owWChh6olAv/zGgJwy/6ckb+CcNLQvWJRtP8DG2sUYsBERn18+H2SsbRpi4aK+EeC8g5qpuwsQ4R
PIzX4qcJOjPbV+Q/Oq66VfkJiOjGq7779Fp1GsdS5GWYGvO4E4fRUbL+lIfpyUmWEZVCavLILvEB
xOfMwYBbgW0iwhjTOGZJphCXpUlINSwY3erot7rW6jyU0/1Ez3kZVihdJ4Pr16sctpywEgr9dtpf
EBuyQSv4UKW0pbXQ/WnS2rEKah1slZWZWOGpBI0OHPLJuLBL6D1qQ2X6o2Mi1+/aCzJ2m8IrUoyY
qoMpa5LITyaJ3wLAXQoGDeE4CsNH6qRikeuG+YZ6rVSXhg4oFDHIWbiIZxhln/C5hwpSowlsnYA4
nPeHNO8b0c/LJVB0L3+ftxXaNEEUKt+yklvWXcYucPPjd3YGh6SihWiQx099+pWuj01TJKcZEOhN
Lj7PHiJ2LwYwW+xa38tV5jc4Uj2B8J3OqQmoyqnweWUeGMk+dHbmh9g/QpMJ2+OotoE8DNrDOi89
vj2WK1AakA+depFGaqVzoxhvuliYB0cZDk0D5sCQj76k9CATiVIc5LlLDPLDJIhq2snh8M4iEsX8
ZjpGaMmHi+CfFs6/MtL+ZqajM6HNnr0x0x+aORZv3KBRLzzyKrQ6x9Plq804JKcY7P1rmbQNfEVu
iH7PAWOvv4AvfLhUF8bLxgj0cH71klghcR3NPccUF7zkrhG6AAHGrcRSzdHd1ltfs0+q4vGwsotX
F/MkNrS5v4sFpXaQvDFlcw9jb304BBN1pQy6FBlkeXXydaE1oN9vgc41SNgKjjXXljbHh3XlpMZy
x6s8n4iuPTVDxDwKi1+vmAFYcsgxFmSjWVmvgbiRGELvtR7ybyAeRtGegZpt1gK9L068uROawGxx
Rjnn9hjfcRAArbT1ELVfz7CrhMEEsUFxD6siwlpgc2RuRh4lzvXQX71D6XpLSGQRAWTkEklh2xtD
sR+KQQX8UyvNjDJSfo6moFMTR7xYktM3Njs9ZG02vDDc0Bpt1CL9VjVMcvDwBk4bUcTxhvbpWAVw
w5Om6o+ZAxYIKc8jxwyfKRW8OFz2+9Y0fnNjHh+oavKkTnPUY8XX/Qg6LVd7jua5UtmS9o7e5qyQ
n0pwActYbTE9SP6B++QbLy48uJXjRl8q79nbnGl2yRde5qzVwX8sek0vflF1IZWiYjZkNerobq9r
qvtxpW0y0CzwFdvDdi+jvA+Dr0BqsqeoaCujIXnpLiw0B3/tGs60s6k1LRmI0iWVz97J1+JnRklL
UmWAs91cUQN4mfTHgH4/lLxPBmiABL2bsgUySNRgdPeYvVXHaRWONyv/d5dCr/KJYvE7DywcUsLW
0dX5gNPzBii2gahSXyJR2gmTobpis+spN4FR4Pp6goHvDv0gtu6hkXAKYaBUXOa5fPWgfH4pmw7r
UfjKWBNgEvBrJAdOPcjiiTnUAUWl2DOPwVy5DFcsSR2SnD+6O2JklWSXmA35Ww6sWAwEBbF38cGE
1cQHQBr/do7fHGvwC2H5Wo8ED1Y8zGHkTKHHFg7dAijlSpvbfnWjRI23k9kWAtUrfy5qtpkyIIY8
Hf9ntop21hH6drsFiP0W6JlaitTrHzB0NMgb7FS3BU66E9nCQ9dKm8RtAsyB4e0OgyOocsNRilZd
juG4BLvUUg7RBM3N/sgwNDvP5mFP8CL1KLm+PX0rDNmXXuYoB11/fAp4/QypuyJUO1Sgdz8Q6Ixs
BS+jZeczVnRGsvCJz/afV8nr5/OFR438+r31piHDkWanbNg9OXznY+DZ1uCReVijVpaJxQ7CQL04
8bVUZxnykTu1+ivsffxJjkWMLqfwzfZIe0uPh770lF5jFlEkEB37SRSpXhQYp18/ryuA0ZB3Fm/e
x2wrdfm16T1owJobMBewgUsSZ0aMMp9Mc3srAWSBoRdIm8rbfK7X9Xl9lpFySunwcOGW5EErqETh
x9p304COJmTQqijgCi1ehfI3q2kU6m0MscNnze/PhIzKjBuQoBw59nmafYQjU/djjUm5KAPDZtud
g/N+TVns+RprC20c1yDONJRIIwxn9IJtb0cDKk0zPETEKDGQHkZ2TfHPloNi4AevGebokwPv9Sla
bkOlIZTLQ1f0EWVHqpx+QLe3IvLmwT1P1Rr1JHHnKp+kf50N8pO7tHAakff+hpo/QdkQ368zKie+
tD12wIbgj9MJBFK61TlrKdWkCXHMmawP42lgf8+IqmbJfEX4MCDuPGGCpl/l5LibV2GthzeZ7KxH
bXYbq/QVt8oJK131vzxhZocd4CgXg22deMWwjWZ9whMi8pz5Yau3qq7RKp7FX4zd0LPz0CfSsYdo
7rJDYRAjxXUBSsfMyReIvXzrnkbEWT1EpkZR4yJ9yA8Ztev7UDL+P1rALi71KGtmb1nrb4zKyHo3
0IaoddX4MEEcM7JUjhLKKyhnZNdpbSncA1QLJkQZV9649jOX6yU26cblS0UUiyLxJIBbiF9mPtWx
de2MR9T8FDUOxOO+ZE3cLI8MeoPApjHXva9b1489Zb9FBD9bLxeemTor8tGqP6F7hdUWAiU/AsMU
34oxkhwUreity8bL4TfstMEkpCIGqJr+xj9NhFFfUab+yr+y/8do//VzUj1ZL66Ba2wxeXQVKQO7
wpaxbuWbdJRxFrHk4m8mx7EbHdDMQhnMq98gvdflIxIxBx/X1slGvjypacV97CO98HJw1FW+3jZV
8XLoHm/dJgch8sQqLRT2d/N6OszSMAdzTgjXthqrnui1gK/IVbg5CTnHU4wq5eNTaR7qqjlXAWbn
WLV++4RcY3TiTxaS9r/P/8HVmAqMHBWTg/ulkIChN1kEh8osMiFC6eogvJTG/DbSH/nnWL2xX76p
UoBkxr5guIvWMSZx3Tt6WXIHaDwDbhtInuxgVj/ZylJbOGa7H5mxLJEclmDzjcXh4B7SKpaGs6J+
VFOo4djKiA7lWxHMp130d1Kyia8E5uXpxgzN13avt5lS6shFctb7xmQ0PfoDrQv8DyS9yFbf6uS3
kIsICmQFvbpyzNeJi09c0n2JfFyEH3W7x4J6H2xS9lTS+f9RD/tgYW4DLnqqNTJ70SKjEWkqBeHB
UoEA49m5OlcuXgk0+mbSrfSFMmFdv9Vry5QWtLSM0GH44PLfISfYud7bsEPTros/xcM/KEnspg9+
mTwlnI9RPzlFurn3+l96m3B6Ltlc80zk8OzuSJwA+s8owl+tWC7SH4ElFaKP0+m75WFbl6cu7Nku
/mFu4a0hrhZrVvgL4vFDmDiviRf0NgdVuvn9eRhdlFOC3+Br29AA6IXlnhyoMlkU5QdTJ7V4e7Cl
yyi4LA/dRO008caOQXBTbJkINyP7WNZYulhMx2Ft1tjyTN4T1TQ5lZ8x4Bj9hachWc18P9wQQ+x7
759ZmrhHzeLv/WKNE43fPK+AQb7vK4CBCoFUJ63sbYH0Y/5StYY+G5YczmO2rTAUQlV4+7pEDfe5
ZyZVJpXvG5yGVi0KiD3UjCNoGECjm4sppqY04XkTc4VspptYBhZV148A4iM/PLIVQsmEuUIi4rJM
dTmyjuSq61WhwKv+hJQKDVjXggbsx3bKr+SvhNtJ3N8SUK8dWEVgkqHUdliRUoQtK06/D0+JO72H
mAjaXSwH7ereyCszWK14n50HolUMc63ztyG8LBIjFOFvxy7a2fbTrldX/h8bx6KmDpVKwr0ZVHxi
jRPUBSnvw93JHn7lB3d+bYQt4mSrq4k5rqox0ZagYvWgX3rjt01tpvw6CKI0Jaahcn5tuZa+h2Gi
niTKUmZ9q8MmcWzwKXxg+unfcxQE+UVPs4bdUPD3U/QnM4m3mAd5ZMISlEqs/SgnGNkHJSXmqoui
JrCGlQzgcfoa0Cw66lC7RBv+WHMLJyPBMTomWMSzpRtUBiQqztvegyMdnThI6nctHFDaw7hhZchc
OICluStrATHY1WdAIUfZ47L7KPGhNHj7nJ/uL6bLZEgkpHK+c9oe3AuwOp3+a5Qo26E6R25Umtym
nwLqJalvH5t6HzR+hMSAnlexcOtYNuXl+gHX+n/EUMwwMj9pC94yHEdSwCV7YqdU05G5q5SQYGza
BZVmUHBjFmamtNOWu/MLw5HXZ3w5j+omEh24sAAKwSLudUbIwQ7xMSH1lh/LSDVqGtuVIvVPGZr7
niVWSZs9Sl/78FvIl1Qks1GtdIxLVvSBH3wY8cF82UAvRbvHMWxHhJ++gGeHdxYoSai7C33AAMyb
/um7Wt0G/NSKIMvT7SOKAHSrzs96tahLGK7/9fSHHSvCpoflgxV4HpQr8xkBL9xwPz2sqzUG+vuj
qvzkdKJE2fLEc7PUhjipLZltiMoTms1p7WbzwakT0GL/ZGVndzMfqzVK41wIo+kvBhB0pZ1LOIRK
oFyihPBCBxEh+Rb40kdnLDZxJVYJE/9JKDuIEo+SYuSrzei2JoL10+AOBxTTC+BwPFNZOxWJVR9D
PaL+502MAOmzL26LHRjJ64PB9pq/HiXJGmQx8p8q6fa/BcliMBgeBiam5Ql63/s7Up+zQrGGEk2P
JRYhRwroZS3KGzJ6fOJOsbpK1v/Px0DzaR+gcQ9KRcYSlldSSJWrfy26/6+K0oO7ldsTGjRy3tY0
bna422BEzplzts0spqWid2H9TLC66ZLUOlqo219trcJ12A76KBZ/nV+/ZFlJCJaU9332t2o9gLJ6
2hQgGNeHURQbDGrZsfDl0OtRDqJi0VwswwH4MRdeNPrq69dt22FHyHUqCO0WWn9e/xR1emvKAObm
ROe9gshVxA28Oz4ySrgQH5u76BzFjcva0hNYsMQ9zRNRjO+rlgFa9X/MrsitkaRYM21lOrvEZCiv
SwYeYqAQLSIVIyZit/LxzxK1y/tzDZjWaIS8+d5ZX5W6+GUIehORqf+DmH5NLYpP/EZH+iBfuC3A
KNIMHozH4hBNagn+W6YKvp5v4QtbRpIOXKHvZIDuKxBO4AdO0/8UbBYBbiRuLfHRx8dgUQDdUTtO
QXc1E3voxIKhqYYUj86wii3VzDUF/5mJ0INIjc8GyOCkyunLDjo9hGnLzztnCPWy1kE5azOaIt+/
ZKc3dviTojEUME729T+Yg2xxRT2MLV6CzyefYkd2Wng1QnTdcVYFj+FmCjy63mI14QcTwBi8o5ah
M125MEWi1ti+LyfEeJNQKi1Nsr+0pelZboo0gSDqPzcy5malu6/mJVw0kzDo3FbpSgFnGaoGN8oM
Dnw+CnHfZ3Rk6VGfCOOpg5lU9irqoz1h+Vb/iCpOkG4sSELwtLon3Z0gku4aMlHs5kVMM/8P5ifX
yaNd8KOXBJb+FVIjAoO2/fX3FaBve+425h93M4p//TnSIP+J3H8NnPeFBIQFnmCgfFPdp+5n7KM2
uxacaGY5vLfA4mXBRj/mV4qpnBKyC8kGB3pH6TmyUCDLR0qjj1RQWuz5VPlPBDl4TYRiUQvBDZbZ
p+MX3tL2ioOYoAwPsps/PAUizhrlJvVG6H5Ur9GAv/nx7b1xNDaKiUa1gjXXsGzzfgWN1NDMfaTO
Tgt4w5yI3jyccl7uYb0BeSCL1pfW42E2SnAdkwvIJ15yU5poGVWimtYshzeTqpEmji078iL6WPsf
2djzFRlVDa5+e0P0g6iOBLst8Ex9On6d2mv7JJuGzBSpG9m93BvAltuyG9HrcAr5Ixlyy4aAzZR5
RmsbmYFEgH4N6g2oeBUke6HVaByyCNbGeP4xy1a0RuGr3sRAZPwrNpxQUsMzNfKJ2pMMDhLCkH/g
4m0hFpFneippsWZhITrRyTXmUTXQK8NsNdAZzVMdfT0ToVPE/3vdHRXSyTiZHBMCAF8TCquPVsZH
rDvUpMEt/smPICbupX0DkfQJ73lDDRyo+Nx17NxvgHocR9ZD567K5JLW+AYSBRG+gAidajiXPQiA
fPl2SPDL/3ZFMIFVqT4r7YYGeuIyz1LakjJGYdw1yalMSDRrtNjjgh8m9JXE5dNKMfHGg9Wo7O2a
efZmV3qQcvywi+6qF+93MgPh+4lLv/J31yGIPAl5+wzfYSGrCcHBOzaxkKQolt8R4krxA+CQFh20
/HrXwm2+QhmEJsSqqqBWeaLbpg/iiasukeTukFxdPExDqQIEfaWiNaUBN6O8zjGTouNpXadum4jq
CHo2yPtItpljQqRD+iZbmhYvvELwueOFjU2eus2/OcHVI3+XpOye5Y7jekABXSjStkQ+72dvYm6P
iTYXhn5X0NPm7rE2Dq0XpUoWONHqRxVEiLc2LXYsj5/bbqv7lGwmUglSFKlCScflDIEqImaRqvqH
u/VTVsvaHk4DXwFfkn6vQC1vT/hpVUaayfWnxTnJGFQYixBN9WANQfGlsR8FCvxMosUSLKo8cuWL
LgaSDZdKW6ZOrYDQ5OEfXalVBiIBJDfQsK1yjoHu+/TW/sk75kHRn6UuHKM1+TprsJgy0RFCUuCl
cyKktfG5LU52PXsRMg9WmbBawMZG0VgJWQtpNGvcMbdFE9t4UamhQMedV0csk4wEj41YcMcdRFk5
GpzIWbJ8JT4tZeyVSFs0XBgYktZRY3f+sG0w9SLmHf8yMZR8Dfp+kAeJn9cMXPqkoRvtL9Uhuw4u
0WCdhUgQwnfC2kISiYnuTmVkh1aMgHJVUzF20vo3W2vdS8LnMWxDFkkWzc8eo8dKxffQDiI+0xqa
uQSrUk9BqFSDOcLcqhjeWaPJW3NxRyvRrR9fVSztLr0GWU5bGKE7WnRlUp2GItYPY5YkrRrdV5Nc
dgL1RMrifYcM9VW3RmOWrwh+r0856p5Zu3ZyL0JQjn9U3LRbxZjv6b33QIJQJaZakuafaSb1Xkyx
+V3Jv/k5G12wKX6vgVu7RWLpJOwcWRzCKKRSoB9cGVK1k9B0TmP1BIqTS0OWZvrju51rB90B86os
hNOtEhh2MD4gm/P0b00mELGYKlRKI5gU7OC2U+C2OgroBlttlvRdHryMm3ZtDED4UeLKTghirvtJ
yrl64QUmVjUowI2TgNp9nZH/ufsiVI4V2djDbWgVW5ywXAqQPXwjEwZ+tvJD+0tKw5JMBbUTrS87
qyyZIjIIQ2MKZWkjSN1Q568d8tKoaSWQOiK7fPwKRpuVfeaSA9SQTHJCVXeN1umCFODU77M3OJOT
sRBiT1gywpTuwSKUmPTighUXgL9FZry4M7muQul3k7kE0D2OOxWpmAWX2mHX9kuD4+FfagGNai5i
uFO2IKbMxNdiVZit9dbRJLjUGQBl4RPihBMRMTPby8EAClgKKkOAlygg4n8oqLkN60XeuA7Y3lpa
sfxOwQF1BcV+LXIa2UWnHHGleNP03UzhRxW2qoK9db2NElVguEhh+lcisenywcdw+SdVw0MI6bqL
HVXKzDAhXoN+PcveoKouRRdqUMNqrNwwlMe4GIbTT/yL1hnUn1CVc5B6p07xqJFZOy4Gkjha5hjQ
eewqXmSEAN5vQWMskVZEBaDdq1qZ10uHEcIfJrRhUxyqRN7uBQ8Mmqc3XZOMyoyA71lUMjiJl76i
e6Or+WV1vUki/z4lzh+iXxzreIK26oVGLGkx2snnv9bbnpeLuEW9nIAsGZQZ703wdobSODjIPL7q
l5d7Otl7U0W5Ipwa4lO6s10eKIKNm/P/8Qb0YUHH5kXDtG/mzKngJ2jW55212aLXF1PhIPTg30G8
jH+wtK4w/TpkNiaXChcLVjJ7DZotLW43L1vs+FefWwZfT8ynTYWFutZ9CNk6SEmDiSSDUMAfmyaq
Ts566hmjWGaOL8xKRi1RcBbd5xUfN3cS65bPtRakmjTbfm6tx2V2Dm/+7i/4n7w3tCArNpDOtWi5
+VW8EdKLcZh9O2xWOiKbDQR3uL2TSOpYj4G1j+neAjI+zuJ4vRaCTGans1JykKu2AR9UZHL52eVS
/tcbvPUxmqOeVVBtYdl7wgcfYG028eEvV4D7nz81c9Rz8xjN1et7YhubtZ9hkWJCrf/wMc2fIl4j
+spnnHm9yN3IHj3AWaAIHy+2F9cKzX6Aw5YEArTAWPkaN7JNmGKAeKAcCUKik0ue1SlPQMocQubm
Z+hmEdkvsYY7VEor+hbDhc3MNQk7E8Y93cJBZRnJSubKPUsm5DTKZxHGsccFoLE8tYb9UkAaeEFE
pkp3rsIKsK2MWLc/KrvWSSJVB7EGFHSz+ZJ80zw0ovliW2JlrCjLDxLN+el4IehCOsr4QC471sE1
ZuAXdGRG8IxagjRVyqZFq65TQM3X6qr7ag9CF8qXkqlxagXBK2BP4/PiFdL59C1LFTW28t+bEaR0
oiBJrjsriEeKFMULq2Q9rcJ2xm1eKIMh1O5h8MLrAesmNLK+sLvGr2lwXD68E59wbdQc85aCMyCi
3qFGJAF+1I9lBRq3QJsOswcMyazFmqiRV+eCrQp/NaQuK1aIc0jCtbpvkzVkdBMfA4MkvTv7DPB7
JgYVSoIeKWRIJQ9/Jb/0oJwz9Lkw4LI5i136jrsq1Xi8WUJFZH23AWMC5ixt2Y4CnSo3l/dcSjXx
I8LH2nj+tQGfVH7KNruCYOT+lsF/3QN0sUbuQ6SaG6Up7Q16V2wfcGZOWtNfsj88gAA/LHllb1zL
quxNbYxXWYf2MRbiTf39IIn1/07U+X5JclsSES5DxS6FIkvTk5v3YsTwQDJohEBWhd/f6/1hcQy1
CPYVNrzdxdtShkG9BnXqcK/legQpp+tEKfkNYl2v8KtbW4SjBINlNHCYX8LH5Brs83/YyVqkyegR
pkcWijCw6d8ep1h8jOE1L3l1LP6KSncUrSRA8xyi0Jlm2+F5Fw0CmVdVS+GFHuDaT8bkS4bZvlGG
CaKGH4fMX++JAm/PMH/LJOU+1Qc6ToDE39SOd75bzm+sg93DCH+uGd8I1LvN9BeQXlCWx85aRdxi
xX1m4zEIg8MB0+8e6pHWPckBVbTuQ0S27MC7Z1kgfKfdl+75f4RA8NxdCrCFecqvLYxVTyyPxwZ2
NNdVpSOjdlwARehgoF+fPsPfeoVBgoe+QMW0DuE53vhdKzCzgRC8p6PBGDsJat5DBp07mbUZM7NV
i7GD+spLBagNyDA6iA8n8mdpK67YOi7mklITwEeP3yl+HEr4luse7a6GzwL7yBlDCY1c5d9f1lBk
sHitzrGtst4VvWSN3CxvZu5KlUGU9dXnVG3bmZX9NX4BTHWkSEkRRsKupO3HL13HYYDI6GxSeOGz
PWISUySwmljK9/w7DtGxStEk5PBC8/ApflDJ57Ske3aYUVjjDLwyiBUKAIYH3y1miNzwzOKOdJNN
UqmYHI1oOpnjNHjfIviB1qtlIoaMlXynobpJlSospjO8UgKj0trZHLuMzwDlLhX8uIj4HI/8Ry1D
vXyBUUHP7lN8RjQxQmBgL4TolhFa5xwb75aOnIIGxLdzVEAwQL9bVKLviSUWYmSWjMNIN5Nwf4ju
aFO11Pcj2sym4y0R2mB9U4Jdg/FryQNnW2ex8kF8UQo+F++eh0Js4G/33NaCVYjMkpy+Qq4jCTGV
i52Kn5s6yqpFmDAzUvPSvlzB2NKyfn5wXlZNtKkGwOWWdLO3HCdAEZ/ZrYx/7y704AwODvngpcq8
oRzQlV6hSiuuNNss/pa6abIiUmjMicwEMsxzFMc6DBGU4fRajAscmeL5XNViO6OmqZeLOfp0yJpo
kvmrN6QKVLjXMZISF8URJWERxFsyD0IwmeXwxKKw2YeBQ+oQQwI5xQQF+Cmtmqs975J6LkKuS78Z
WbH7ewx4dzlA6CCc6k+RWw+c5ufdxZfbK00UJY/UwXk3OVWeJhC/ghuyogu+n36vTN5TkjeGgs1z
VYnCpAcFSD+JWja1eKgnOhYZ+96ePXwKD/u8vfMoq60PkmO3FpUd7FTAEXlbnHiKA/jLcKOAkMJs
YWR4J0gcCXa2ff65hWiRcBKVYefPXLHYpXm6dfRf3qrC8jj/R/GBmNSu7yvR9LwL7zFFYDjnbu63
eKkHO1ILfksdbIU3uUefExae5Eok4sWhnS9bsXa9l2vhZQGKpFt0Bfuk/Mo/2iKE5r+v432GDlsB
JtJ4eNq364k3DTdKaPbRZQzU1yhqbVngFr1TLYBBcaaLAuQ5J2Ybs/rs874n/c3auYVDCllXIRrW
gXGBC6OkWqMwM75lB/hcBLOQOXZ9Woq0XoQUJu6AVwhYlKXysy9r0Mz9c5hHLbQlA7e7duhUgeUh
1QRZ/Y0fv6/Ju2URoUNV2HZCWAjH6Mjeu6vBtYSa4HzBvHiMG4I/pHhYZa8gnxcwnml1Y71FTTEk
+5ql57ShCdmujkIvLOB+OFU7S/GDYR6cAi3vh9U2WJoSMkhudbMbKj11LRg8bF0frquFr0Ry8Jy1
eBq7J5os7POLqP++0wjxWstLOqcsPzMq9dfx0QMMDViHqC2j0KaPhc0+t/O4/AaVqXKkP0XC9JbH
LOpZss0NwydRFChbggqDTqV3NghUEq1aB1bqHdnQsHk3IZiOY1myJsCeGEA0ACNad8TtYCdFDw4u
aQpYxZoXppWs9Rd+/m72riPrH72ajQFskLfDx5faWeo2fqfGHTMTDQcpYPQGUoiw+W0mdvLK7iUu
IMBpQKUc/eRw+XDK7pWeBse2ND8mUchw81umhJlsLZnkc7UjLu3cZ9InvCyc03GxtVokYxBJ5zFX
7wuTG2gA/A+P3MRBFs6aiwZUi2IHlXrBfgRauZFAyyZGJh16wNrQFJMn/oD/emHZUtSJSU8w/8oZ
K0PnTz2OMAtETS3Oq7R4t4hKjhqSlXjmCGD4PpBwoA7jDZBoY7Wfpf3/MPlBtmX4QiHOYVhwYmd1
30FJPAFlQlV2JMRBtziWjf0QtDmPKFAcuUVDmg3q7EfGtQxr8gQ7IJ7H31bjcDtG/qZKP4OMeU8h
dXrpAVbk8Nh25THOSx82rWD5DDh0IHJbWWYUnRhE37POxNafFB1tEVoEBjoVdBM8zEFIXu7Xnb0E
aLQbthcPoHxDKtu2QOcX4WEEAck/5yRgCkK7+kZYg0qzfkQLjqkJED8BxIwWdLODC4bLahedXtw0
9mNa7KiryUNGtgOXB86pGGzzT/y0KQfp7/AOUT9sqTRF6xDuNPHWh0Ba50oMd5pExtVGxXeI4rOj
1a5VZYvnWLwB/JeMKoFgadKSCuj0eI8bwsHYapahB5dDzQTzs3gRI48zCATHTJxZk5fvL4yjSDPy
n482YoX5fohbGn8MT75M/d74hmPvnrkilJx5vo7T37AdfYC7zpVeBbj3Cvtb6aHuu8AislzEobk4
sa8tk0mTfjUA49mbTHH9ef0Odxx9VwmHJT3aJ3kvJYK3oXHqwKIAZj0m8Zlf42TTehIMhrAUZyzj
7B4GAXt60etX5Hw0HaDxFumtxL78FRv93Pqr5OusaySdkoABkuNTj9q+hHbvHNnUVdeXEWuIQTCh
X0Jnbk714yuA/zpS5uGKPrX+DD+qdiQioI8eP18gN7IEa1EXXYRgQ4KxL2Y/SfJePEHW7GH+ML5P
4W0NLzJDDwtrTgUIg9yseiei3CqMFcGti93SG0TPMKoBCqXmkSm7eBMEqLSFf4kc57YOa2vVLP/g
qPvaQj1hyphNfGCfNTt227yQq7ttSrKEbWMKRI/fZqLsbvQ7sMy7Kypy2Uiqnrm+KibRPHwkhFEG
EvZ+IcAYjX51s7TtgS30BcdKAOMrnAtDMiSeSz8RBKy2Y0gg+dfBmqw0izrOyJlj/JEwPF+e6mew
sVLkaFF+xaoV5DITV9o+xrNxpwyrNCh3Hpn+fNb8npNXrcl05vMjvpQwzQZfFi/LvCY8mLqwYaqO
h+UWGowxTaKKzB0dhqyLndgqL7584kLOxvRDIA8u6GIFLOD/aGgGbnEUMzuxtu5/RTXU77GhdrM7
gZta2jX8CgiJSjnVoNXm326NLsPfUsMTHwfd4rxaq3m9WOcQ/UZB5/RKOIbgLG6wOorGk+mAduPK
KPXM5iRm7cNWuKJ1v9GJp1tW7Dpb+rrxfHQVjFDN9erXOj8APTCsylPBpNiLPXke9RSxV8srjt+X
astNP5ZEm7P3gv22AkyaGybecXpYNLgELl/4qr/qfGU3NOApD+cXRIxYs5xI3Z6GvOZbm7jjJXZu
14aT/3wDsH2sNRp55RhUDz28GxwiLlV4ldRE6uUGET+3YaxVIxzMgZ6Jg75310aQZxVfnqP6aGwP
Z9iPNmJYef+fKeNrqf7/GF4/nYGollUKg4B7SDSb9lXprcghn72cvKEKILVEzlRaRhlW8kac/bcV
pvvTi4plBGIHESJJvu32zg3zof28w7Gp437HCAVL/ggVPT0y2nIEbdLOGsIEM/ALzzt5w9Ayo4VH
0DcBJuXNuctvFUUQm9XXmUCOEigOvACVm0GDBDm0NtFqYtgdJBp7VGGZMKvcTWKmG1BjMilP6TKh
YanQ/2R5h0hnJLmYhChDb2VLAhLUMqErIECvLhDWTNUEjxnaIMDKu6LchpejdplXEGEv/xHvtcb8
XViUCcYSUFffzbkt+g1TIAWwenjYhcIthB5BXo//xEqw2YLywxg0S5mXc+YSAuE2aO1wu9wwASIw
cixHF5Xu35FTywwQg7lRPlrZvj6V6FaeM06bkBJSMGUP8tL6a8YPXOTVZNg4ioUgR6R+0Q5Hfkak
bG8Zq0/ZxyQd+kNg116WKzOLK73X79muuTpHg4C0t5Kv1YE+OhAWskPryC+lDaNQCp0ltZnDgGXE
de4+EJpr+bG1GVqS/aAWk0EtCDtV1234vAt7R+0LWumTCLw8kjK4c/4tiyTEQvBklt3mDRUjfHh6
Xo6lT0fMdWnVyQ0uJJA8YbeK/A24Rjqwtm/ibUFbXT78aq1D/j8fKz/VN1ZOJlw/MhD/DxUfK5ZR
7nw5+ehsfT3nGE2DXiQiGOlayr3KAcE7u6j5lpzSJpYK8J3orD6GmW6jIlTXy7YSlBYCpwg9VyYy
BKpH80GbwiKIowejj/NNL9PjE3+KWqT4ZYnlbFGIa/BgKLY2d4NYOjziunjtHR0kFqL8TrxU5h6e
nsOVOliu/3uXxtYP21ppEO43oH4PJLrchRKFOtys1G8oLtHdtIkeu4cBNnNkWBtUsHznQljL7NRX
CdSs+vbopj9dJkKz2dEJRSRZcAvROpapk6ZWTwy9rA97vNoYTfNeISoLWb/f0mgJ2mgaBl932lnJ
p7Qi86PWWEwpY8FBh9Ew2UZKb9vXO9C83j+zjzJ3/BZrNL8wjiucF28okLghTuNnVK/DUtYaCj8v
3WoaE/6CSBhSnVw2ImhWa7sk9dfQtF7pciTJWOXcz6oi1ALYyEc6sM7ex6B15tcGqzh8uA9t6PLv
FZVA6Qluoc1HYEUJejKWMRZaPVxFMoYRtFTsdHBlDxsxeQ4g6kuRzsPJ8ib2JDgKY/VBvsvvwSIT
LlpEgdN8nZcZNVqQ0XLkCUPrXHBc2bzQtO7lEv+2+kfUVyGz1Eg0HVnNuwSGGitWykDlh3ijomB1
zPVFi2wouCJGD5cNxct/cBix/EjyF0lfcq7X2GRRPfGduviEWGHR/cqZkMmqCeERvctofk08vhSv
ntOgXZaKIlOXRyGTleq503DhjPj9Ry86zUyMp4yHO8j291+xm6v4ZNhccbna5vMVMeH46KCvgijl
Kf8HjLl7x4x/B3plEBE3jCYh0GeSb92hfIjjrw3kJrFd3Y21Y9FLi0bLF2x4jzMxjFr9fdqP0VJq
V7XB5kIc05Yv3XEBAKpavwGgyT60BNVRGQDZXOIc+TB+xsryXSg4THqz4sJ7H5IXTDBf9jsMwyuF
gb29Xoy81dV9g2v6M2FvakY6yT8Fh05VuDSc9Axtb7R/uaEEwv5Umt3JTgNZmRFpo2MGNkh9tvjC
UYaqfAIjLMtb8lF0RIC8AmZjsrVYPvzSOyj+WseO4ENL8zrK1pwWp6I5pgYMlFmnxsTXY5qBC0xP
frffT93nXSOH37zHoTi1AcVjM4jz4KrcYXCwawn2TX+FiMWPY7apClPxKAT0UblAvGob22e/FiXx
9AJlRff7ByjV9KMeFgt7/rL3nMsOvcb4J2roNBYsCDjwlDOjyMKycVQAqJmq6i8LJg7YjXoFC3bc
h9tl2ao+Z8700wnYsqdUj0z6WWXiR8GzNUS8niCAW5VyG/dRSR08ORDBGW74KaflkNF1NoBMJbQK
iAYqX/fCHay0vT2pj++LxFHeA39+jXDv7JRHc9DLr3wMOYAhO0IoY9W1TnhEB/X+foz6KyQeyU5s
wrp0411Cza1OZyWCme9K8w6UEhGToM4zaqda2yj434LyAo8sJhW8nZcdkrUb4uVrvsUgOAb7r249
xBt1rYJhbTez2ZjfO9rG6WJHjilvsow9TefULapp1E9D30iH6kSFLT+hpxEi8FKMUB2Jr3/qS6P0
U5VGSfShhBUzPe1RF8Ep5aU+47O9b+hu+lSpp8Aw/bxhNtAfilynPR0QG5B654paHbLHUG/MYAq9
cal/EguzCjn9kbPqfI7lx3IrI9rSrSOpcgXFCalgjxwpMaI31CCJcCmklpPo2N9gKn86lFYRg8Ea
Zx0hyXwl1/30RqQWrKpvx1yEOSfNiYh/Y57RAnDoqD6nTsmzgmqt/E7BNN3bXyzbQyECeJv8CKWg
or07iP8c3TQO0Juamxt09Oy4rb3l+zI/qYW6VJ8hCP5CQZ8spe5NBgTa/d0ZPHShZIMc4NAeB6QD
tNJlYtgfhuSONWVIoAGoMNOVOmud+cNRQwHcTetDnlOvTqbNouu1EDsZh+YFuOTD+6CTW0ehcdOX
eXF8G+up34wCMUCyexgEXwpEjvT6l30LhKtyeUGqLezysuUVpJjlv7en+oXU0Z5gB/31HxWTG0cs
EPDWNrOCJaK6BgDRmAqwEOdZ4d+p3DPOZxo0P0LivLS99MnCTsxYk8Fny+ep0Lux8DL/agItfvXr
qfLndbRD9tjVqxuuNFiSkneWfvIARIJGVWYWanEICLFm7sM4C5Hl6jiMOxb1TxsQeQ0yg2y8IkaI
dZhqJBqQAbMaa1rZjwO2ARWU4lh3EK6FS7shalMqlnmf0Jpb+PU55G4DoxxeHSw8IObOknvvqk/J
cZMQV+uxHiHC/OrqnRMtjGlI/WPZOK7Yiy9N9d42CmoxxdzVmLvFIJNyH590M97WDOHCLYGUkic+
qEkKYFsf7zsMalv/YW6yuxRXXZAaxujbJiDveSBjo6w6Cd/qaI9qqVmbtHsk9sEKVDxwr3e2A1E0
/1qTKh+S15NwqECbLiuKVuBvSW744UcgdBfCxu00gHakQLv42kc7oCc4SF/ukenlxSiEBsx/hK+8
wE7C6KQ1gfIZcXDha8S2S0VW56tLpDxAN+4l3na6+BX+SsrIofbcwcmRnWazG77TC58JlkGI7ju2
iV5I6lMSXEcQDmop5bA9w4O7vjLSVs5SCBFq5190OtM9UEPjy05S5xjhiAvsfAT4VGXcwG1n9WK/
9nzeUrNTYs9W5p1DFnmksIXk70O/Un8/yMXMv339pv11ETZLx6wpdmLsGMANyGeFtB6UFwxo0BkZ
d3oCWCgxTmQdGH9If+Dur59821ZnZB/VL1GXIS4s2AUAsh76WFplLxr7DU0xkowuFo8C65NhAz6w
5SiVAdY+YE0ZcS5jF+2sv/uFIeLAwE+ejhyLckcmZg9FKRbWF48cZTAiXzerfqmN7sUYEztEm9Qw
z9J/w/ZMgHpUwA8agjPRAk4/KB0fpk6Ryez33WwrDt75jj2/XETz0OyTIv3IVo5fK1bpRwIJpmah
RiLmX6QLf/oN5rDLHBSWcyooPJ2S8ghLuodrOsUvzHV573202PJN9p/YJ9Iee5XmuaR+eqvMMvu2
o1ScScB5NGDSX1k4qCWw49nFZcMk8x8D8H2zQBH01pp0N4d9ag3J86c3g6HMGugKYFRPO0qDkNZl
BtEcYibTFloiD7Fz7+4a3GU6DqXIra0CigezG2CwKFyPv2Nyy6Im8K2LIiS6pheZj39+wp65wBEo
NgZz8DTroP6Agqhp+fv9jiBpRhjlXtG3cbMix0vZ+Yr2hI03mA5O/9QJD4so2Hy9QW4D/qVU0l8r
tFEZ+6waZ7TalVH4JSVLWRzWknYLj5y1LhpwKUWjouiuhUeAKJEw/gqeOFG4SJXOEaMQayOhF487
LjHi8BlxaglLfjSlhQbr3q585nKRpXTtKL9oPo3GnISQ3XKAbUvLZ1PdqY+e89YEOg3SW1hndpTu
OBp6Ynq9SFT51HgmUQ77MNajrGJCH05lngDEzDNismS0XeIxhdo30PeQZf5BtQL5c8lyQZyQmc7z
+sYWYpu+z73pRXb/ghbTcqnE40Yeqn7WXw5YAJusT3RQk/RxpW2XUO4Zl2hjDsCzEu/efOqhn3IT
pfmmzi32gsMGR1ArhK2x/7ku86dgrfyr+B2sZunA5D7r3Lt3h3sQkFbKnPumLQncFxTiN5N1+CMw
jJbucqp1fYix6R/MJRbHMMHECnFJ3MEN8lOsjgut5S3PGU3yvd756zQ+waQE0mczw/tomXZEv+3P
A1IsT0e2j9Bh+v/+VtiraobT8RKlSTDXTwb8+XQxv+VySokFo9m9OuDpy0MmpHFZMxDzFt9Irtx0
WO/cev1blyYTc9mEsdPAPUnoojuppzI3J/144szvB6YUiwVzcy8twjOO2EWLmVlAYZ1ghobzrfmJ
WmBxu9zP5ebRDZWWjhAHAkyfXazbKH/kw0zk9nK8OAaZEmieED3etHzc5DM1iGE1BcIL6EySpWRw
u+2tnohAhWNGX//1WkLuYrItb66UGukDWAKsjJDYDwKxKx0XAap29v8SpGj9fjKG/IGnViMMOCQo
Y/7ALRLJyPDG8cK6lU+VK1uqD3VeBLD3t31LPoOfPM20cgR5F633IfA3STUDtZn5yAXzgBPQ0wv+
iqs8bLEpDq9WkiqUfaA/8XW8o4m9mLJ8GkgH8Zi+ZBe6wMwcdI1Ig4lf6yUz3TSXv0obOwMVHZdo
wv8y8315uQFkLaY+1O4llWKYW/BKfkjhQ7PQesbHSVKPTW+DIDX0VAahx5PWJg21SlMPM76XoPu7
oZRoHlbhqYFdO7hRJjunPtrMYhijyrBZ4xiz32w0MXI7s5NiN+iL8B70HueyDNIobOt13s/7sJ/j
pE6naVQB7IOcSrBBaUxGfm/2sKVw8bWwpkZqXOjvEcgZqPr0jGiaQqsFf5LjU21sV0UBzn9Yy6kN
Q0K7KbtnbRTmBXmcYWZr7mOZKdLRDoQtuoqol+c3IBf2/o21xMoD++2zUOJV7f2YNJJ83EPCQ/nO
6c07pyVuXfLCMgbQE7SkbHBoiuv23peBSooB4xu2gCUDPIjnS40vz1xMK+1jFH2pmAweOGg7zhM4
vZZMysaVKeG3S5bAPwcVKnYp1WoW+YTA5yh7pAAlk1IDH7n6S6BcodnFuza9ZnQnMZHoreGBclS1
9RkPYzierDztLExuXQKY1bfRuvHqrJu7goFtoLF+8OIw/Jk8Qvpu4jS3utRsmj3BVyGlzScKU2Vc
FYTwdArd9ob03X7ZNSNFYDQuAQEoLjap3a9P04UA/cEzDQFEV+gsbKabYoKirJf+Zd7sLVhCtUQd
xnDG1YOjdLKOMnJeiL6UDMVGK4EwyjNQzdJKuXCU7Wix2pDb/BFV9OxyHAHCaMPhV9KZjqQ7+CY8
Uxqx08mhgfgAFxKSeRBYiJs0OcpHkab0fKVLtj3lA1vCx30RgkFV2L4pROfl5hVqrfak79x3PPgf
BMGuwvCWXPDpdbZFD1+2VTu5s28vxSeWMvPsnUjd8b5f4a0Fnq2KWoFB6/mAFPQamiHzOxmGtRZu
ik+YT2lVL8n2wPqVQMwMOQ2maZThjJCLhw8V/fTPNXGSFiTEXnos79KzLSHjHzKjlM/CTa8xIwP2
1uRwP6/ZOxwEUfqX8Ml6sWa5bRj+gC2Fq+2wyUZw3B6t3tnQ7gwlYPQmIHGJ1j5WmWpRJFE5tzJ5
N/S/ZPJD+InlEKt1o2HNep3LBCQ8o/3kpIAAqKhcpPzC6x8wf72oHwfxTghcNLupqNb3K6UabEh/
baRrgH1LbBrOubS8NeBHEGNhHQrrpS4FkA4UdaDaI59FfExRwpnxcHKUv5Gzj/6/h5vTw5iqR9RA
YLkTI6SWoOQDDdRls1vXTi20pQX9ajD0UCg59xYid6HZPHIea71q3jF4ygAYbldjN5bNYSqreo2q
fHB9Hka2tCJchNJDePhkPcOvd0ETm3xbA0lNP3lEtF0UG4MH/m0VfLRfYznlAME/e5Gr94JvraPo
/WY5y+gDdT/HOdqx6/hIGGiZus8Ay3GKxIRqt1UpSiVfJzTnGkSxr9UVOnoPIPg2uP1lnxsrLqYT
5AQmDJRJGRbP7Mx9LYyP+sJsn672RgE/3+JpjgGmDhsjxA/nP+TxLk1lpcoGifXGNqs6N0Q7xF6t
Bzq41NPxaSA9PyHm3xJX7eYmdeQTC3n69TJxPztJ/wtgfngtvoNN6hDHVuP4Y8ENa8oQIUF9SlHi
QbcoYLjR2XD2BeAPF8qPwGHLL670gZ/KafPaQ8xKtSNQei8WEsUA38blWPpIu8vhVP3TYc4PxsYc
CVZL69/8ll+bj2PQllVAncpBHEpc6vzHniLmYylwvm+YcMeK7Fa6IX/xnYQ0+7xRyrKE1HpEO/Og
BfmQ6unZu/K60NlL+UPt4onj0RX/dW+thHjC+Q6KdzunsezOPXTn93wLi806kNJPi5GRX1iWUMyG
yqDZnb2KzZ1wEQz0FAYx8pyMOEZS88EyY1YjSmOy3yqFCp40Vl/lgY/ylbY0sJlTVjpy6uMNC0aX
qZGAlI+1hRvIhhrRpt8dkfuv8kTjd0aj7rxRfaPzjDoq3mvl4aDOR0gaQlxhCEkXa+2Yi/6BwwKv
DIuzTtQ6d2dARB8LI02fXtTkL0AsXEX61skZX3po4NHhCkDsNua1XJoFhm3MIWBFgh5wo5Va9VCf
duKT/iML8Da2dZy1SoAoCsbulptSHCx1GKzu4VFGBMY6/kbpmBYX94Icb5jzXSe8sCU9SygF0A9H
dSAfsBokFEJxQ4lJ1wp6lwlTI4z8oBNGWKyKqksySP+CMixW16qQ9qHDTukt5CLcp8q04fYvecZv
9DI7lML49pW6WCH6i3UPmJBlQKrlK4u6WzgQpQVBzWThNumxt51yB45/VIXthBA5gM8eLLukI4dl
axOhMbm6S8cwkeKQE7Ll/cK3sxe58tG1ugCLGKhZHZyWj4f/nitI4N5QPt6BVdmUkr7CeGzObgaQ
4tlGqH1PLF0ZOhLYl0wmXDKO+vxWh00Qk2lBkEd50qRX37/diIcK5tkr+pVDoqx5EEOf/GZJMzxS
hhb0si5zhQQYnLNLcVEHjCndCGlJWqoN/ZZLz4E/IAOaFugQ2p/2NyM+PTQLYXoy8jpT98ztmfc2
uoA/oa3J3KfCuk42s84LBfol2aA1buwzlRCQogUCEONAuid8htZ07/P8UQMrHCwbpHbB8xVaLAs4
mib7zY3DM0BCMXVOXf7S3v+8Fp/c60bqXhGYWI+1v1fPcIKaXUkNkF1pfa2rGiqciHad2/v/YjgE
+/SnvmZGDnLiP5mZKrKZOX7z6Aobj9iJ+eAkEZ+0od4uU3R7WyggwB4299stBZDhM7EXflP/9U06
EiFFSkCEkQ2xvgn7se8b3940WYovS6A8mibd5dpTSEj5AoSveuFkiMPmm8fQvyBj9OF+rxKxSo8a
MAFAja6VT7X1OnXvH29z6Lz8sU6nH4ntadhDCd3k0+oCT6BDUs545Nrvqfn1a+Vl6Lr9Qo19OgZW
mziywtb6FrxBKG24jxNRZAEchw2v2UiXybUkWLdPFk0VzvqbDONqLFiIk3rZtikMp8l5gfNjwOGl
Y/gUt0s4DpVELryt4QPKvDXlVI9f39lrLDTE8RaD4JrGHAxkPqm3oBBbceKOK5FomC5pRQsIoDN9
EydCkdsI80uCErJKBrbXmCrFAcE0x3XdeoJ8vBRuF+rt4FDihoF+QylBZonEO/JW+Fh8qwMyA0Ak
EgUGPk2J8CJRODEgXFG0APwe2dWsparKHlrHWsVRMdXATr0C17omBSo8aOaylGhjZ7OqVVvocY19
RT7ddo5aNFpo7sFWA2L8Xh47olBxY+t2j3yM9tU0Qd2ow4i9zvBFr3TEH7hx+rW2tGeq4wY1Q9Aw
dSdVofh/yFWcvesnC9sBLxss2Bs9sc5O8D2+8m++1oD/B+4HpMY/zJYMHAsvYgP3SxnyNchsXZah
6z0Y/IPYZyX9lfYhHKs9VHDQjuEbST3y2bopsZrj5ow3XHd2M2w5DeJ9hXZsDCqJC0Ti8/Xngjge
upjwvGiBe0FSLUIK0yVo/+OpanuHA0BLxxJJfzzdn+fpZQmcQuH2KYoqrNXN+YZYSC1P7u3mEc0y
umr7mw7A40X4c2mpxlVTfi1wuS4TgMhYdxXwyE9CcvDFphZVpZI8uzUg1A/gEFGkm933KWdHZzk0
TWmPcDELoiHFWTFU8PxA4p3K5yX5gcUXN5g2TyESZ9pJQvbgxZVHjEzPPMMRGR6fqifIMFVqouSw
dfpWmkvk/bs7JZ1GI0JHoU7NtHBfUA/XQIHpRvNjeW7AlkxB2v9eSPvXlV9N5qGxNkMmcmNTDGQn
5ePqz8lMF/nhaSUfEpDa9Lg4FCR8XWf+i9ODK0nnmn1XOuW++J6/x0CvPtw005miam5cz/AzW+XG
7ahBL4bFhyrMzQGuvmcXHyPO6yXyFt4ZnNoOQCPZY/MsljVuCC+CLQNZ5DcPj3YSUOPSdH+OQ0BD
03wgN16l7qqbqSAPaDlaYwk1niypM764gXxTUwRGPWKg9Crgz7Ta7U932HXm9uOG96xozZQ9qgAx
pFnVEuI0AKK/39cYwnyyemwDfCatP/TVyA9SYynDst+ACXYGave7XPhYI2Dsn9WPsUQasEwvdtgn
4Ux3AR9lb+8yo7uiMStYQt9YYwBSTzVyPtxFW2HLUfW7qGgpnSvRzDskboNBDTEvJcNUPSShParv
vDrBKeASLrFmimu6/ZxNlSpkSVn0qUw2D9LwEmVSBYaamAsI6SDt9KTZBWNMgbk95nrPvdLd0mUW
vbWOqf4HBZKXYGPXlXluyONyKNnTM+nBps/yRpqmTNb4PdFerENv09CzzAQ8XgA3W8W1UqMQtyZ/
snm7cuamLQI2cSOpoxWHr+B0GueDRPUd3y2eyu+BBtBzYXuu4eEcIcxxL1EN78KX3bmTkbEj6v9R
slgcsn2wtlbQ80DhfYafetFHiJMyvIuDIXP4uvWEzKNL7rriYlGJt05G357L8klsO4k9SeP784jS
6BSckWggx+7DO156o8pRDjvrqn1MmVm/soThWDAM7wOJx31bocDtovtaWsJDnVb8vEcUpj28153D
JeRolLHQcbESLgKB1MZCuTm7seBgTrKpnESJ6cfsY3ZzyTh5tx3zh+6rA2R7yjxpSTjzAMKqb3j8
yry6leQKw9z30ae9+NFOH5OwcW7t6MSuGO1LMObJcFP9WypfwRGXEOACh1giE8Nl6xxfdwDYVdmm
ZEdBM6KgzQQSopwIOEa3O1XvF8M5u1xHPghMu5cMhjJCt5MtvPxrA5j28hB3upjZmlYEVG9BkGyI
32uSlzQCERuliOahpTJep8F/mQyXxGNf1/yOZ48rSSVrBTwlC7Kh33M96sJjXf02+TWgoqAJ8WJN
w4pjXAiwuhPICYWQHzP8fdkJ47FOl8uwP4m5PDR/KdMEGYEaLjOb9Toezj6d/aH+BW2mtvW6RwFZ
3XIdIyySPK5sVtZeyhTFOkWKbx3aMGlBvX7KGkG8r8URI4H9lVqXDsiJm2njGtINSHoakktRe2Sa
iODrrkDYVh1Orf0t5vTzeb12HPy5oVsAgv+u/Lm1Ifgsjji/qiQ9C71zwTv6uEnbzhsqC73hBGll
q9hbBxH94GpFHVIqxJnUIEG5KtNm0s5xAwgld1XBKb4yCx9VN6LaANKEVRCoXejvUc/mKXiB7q3j
2NX2/GTbYWPd3Xjf/qCoPbEBWLIWB78P3TT7+gVqI6NGdp0ugqWGGXzHDS+ATVpgHUA4WOYaw2pV
5YhdXpNpaigkx0ILTzbA4iXp+GpEteeuyl2sAcDQTtqBG3U5xjlyXYR3zlPk86mypZR4IVMCzjMM
ZYUfaDpJTpZeXuPLPPabtXmm6x7iJRh6rp9EO9EEQer/ixKXd14KfLHWzFeVzpiETwjQ1cOfw6kO
Y+gMSO6eRTYn0MVs9vSO+TrMm87hzKj23iwb32zk6inmtb10/iAOGFpjG1XKZ+DSIQiD7z9Ybn0s
/PJ3GTKZDId/CkKEC0GPt3BKjNq+23nkzaAF7gV7/dZATUHb9UpfkzQ4rXeNokxEz5mI1SdZoaVu
3MJoYaKcWGCgZclLrZ5sA2U4IrtMrzpzbJ6T3MEad3FHNtLCmvWuyzdPaOG41ZbLZnSP9cYMQ0c1
5YfQNUtzWcq9PLgsddfedfwiC4CHa4Ia6lLOh44zfrxsKKdnMYgq7CAVlt/aEcRYUJF9YTTJw+Za
dztddug+V/1/fbLEW/+obIf2AH6NKLHZ/WPEW1C06PZ4jd1NpOXZOTvGBYCxAXXWUoxgnnhBLkEj
T3FC48DfvBHhgeK60ZWoyC6A35FBrwXPGUqRw8FhlLuDVgkVBircAE27wBHR6mC51C6N6TO4rWHb
7O91RJvwN4TW5MOVkGSbelEWohiKnb6CCgbzrOQFVtZhwQ0j4rlXsVLiQchjusphPu9FBLxpq0EI
w/JvLWxvdOhSWS/v7wL4LnMquIa00wov3ovmJCB5n0Xlo3cQKfeeRcWHsLVNd0ECrbrs6dLe2N0u
QVihmrA6/hEzBWgrsVihsKoG2W98PJPjXghKUN8SSuZwJYqMjhy06tKS7aTD92DYIQEoSBv2yYjw
icRwBHbJPw2GnLOpvpTY+TWnM47W1BUfoKugIWzq+Bdah2pAUzxurFppuRZlLaDch9s+pvzaJOnS
zSbUhA/ZEnMm4KSU4J6j5b+xt2G0Y+UkvZwt6XlQ3eZXq+dUwZ0Co0yT4DLD7aE45PeNTXMj52K2
Tc/pHIu/XrPxfA+JbfZ/H2gHC5HReZ6yrCvytR0zQnYM9wX042TQTKsc35nJ37L/dt1N8kAoGDc5
RX6Uh+upeYUPkn0ntFFgs0wYSMV5dHswmDRB2VaxUXcsDSp6MjgKVpT4uoVAJKa4mYkua1kTYhmg
mgesSHW8Xhae2IFgaoBmvaUAFAWK5sOBrnXA+z7PUyBm//1ijgTiAzXBNavMBtCzubp5uBIZf9dv
MR3hAbF8kNgONgCupVPFQT0Nowy/WLyK9Xxo2BasaFc3djGj34aonZMoUhMugsKBSdAMWClPlOOE
HjTwI2eIBpc0SRGYpu5XQmnEnlanllqptjEr6eU5AnLx/gC3YnoHmym/04ONQ9d4QID1aC1TCPBs
mCdbwQhFqJ0vxq/6ZbdyXLrdmMdcY90mHeCbeyTm+RvqKgeYUn3y0NxRcdFqJov3VrXRp6rYVLgp
hHYb0QpRabguYCA2GbZ4cwI3J0ao+ASfapJ2UHa7lpSyvg2dB0ooXQ21Ojr7HqwykxGO0AlGtxdF
ddn6/2n6aIijkdRaTzFWgZhTlrlc4S/u2cShgUgBvXrzmcmO1UGVH/V0HEfcqIOqjr0atlW5qE3E
uqEGfAMqBKhpTr/1ucoltsmxHK3G3EwhBetotl8fwJceX+KlP1FqWpM434oyTE0lV5IOIPs772mC
IGb0Z9zIsKHEwwp1+I1YG/czLRpIhK0mpqwvk9EePKXcPMRzS+Mek6Fc/vhs5d07xmdIii28kDoo
/2S2zeLUe4pBRfpAkIZ93bcPTqLzL+PVjmc7CViCpuGw5/Vb2VuQB7GDN3/ouis2tcUd8tXndf1J
57UajPlu8cBfz3Hf+1ZS5VEG98x6om3mgDRpbxjZ/NDcav6HzBhZ0SuZhqMjT8POHzgPC+zAF9ZR
pxz4w96KGfXkSDnFWS1vsPd7WLS2n+F5AWcnwJYDup0dlJqhWgDskyPb4/jrR3IIb3oMObFT3CER
Oxm9zpJx6MmI/voHLcX0W2h+DdPcDImxlEX6PdPBasYFy0n2Mx/ny3GPe28oWKwhOyRawT5ilG2e
SiPFS3TT7sMdXlBp5JyanpYHiiI80S9pmmDjEUIADM2cKBxXm665j5uUJCFqsOxr67qddw/Hi4Ur
au/FbsRRHdxe4Rd2zd7PJxB2CYtisP2VjjJ1IqyRWrIK/R0pWvoumlrWvpOkrZpE1FuAp0r+BWtu
sSf1uWdxoQkQZ1Benxt5neVudRD3j4H2cX2NKGfXaIqILAovxMN4JuUMM+oa3yL/G+kkELvkJIx3
mlmFcDiJTjes2fzR5sg4NEX0JdYciNBM56iWEg7NjqzBj6gUHqZur30AhMItWfQZ5FLMl3SPJaXf
RvJGVm/Sduw32d7lfBFGmLhliwnSctKHvNZ/SM+/oGG3Bgy476SOM0UVjQPp+bKnr1jSDOOIfCPH
u54EkXuBLOJ6CgqAgEbr1bkBGIlr8pKLHQ+R2WfqT4qbCCcnrRR1p5pgqsku8oz2f5DR8Us70zGl
CwAvA3wU8WOiRGUp2aSbj39Xs54EjpshCob/tflH7f0C0UShIZjB53JiAUP9zZN8Sl4cYEZEGWL7
tvKpMse+sh9DXfnCteNMEsnFChRnms/mmgQpy7PTMaUBmPoAWAuDc/Px4wbMwbcPIPjwyfDISulV
x4esaxLhfh7pzWR1tV+xrRvzIqOGfAH1lr9Au/3qsWT32CkfYxz4UT3cl2ddxMlI1KoCHvw8PdMW
ZlDjK6lmwJEzhaDNo9NKI0UD9eOovb8mVDgqHdAJ5eKCjYXOkRRiaQemQhWTzQ++HnMAanG/sFlf
InPIv06B+VtqgggxAA/PAUcLqj80H8aaf3/H/R5m85zESTh71ld/tJHJp1vS8zFOFJx68+L1vFjY
Dqt/9CmGQAhBRSpny5MRKN6LYAQqtYmO++adLmo79ite9PRsyhhXE/6v8YBlaDpEr7imgC5Qh4nx
CrT69l/9jPFu3OWh6Tk0SVPWgSEBxNp1ukNFKJ/Z/b34hcKk4o8KSyEU6ybX18tZHIuyjfR1qPh5
ZiV/WNaEZTKvlIONetXo4I0N1uu/gD3rjKQ4/Wa2s8Jxr7yBikGO0mJVb0TbTDKAZE2Bx++BEhbQ
lY1CJGO3azNNT/pQR/HXJp+OyW1yEYLhJ3T3Lndn4igVLrtDWJRIiPVDILe0ocmpSBYfjvdoHzHN
JeUKizUqn1C4hbkVjcF+iX8i7sMuIZJHOGzpfEUN4zCs0daltQdgn6AWEYmD3nqZofdpGPtMvn4M
t9s1RZhQiKiYFfzxvlcK5rS2gVnR6LmWlQXEWLWCfBrCuohJmnpNo+voEWzwV3p5wmcil2maU9Xy
LimA0DjJIwMvmxnvDSQ6LzsGl1sKcea/X70y0U5QawOPdZIYB5ojU/zqmZ4/1pDwE4uUpvGsS7tN
EZDmDmIKhjVuSs/dAdqHkfDMrO9VUiYx5cFO988mNCvp8xPj33we8k9mdBWQmJOYQHQN/kypsLO4
pRIhO4wCmZYpmYKuiKD23ClgSJLyUBgIVzv+aZSvC7BtHfxX0RhGxEhuFPYa8efxV2tvtynQTArZ
dIAY3o0lhqDS6ubI2xU6lve1ZBvqDvLwY9qYCdDeu1g1ydsDfW8njvCn3wcU4sNxVMYnunE9AHx+
u/M3rkkinWZXD4Bo/53GqVtUvOcVkHIh5bF93l4zf7+/UbFWjqPbvhp/M4cHuJ0b9wIQAYU97bJB
BH/ui9dlgxX6VNy7jN7WxGjlK5HU23MJISxskhYwpV++8cq2CGtz74PSMidhgLklZDd93TiPCaRY
ADFhKUw0NKsTi0XUDkQHba4TlBdIrf9sW9C+JgZ0L4EkXtgpqAEvFjT1NyYynO+Fh2Pb1rQPi9Nr
/9ON7DMo1gMOfKKYwJKWT0eIS30Nn1Sg8aKTTBN4oIHs8HxE5MkUmBa7zatPq1jEnnkbJIiKXjUJ
NS41weQBDpOTJT5rWycgVHqIdXXNKQhT7hIibWwNpF0HzIwNIvtAQgiCBeaZlgiDZ3zsrh55LTgO
7S5rolBzR/1WyLbttjE4vUeeQ21/Jiy/RaCx9hzE63u+f/yo81ReOi+qHhJVdGPRIcp8EkeYZv/q
XHDztsRXBFplcudbhC10spso8KfN9DSN2F69hr+0qecZhGEHoM5KGST6wQgZQ13o3g68X23sf705
4WKqWUKdh9IHhTmYzXURj5F2sqKe/aOIZ0jln6oq73LhEzoK76hQGSGe50W9JBRICPngaRsgVuOY
K/WIFfNpKL0KUXs2YQhjhQjPwBX1DqpDqqOn+e/sav6YsxeVgxGHoKRXv0kiRNJe5U3dDXVvsG/5
4VNqWzSqHkSiAw1OQ50EdX2gI8BftBhadiWVXW+AiLKuLNRQz6kn1VlqB2QBigEPsKMCq3u/a4b0
LWHZWasPxqYxrfObfAUuE4sOeo4gwcwhTspFDAaV3n/dz+8U5Tq8mBX2LvfF4MWbM1/iK25bYYMP
IO932C1wUHxriCRNkVQvee7111s/bvullMBQsxPizXmFZPD6AI0MNAunjmWeO1noFryor5QkYXD7
fIliq4Xz/jsaQOG7fRn3adwxjCl6bvjNru5D5IaQfqu5G929JagJYmagpHPu31PDiosT4w7Xvvnv
Qc4v+rs5Kqu4y+k3/YOwjxQnNWAdtpZz6HVWQ843WdE//ad8/LawHnCCv3ck82f4PdBMmcJbrCHn
WWViJaIkhcZdx2DyC1QLx49itYf8BtPi/qu84MrhYybucA7P8i7uz3YRVBdOObuQEwxIJ82f/yjx
CsvSHiBs7yhcV604AMpOsOsI06UUuq8tvyIXYp92LLP+aLx6a50eThp8yt2G5b0gA88bspjck4BR
c2SZQBo6ZVpF1DOnDP2mHS8L7SfLlLLtY8N4dIA5vLLl1xkAfeCsgM3bFwRwhmoUorqE9SGOGE1J
PjHsWpp8rvvAgdxaW03egR0BvF73yzM05t96FAMZLXZ1PYf6Vnv5K97sq0SVE7aoAFBqFg62XlIJ
Pwa/kzFhGe5QRmmprJv33fgeHaCZ4XgWF1XzzzP0PkAWlGgycGVgGE/BLVzAOc9n3DCpVyGLqd+p
Ben0r42O5HFzdTX/BjqVmFLukBMWtzh6DZO8S8GP3rohnFddTCHrOiap4AQVz+mTwnG1rExR2kXp
Amh01c3FoGwC62fq+gpmzEQQXv39rzKnHbAqQdWujnYK5EJp6TLSg5nwtqd5T8i2l7uwJpWAPgvO
M46vrhDXeT50s7JDcDgI8N9k708cEpsnt2FepwUY8uTmA7AmUaja3Dj3tKOB9laSHnwJ8xnjfpz6
Oqodf/tnollYzOgsWY9rdwxhaDeRuMp1WNAtRoC42f5b5jLuSlQVf0dtc00JnAYhKqxqMzrX8AQK
TG6vnLNtRow9BHIFTDv9eK/VVOvGLwlOQp1QJScA9LkqDACU2FW+oUErGuLVdfmqDCREsTzwR+28
UIyV8Uu5lsyQNdWqAnBNuauu+1xN+XFhAspfrQOd0oN98wbiquIQx53XQ98nbwWD18XX0AK7n/Qq
wQRAA6dM9NQDe0FtDoXmC3TIjTswEVqKaxrICRTAOM2TQFAFPV46sAf6+yUY9DUqRIOz7b0M39cB
vb9PeStaw9+2tKgHkOBdUT22rB1G8SJeqrGES9xZDLShFua7TJz3tpVKnPKk0c2kxSVmidW443DP
F0RdDV0f/0zvPqubKn27uR0zIJbGfmQCBEu0dDfHIh+YBFHab1RU23uDJgDTVp0ZBFwhx3FQky8c
pXHV2acZeiEMaT2vUbBzKVGmSpz5lveSC/64vonT0wEZTVqvKRuNqRSqw604/bP0PZoilFjgX69E
KW20XK8AuiVDGlD73ggs/dQsiGyMkoYGipyGd9wjCNNAe6a74IxGEq+fclm+eEpf734MNENqTvQB
racRSmXpTqdfwdsAcA+hAZJv0plMV006WoLWYDaXK2KkLG7OQhKpDaouILo36cuiMWDYN3mn8Jih
qt9d9REXqb2WhJ4NH1G/VXvZ/ewwe7NLk0HDWkSFqfesk4Bry/8eYG+20m2E0hpmgF6BHZBjLlVV
aZ1BE2ObZtuZEThOQy+/+Eh3p4iIpjawP2ydysJJ5+UB/5SopoTob3DQ4clRNhOVqlSZISrXo1uh
7sN0U4c94IUhjk1Hy7gikErwlzFcKt85DpbxDPX/wHN13NuAZYXhHjAUdK1E9P8twKLMgai2l26X
Y/NPFb677CEL9iTPukJy+Y1y8SAeNtjobiK/gWbTePx9iQ9Jau13S+hVI8ARpjnjzgPVC79/kaP+
0r3KHdhYNvptoy94FB/mudbOwwvlurAlsk9Vz58UkU6F4SYAaYKLAX6LaOx8f6/lMtw8dvklKvej
AlRJVXAo7gjByuIFBxJ3ZLdeg0wlkbMxrHrooji022o0MtPbyVHDqxXJ0lMDELvLBGgvmkQbWSvs
NM61MKM760RhqAirK2llnkM69/tjbNXxnfVDamOZ6ly/mOmhzRDYhGHDJxeoqCzuDHAR0baFk8wv
gG8HyKsOrQ4Zf5S66gRHhK51O9KC5dsyAge6RESqel3uq1iiNz19NKHf5ufQwWb5FIZDk/jvZLhw
Pjqt1x3TgP3uN6LZ0+WodAyyvU9mSJF8gD+5vsyhaIwpuzuXl0UI/s75+XwA5wiyJ0Cm7ZHM/f6g
jTTvbge0B9FUbTfmqN/1a29nhmYwkb8muElBcbefrCe80Czx0WJVEuprqwg9DtbRFRFKMJVB37Q0
K6oQESn6O7hcUVvM+zO6f5E8DRdpIyRDKpOp6wVwqW39WZEhnuT7ifblXYKBuCSLlHs2V1a1CqdZ
mwQqz2lELre4efB2zgXD1BuDy6bPBNbYnXS9hUwS+icVh7aduMWdfDNQhq5jfHSBqZPGkzBsVFGO
M/d9TZnS27qN24NDWL7mlMWSO4K4w3b51GHTFv+XdYY3R9HA3zQRFiL8shMbSYgzVgbYU4j5ejz1
m4y4yjfmPHabyD/7Rql6zYYYEpUpYEjOl3Ae97ssYYFki+Rr44d5MjhpLq6+Pg2eqtJZYLGaRGFS
865mMSSZJOJzaIINzHPLu0+f9Sw4XoNfUoOIzSvIP5S1YeuGxsa3V4QZUcvednexbZ/knGKQzsNU
gUiE5B2bQMgXfJM7HGEBK1AELbdLQOZJLKte+jezshaOg+4q57Alw2tMWP9uLfbbgX1POjS3stoN
TDrhKEqXcHgN0NT+7zkdV6AWTPqbTl9djOvogjCGgX2a1FVIhq5TQIQsTqD5+KfJjInjrOW3eQlt
P6n/35YHrW+xhdyX4HorkpK/wcTyEKjmTuNwgxbWzxM5+4BbxQ1bQgecOV5jl+L8r5ddBDGPPhG1
VxJP3PkX+EIKeStaGVcqMf3Ney1g01hZ5JmUgPRWrMvW9d51Q1pgvqaULgoGaD5axHkAsBkF0GwA
X16/KaLmC+In8t9AXMMP29M2jiJhMnwGE8duca7VDjhB6J1kt7vAZgrlCHZmMNeV7Y0qlwKt4k/R
mBzNYQo/WVI/kByVwzRfdCamw3bN7nlfdzXUwZuuJK1uXPRwpko8dSaud88BGDi4oT1aDMx4dASi
VflyaQ+kM7hO0Bw7r7DgupwpyMadGswJIJArjuGOsYxzGeu2TfYuZ1gL61vp0T0OmHzCgEzc++Ox
3HCGXKB+SLcNOMnc68AS0jjsIEe36wtQygK0jyq4hgoPiq9naTFm65PA9rI9rDbKkO36HpVQTyre
adiIeDYCYQsOEMuTi7bAilruE2GE4db93+PEcCtKMWJXr26lFsUsMWUNdyF1vMKJiPSQaMEYdAze
jaxJsD80PmeBDJRl8wnRePzWX8D/4Y5y3wGzR/U53NxvNXRJQIjfWC4mTGJqTwKjJwcefGubRwCx
B6Y6XZkd39+Mg8+MFavfeFENC7A8u/Q9up0/Xih0pnBlbHkKXqVRyGL3tlFqPVV87DAm/+3OjJ0s
ex4azfEPWojJKR+2kZS3Fp856EW5eDF6igaKtzd8D8w+NG5n6ci/vl8JnBt7h3u3GN0J2DlWILDn
y/ePakQynCEDw4tGP/aAkhn517PKBJkNjXkSMRWlZ+o6qj9a7ML2ck9cY0Pbj3ISVK6dYBkVXi5E
+OLWf4u2omMv2N1pUywzFlGX3XjkDk7+jOU+xPqPMqc4z4D4Gxox54jW/yxg0uuC7KBDKq3aQjcr
b3LzEOeXMH0guyaJMf+9NQHPlhhOW1ugBiAGxXPs4MxVpLPBAB1QLGakvNDha+pOYFRHDbtG3ybH
hsT/+l22nLPWbuQ6wKWpRHzzIM5EbGy4NuavpNEYVi/H24rtkG+NURkOjBA9hTyyFXczUuS+tMoa
Ta/1TmNE+hQB4ImWeSqQda459ARdAB6GXSyP+4++kLaVAu0GuD+HzMGvTgvYev0v/ola9VpZt9kM
uMQt3XMRLx5m5ocrM4fT5KsMzLaqqF9TPQdZudo213OVVG4ndkldz6J6ozA0pxUUcKuOzmdUooOT
VUFylLgd3+/5RIrsK/Mwe1siVYgIrp21xKAnPShYsAsjqOSKLVDnb+reHR6X31lmnz2ZxjrjFUEq
ZKGeqZ0Vd82X3zHNpObQvkxGutJ74msSvABDUsO6nV8L6VrYp+cEq/tBLoYYdLk9nrLEqROdnDEb
CV8vK++onvYWDVvWY9vqIX1l1K2uv1+FyrK3mvvVEHUF+GeyQGGV6YsM1Cew49FvGo8BVVDgv8BQ
6ldFfLtafz565iyb6L6Gh+3iVHqCiLaFXeF3L6UglY4wp/15Up+lY7SYCPP9v30c5qInuozxzYmN
TIEvxPjCVetCut4ujFeQcC3z22ZdgylHHqpyd3R9iqQloA30kpqbtVfiWDtN9vySO4cQ5HNrb718
32S+/x/jM8ijWQJhS9jJPHY8nOWau/LSbRjnJsb9YSE+fW61lW/ArD1/BFhXFpeq5I32qi7q0itZ
RBmYlEKYgfQwyouBxWIXUd1zxa6UWIB5v9OhXCHrJSRV/VWDHyzaYdWJqJeiPyyhYsBT4j3Hfof0
Ypk9K3D3pkN7yK681PBosRDEmoChVD23dhJubp050S5jPxwGakieu33A9bPW1giZZjMA3nCoW+mt
UY5QGdiOUhAy0+YBIvzi0r81EnF4MHK8M5JWOyVDNP5oxZVtlpPs47mnJyZ5/7wFQXXyLuIOMm7H
pzfIP4qpB3qL+8e8QZCINaPmnKz27wq9Wo1QnDipf8MJs3Y7e1NJOCzMh0aiMHfawraDtma/25CD
k/R9Pd/iYAi+60yybjZiywrfG4QqOn+g/ATE+UMQYsERwWv1bSGlKK7abM2smii+LhODF1zdcLen
THoYBV1dhigjgVQHpUa9qUXiVcjDCB4v5PCoGapmA+s+4RKXHuz1GFBdEzS1zWudTYpSB/CAq1ej
JPu4evxWREAynVqIj6hZGQKdrLyCTV9Zahv/UFMt0HHtHDO4hl1jnDgLs3t71POMmRlxCvuUabVd
owEeLvWAF3H5TxyzJ+5Eslz9d3x5mGjYoVFEDGIN2ZYiRfzUGEuLIPvgwPlqwZSoyKxc4H+G/YoA
RJwFkS2npDdZviNgOq9FmY9zk3U6lQo7OEbS9w/1WR7mngjmwx29pWpC8Wv5v9ex6Ii8rzDeig0O
TrpF/M2UVxCUJLG9lzmGV0H8MPktv3TnPrYEoZGblACs/yd7G8XDZkIIa0zDgBRGH/4XIrA2+/lS
5sQlljoy1LZDLKnhDgh9y7+HmQeX+vS/uP7CmVcd3YunRN30LOfglt4P7kPn3xUl+URaKODGRUHg
TG35A3AiWdxGZ9TGzm43T9KJ+8aCluBrI2dz9Xcg1Wsk3MXV6c5sR31c0Vs3jed3sz5CmjEOiYzz
Yh8yPeW7Ubzy/FpT67CXbNJubp8wfGEKmR4rpyO2LEytArRNqdN656BX4RhoEGXWskbXszdFNEfi
Sz5Yt43MaixIt0CYtd91SBeCGq4wX6nFL0O2CxPhqI2ZPJby5lPko2TTND8oA/6wcf16+1gSKb5W
7rDUIqVIlX2mgAxTcTFEJzqkSfazcoUTu9yZb+q2QNoYK5vBImavHeRmyfNX7n1upGKXHr0RXN2y
sA+FYM2PVsZvPZCv+9kWyTqBadUah4Xo82aFTH3i8LYWvyHFM5ASaE5oPlHCbce89fFB816R90Tl
kHIa163PDd/MCq/nGjkcnGNt2bHLfcYNN1L2SyExAyM4D3QfUD4pmPWMsNpHV79oIP7crrnTBq+M
njld7EsQOkuLCpGZgashko/CJxmmzRxQIQzWDUeDJlVkYT9Mdw5B4hvAKOVV02Yo6rQqIHZnKoju
KfhgsaDxDIFg4i99/t+UBxqmJ00SEUDYx3rfy5x1CMpcPsbflzIKuH2pYMMr+e35zoRantyQ9z+O
i11tjpe9LOhkuMRyt9WcotoLYyw5/to+AoEEDLvwDIl2cvITyaEjdxUHFB9DkM99pRIveeIRkuBm
0qYBOeVDMh5GeaC8Oyj1pw1li6FiZJJyoGN0ATgX/KTTp1TCF28NS3dxpS3fewiRXTCoJ9ZtzOkd
tCyB8QYWlY1HmJe7uwTsziDW0jMLJ8hLeIr5r1eDy3kmCzq2lyIY4LR5WEEXxzoiEWW48trppfNl
Xo5npHSaKLzUGk+7I4dawn2zBlV9WuLT+mVWCPfHIJJTvBzLdZxfV4e0HVYUYqPElkaWBcPHqH2S
OIl45vSr/VbjDt/Y3M1Uj9YnqZiEfjP+b7QbkP55AsKuOUbjf97L+cYzzP3UBoBsrEPnBLvtpivJ
hFtm1qwZq1bkiGS9qzOutOBQMEX9bt7OrEYcY06JW+JIzgECIFLqc6d7OqtGdJqaG2g3LV0w5tey
ExEYfCvb98wDJQr0dcJ6lflNzs8BgeV5k1COCfDn72TqfR7a8/BCrzbaMJFc6RzW0Y9pWiH/+lfL
TeIfszQelX+fABY9CL9o46gKBI3YcW+NgY4ZF012ocgB8sybaqlUWfSqvw9GIjwSwCyf4OxHdQfx
ALCrClCMiWjAcs2sIYB5FVc0G+SQFaRYsALHynS+BRXbZypoVeAhWKQDhB6uFKwce0mJWB9CaeoS
/B6Fa/OFuCRdhRGy+gK2/ufZ6t60WYJXeiWKn8Zf5qv50buUyJzk5rQdMWDeQwZjdhUycwPo9XaJ
C/61obHjdrNfLdAXwytzpbii5pP8qNgs8+ZeiXsNUmGYRro5+uuwaNxMuCcdfIKVvMYu4thLyuy9
GtgmM7bvFWIKKqw5j6IVp/aexSDYqL9UZeRWKrJatMlnmzSFcnPgGMy++2CgZ5j3fKwIzk127GKm
Vq3Ebt+/H5/VEKpmXdkAaRcxOT1/yLF9LzF9FG5Gg5gJ1zfpq665TIAs2u+z3w0Ghu8mVS7NUxp0
95+Frsjulzjhkk/P+zwqaMGrwDesbbpk0mco9SdrjClGdVG6FurAwOg9ub436PgWryCf+cxgCr/9
dTH5YTC1n6XP1v8Os+vwzc/IZgnNLO+oPKfg8eY6xxQNuxlbFr/TO1h/r2UOHWwcbXM3u/KF3lf9
K+clRpRdNx/FY4PQOg7icJJdhRTOMo+lBKjrI86e6M+49+tYDFUyHHByDotrRn6EOT5WZL3XIUnA
1qkhn3mej34ZDwgGQeWf2BJBHaW5pIiGySOVGvGcaDm8d4AISm1svYXZgQ0tqC043zNbcezk6D3R
VWZDOgUCmz2+qtzY6pLKghUUndmHVS3s6TU35GZYBwJZKfo5LDkk3664VmQTSQyldORpFxbhE2dl
OPyArr4eznhduFvHvpO9DgEa3pP3Wu89su7vb5OQxOiGrmiJexcIk5enQjZqpuIfLICxQx1uzmkk
AWTUfiWxZLIsGHoj4Di8we+COJwROSbmZIdoOy892Wg1hB9pEgZxC+zmGKjWPeeDRachGHSQxm8g
allLI9wHOGBIVylAKQ9s4gvVtePKhx21Ef/s84grroYTwgW17VwDeiHSMxXM2ziTxogqSKN0iLsC
0NILaejPBtMDsnLl6ok/OIAswRDARFdQGlB1TRhWB/80xeziv2Qb0sMXPK2U9CNIdqAx38maaANP
xlNxejw326zEnpVkx06vJtNvJS2fnOUuWGqmAbzqoOMY65PgZzM+5Wcw3eBKOqV8SKs+8lCkBT83
5HzZrpUBYZ0laqmn1dH6MbKRDbSXJBj5g0DG8+3NdlJ7Vfqu5kOuskQEbSnO6zhzgKsVc6DVyYZ5
pVYspiQcQS/GS0q50uiUiePWm1gTakDSlQj8JjUoE3R8gjb3f/tRQhpIxsGDDtbk9Ng9N2vf9Y8F
tdElwfk79gwKLOaOiPw168MA4XQZWdYpQBTW/WdWBA3fJ8SGKlz3djRbN75qFPpilOP8dbhF4wXx
qsmFp9ad7vyt27iQERwmiOnpXKrrHl069uO1HaRBQ3K3z3uu0AmPnZK58LaTDBlTESj02qUX5OYn
2OIJ+GLQEZyaVuUT//U0iiGOQ+W2YRm8vETCQgGraTmygECXLfeEo6VwK1pVA3Fa6ap5VRiPufxt
h5h6fW4UYxK/i9ijnn/KWTuJdmitaKr23UHTFIfwhiHmHDQ+r1QeBFxKtyNOgACBbZAVur0wl9Xl
K4WooAC0ODVwCvKFuFGm17f15JE2W9z1MSjgYMavOwBcYH/IePCxHZAb6KBFkaXSVPVu2gjbrecS
wuMlpFGqDn2xlgzSMSfO5h3A/KkSXp0P+r4o2XALw0xGCwhZkHA2RlN9q8V8a28SON3oK5qiWsPx
I1nmLCVlUHOAb1T9sYtbHkB13uFMs58Ntg4QPjtCNlESv/69P6hIfUjoXVFQJx4L5KgFBIQTMi3C
38KYD4F1vsLsjdC1Tovllm8s3Szesu61bg4IkpqwwQMA6R6Tz2FsOZl0g9pt2qOtgdUryh3vtD2H
DbXbALcsoR5W1HHOoUCuF6IEI6LZ8HoEgCDUaFtLvXJ41oStLmFiqb9v4oLu3FT+s1TqFSGv+yqZ
Z+BsJlgJI3HIt4EMG6+x26Ndl0RoYTAmcBYj4gP2hB/5gvzP7w85jDUfi+FX+ktZeXax0srB9oR5
1XD9jr1lMubomnfN9KM8UJ09RrzHvGQB5+/iSNwe9HxPt5DsqiLiGkLHDN7A5CkljIkF8uE9Mi0n
3luX7PsoXhTE6IcZ8KMWtKpk5Bx76vB1fcD3Nckoa5+um7nT05tEvDjLx5Ly044dnP5pYAiN6Dr4
pZECRpu9cHnbr3FdbU91qRin2ebabCOhOMtQpe77RetQVDamb78pIMeNH90ZLLqFfVySLglIHLKX
+YHh5oK3moHtsgF4XmV8qrRODNAVZ9d+CHV2XgfkudeVAOivI/QTVmTuJuVG9ORdQaw5op02QhLv
QF9QiZV7Mae47P/1Sn7nbZnX57fvFRme8Yg462tMXM4SN+Mx/3uw9ctosGjsqXbrOCH7ah1pl08D
6uMRQab6EBUF7b3LteGH1bJSPvdXNc8TRpWlv80PPlCIkXU2MlrL0fUSp2F+vShZTjrtqgh+neoR
i9nPrR6TDOJKcUfwuKY256z/DOSlIwC0qONglljEk0quXXb9vHvTpx3lsc9/RzGEne5WOAlLAbmJ
0F59G3ZrJvFCbrhUb7jDTc9AuSZeKP4OPp3UeMubnb0kecQCB7FN+VJusiUifqRHivnWUCemzYuR
M6sKG1Z+XzkV9dsmZRG3ebfw0TaZo/7PwnCMbCkdC4359ulkUNEQxMZh55ol8FRL67eQhHtgDen2
mE/mqftCWuNR3CSdjGYWrKTc3FxTBYB6WTGs35PWW4nBZord58/OO/YJA2h1CPWUIAra+D5WzpHw
r/nyoe+TpD/uTeY5wv+WnRMtRTDCoDQQ4UIlYc84R6GnoBdFPniVwFYsOiNp3NQpF1rYAdqKvscL
BqG2F8GkBtVk57C/zcGCYbzsrfUuQW2GvmwDM8/onwdXRfbw2WCXy2yr+BLbeaY+5OeGMmqn5blD
UrlSCUAo5uvvSO5xmYul22HagZc0qHNF3+FVtLWkWeWbmKo7WPx8+QlcQgHQLkEOS0/uirvvET58
Gzxm/EfwpLramRw1aDe8u38JrFzKzl4nG3pJaAOR2ni4w/VXwJVjZWOO+7yiUTajs9kGmun6aCid
deWmklQqz311blpn7fn5pCOcCm0UUjIDGMVsWu998NyX7xDC06mi+wQbByngFMS9UaocvGnJs1/K
qO5Xi7SDfyavp1jxG1gpjOmiv0LRJc9NbrhmYKbgVW5Z4AwDM+ZXu41NeKnzY4c1B//ic2bEdBT6
WT/kfJpP9aDZps2wsUGSJ9eI5u37RC6YhVwGhLQ3kQDZdLglj0glz6NpL1jrkPaACPyRaSOEQwej
xRxSxJGyahDU4fkGKo7PoEQZM0bKhI2DR3mohLMhJT7V3vzCFK5IDkBWN2xLjx1gsrLIW0k+poTu
+Zy7kUw9XMAZKHQSX1LTk4Gm7JQ/bQj/M/pAPYwV6VfM+3ANprIWmeMYG+KJbZxhGYAJFQMkVJrC
b7PWsXHO5KAfIE/hF/ZZxqB/5AFBJZufHAP7b1HTAzfAFxGMWkG4t7ikhfPN8HXObzBbXU57dPsh
iBt9IcbGwv4GNMGfJby82PPERVvkuWDvjzuIxYMCGhTKGbrN/7i/kde4eChH99/mZVxBo9cUhltU
nYot294u1sgDOnAsIoyuvXfs1m0/TDZ439o8IK94oKtcEVRGrJ9umnPA7FSwhKuWsFRDv0RC6ogg
uTNQ6K1lxn85Gt71NCQlmBPgLZKPNkwkIpCjE9+bzT+F0LQ1vVQt4AIp/D4mUu9VKkgCo8nhwHEc
XpPp5zb53+ixb22mCPTVLEsJMlTrhiNA9D9WBenlTeZqq7a2evIiP7YJJ8zsK3KcxixJibTqlkCE
9ps9sJ+wHYDKF2jdFpvpgfe1PzGNwXyL1TbIqxq+tzuorA2rcU3EBYD51AR82KYNZMwFXPyMukEj
vKMajzJAfnoR7qIhBmqVablbjuWYf09ZL993NETCoVkwe/0085sMUfw4EsW91sIkyfushzmYIvPA
f1im9GFK2PEyjvJEA15CV6SlUM9X0IGX/7fEo88txKBb0Z6Dm4tlPXxEvGMZDrEiy4SxfoASK++P
pigKBiGiiSJWYqQlm/zOOECr2+KrchhRktW0CbVjViaiKY5l812/h9tuoS4Xhg4IbBOzlXJ1w761
1HvQFMjSUidP/VVnJvurH9eQC5ksOj4biSqesQu2Y7n2Pz4uGitDx04Hyk5AjKGSt70BqXYGuPj5
xQ/EdgJNG02DnF1XS9qPoPNxO/TOaUt7nW+e1yIyq/QIreoRVRg0GLA3eijTPsgSWA+gAD3DAKt+
4+Qs1XFQDWIWaigTq1Cjiv2+YQ0wSfaABgOB3j3EY0Zvl019Ds3nPqyilSLrXIZNN8MVERmfij5n
ZxuHadtEhJSsSD0si2HaZoQTiqgJwlDGZs8bfayyZgCJ7/00Z5fySheRq42x0s98K4IHn0aXS6EP
lCKjyzJwTMCmqKkYj1tHcgtPYe1Q/KeVegHELbxdyiCJCeMsPnlDWo07huUJJPMN5MM+T5jM1OKZ
VJ4mFLeTUJVmxZtyH8LU3fuPSIlJcwVgY5jwCp9XqOOGLBqoavQ+jeb1Hj1U39FAWx9YEO+Xd/Mb
FuKRhG98vuBc3vTifZfJah/USt4YEZ5Mgc8Yiw4gvZ5gbCI8TfZUvj4a9zGfhZ5wSPr+S0bFhqay
aczkcp6Arpm+e70Nx1fHOEQPf9Xuv2DI8Jy1vi/zAiqMF6WobF6gMbR8Y0Xm7ARQrfu9Wp2juJUY
nnqtPNXv9qh5pXy2ANoEpFt1kjvXGgNGW4kXMne5xLwjhqIbcCYfQgP/St9Af6kgmsXS2sGUlQ5u
WP+ijXI9PfR3OSqrubybm25CVTx46a/30x5vhZp5/RV+eqic/57o+qg5+myGchJubAOlcxfPyKb6
XiBbkI4VJl6bTvM7E73RmunhATukZoim+JV8HE90U2Q+U4ruqV4WBCHHUrNaIucbTNWRt1dUUzFP
J/GNvw/rp+B+yj/6c9AW8K9DHi/7J0K9+6Ty+AcMovEup2Gkgzf6/wzTzpOn/BaO1YHev/xk6Uqx
La8f+UQKNAnfEZWtV+IgMSA+JMqYy/+n8rpT4bpjxozLRdRNIubTnj1a56xvnpTEz3SYL6lILAtQ
sm5daM8rwqsQ2cYRz3iZ9qnGKq6VTodBHMVh6m+r5vknQTaInYlNIOAmZ7ReDMmZPZLOPHqaSPpL
HKsJ4QnVvAXiYsix/oRUjJjfpXTo7nsAChQYE8A85FUPmXQGCzn3cp/YAK5FySVlO4zKnknf6X8z
FumJkW1l4/xv400jAqIfrf+Dx2vSyuRy2dzgubY6pU+vN6du4v/Bj8W1GcAucEv4iatcQ05n6NNk
kwluW8d9zgPnnuQ3WRw1eERBuOKm7MyC6UGsALU6dy0RZ3Wk7uHnGJfr0wur+lN9ELEudQ4OKvvg
JMAoHTIifK0mvwJKLrRiX9m9jCrpZxs/rE4F/TqfmabHB25nbKVlr1VDuzCqzUOmPtQ4NrrhewyB
8K14QXm/sQPwLQkIcBYTmcGNPl2k3WesQ8lLor9l4uuVT0FPW/HzUi0vSlAO+QAFXYoglPaQ6NOE
tbBzCHdoocHQXblE130bky0+cks+LOn9kDvh4HhXlmKR+858fGv/0mHWFe2kkiUXtD5eX7F1kzXA
YFzcztf9GrHp+juOHD6yM5D/vOtooeTPBX88VnYSY6dg2G/glL496ZgIz37L1vw6MJeHFj/J7wq7
lIDDuALV8Vq72T5s46di+bQJSeV7Msl9+2WxbppmkSBffKhSYHUAaV7saZJ0h9XXP7kcv8TYWSOl
X9PQGIM0+bxvnZrLxhmbJ/tUcsMIzJfak4oGKo4KSgfcw1I02fvS3xMy+V5MDmjcbpmru4He6Wcx
yc5aGJ63S9qEIMGc4GbH1DdKRB2Jh93t92XbYR/FfFPsuJQei6zOSPzOKqSwrPKtA7p5PYaVBF7H
j+gU8dl3Jj701bU5VXp1nngOChee8W4DT6P5bdsDBjGoJMqmSl1p5q3H0yTz85r6YEDzUF1LmCys
ECxB/SxNBow3DFHDCTw3GvJVpJeoDTM1YS4aoRlkTndgAarzpQHmlT+8N+M2NzWnmzQqZc4+1MtW
WFSCeAIJfGRaTUM7SFkd81D6VTZzquMz+I2DPYgYdif42+ZxNzvmZYFAJ7VHk6D0tJ1ohk2xjLsI
70Sm9e13d2nf2e0JrJ+o1/Q93vtwajDSTgsYWlM0Fz/c2M5nZhXvfaB8A7h6QfAVK0VBiJDZhOJR
Y9sBJIVhPPIe/zEA+RCQpY1dePxWv2kRhduby3oIqhNOvvaD4/0PyUvRK2JHMkjFzOJ/NZlsSdje
igkzRyXe4QVU1ceykHcAHuk7/mgcvHTqsvc1+N/hk/eArmxlU1tocjo+cTssKiy7EqDg11mcamZk
zbnY1G0smNyYOmBxiik+Gj5Jc09L7FN4Rwn5IgL8Bk8neDzCQY2H4T+LAbbts151gE+3k2IpsAku
DnElMRtDT9SZ3L/vpR5rOai2PZKxkS0rUtTJZrzso9HRdQ4gFv2pNyQP5OJDD16s7KzU1jfOObJx
moRkAq84iIFdmL4AuQG+yKdA697KKbYGrnA2fh4EofdWgL7AFyJxwuWP38Qlsg8uAxmsV0cW4K+w
2nvK83bH4x4iRLVlKS9pKl+rtDinohi7KRTFG+PSZ+icSpyk306/mSTDCoCXh7/sfBWRBugj+1CH
o0ZgVAuuHulqPQwwwD67pTsEy2xgVnAPE12NE0skLutfbRplcKeFPnPkzBHhfN7yhXAWmNY/pMHd
kfpAfhWTD63WmzHQcFMATMxKFudRdBI3wpLx+IPg6oQQpiKnEUvdYhA+9LwIqllagRf/YUyEPF/t
KoM/Un75GVtBAcAAoq1UxdtxXtoN4c56NyOMjtboSnqYYEE/Vqrnn0I+ZPEaVLLN1UYpCW/I9DcD
U/eSpoE/RXgadCYyWrRRjBRRRc+c1lHXWRoV8WM3OK5pt2WHkvtEe7rlLX0i2uMFr2fsEPMQ+mo0
NKOJ5IBHnUap4JbQFo1rxfDN0PUPWheXRHy3h5ZsP1o73Z1+sqYGOOBQkGMcDM95BPEps8p6b8iX
ckQvGm7UjXFYgL7YGaMEKVmareIayO0ZzJMTzAVZ/8TKMWEn04ZE/Fwv0w8bSyjfU7SWlwN7Y/UD
DBXUQwfFAUPb63ovZF37q+/Z0jaNsF+KbA0fZkG/gaNcU4aMRwEe9s06235RnTn8YIBKLC9el3t+
hPiec5rIQpBr/ql7lAEaEKpsazR+HUb9gCV8CSA7EW0PwQgkhqat8yn5b7Z8rPQvG+9kAWAQQonQ
nTg8q2WIEWDFg5Ax+4fTOJDBD+Oc4Rd37iv/mAoGfMIfGcfCpXOXMiwXtUheTjsvBUdVVQ2kGpSt
t8yMM2DNnmGuKmh+dJ0JlZZum1ymiicfWVRqNE9QHPiuodJAwXakFG+FeH/p8A1ZLla71VO5MER4
Jq/lTcDXUQy+NbHc/DUnnkOjRkWvpL62fr4uqye/xu+jdRfodrTqPSvyWAjE0doa6ormxWMoJTPx
Rxz+ErKtwyyE9HIfEWPH1vP6GL3vqhlomP/kNLXWUS0o04FdhfbZWH1ozRF1YPNsdwd2owGSmr2J
Zog+0cdAHsoishLA926utwqNBRdcQZnSWmXJWLX2pcSh0q4rOgOI0jpONXRL9cxz0qVQAopSDteL
GX0eqWjWH0f0S5Mi7vV9IBLcWKUngEzuCNeCdu6aJKhfpw55FlcTSr1r7xlG1bhESDe4Eagvk4Dx
KNqqMmrSyDVJTQHlwPpxO2+O9hNgXmyXb5V/7nLPPI6Ls3J4zKhX74K8TxKbOnrWs04D6GcrtRQU
/uftm7cOCmZ+S9qQr/8Jz3YtNiqZSM6hLGQ0At2umcRcNex5KwT4Lcyj8kdLrPexqlnKZZOjVa54
JjbZTJtjIDau2LXAflr33yjM1M3/xp1XlTGJPt+3/QUm5ioisOmH1HTUUyolGbigwTu9+5IqfTW5
Kji92To8tDRIPFN0J06iHDkVFMmI2RXV041dLRDesT2kl7zXi6jPdZglV5FI2TAgB5v3PY4IqQft
cB/rnObzjDiO81yc6RUcMJIBqUeXURAI4id5NVT1r6v1HEpj+/FD8iSZZo2uLK3T5x6JX/BiA1xG
gltxvBRRcygQwfyZNeS+mXOhpEM5dw7p1jxo9KT4SFu5Wp5DiFhyK7A5Paatlxd5m19CE2/W31pq
H1L70O/mJa2knYLIvJTdB7QJ6FtwrTkjMClTD3xOg5nTBvsNKtfbg2xXf8Q3VB0InTldAXLug1Dg
b5mKuluq877W3nNfKguM9gWbeFxjrOgPyQvIM1TtIa48jPrl9aYPeACcEKYeBHQ8PNzf/ikHSPY4
djSH9d85d58Or8ORQbgCoAMBgwlPsf1HA9MSNkuYoLJrR1Q8Zdz25T+TEkkpSr1QoAQsxvqFKY8a
IsmjjsPqWF+6zcPcFFQq4t1Q128Katg/m6nuiTA5fF4tLyc1O8bTOBbo3SI3bq4ehj3E9vmJWQEU
553/de+W0ERxwan2l9gO0Pw6YS/hKkeSCeEX5PNRNB8JI/tr8W9SpVxm+BlEUPWkSlcb7Nwci7+I
AwuUEYnc7pwjh4BJ7nc8lAVTCCG/y2w5qBzeTddtnnO3SWH41Cv/DRppeDTPyf3v1D38B3NPuxN5
PRrXlkKehyi5wTw6Svi4iIkYsJq3MDLMSXrGXchqwbYZwvQoZtUwgk70bLLcP5ZRieHpJjj5m/id
mhed75ri5Tnp7g0w7dlUVCYlE2tH1RahGTJtLmvn5gwC3t+11DvxqXbvsePqSq9gbMa+5kQ0QW5A
YEDs58/56U6Xv3gQofhMyPp2CblITWm/bmeBgd70aq4rA5Qg1XNqpo+hnDQjrY7I8hmUSI6h3eB9
kFv6sx/m9xMz70RBV+lBNxDj7/lpv/jdG8MhQPs2hn56SbT9kqj1rk0ExXAvmQuX0OZhFbDQJb/+
3U2xjiKWJnbw/lua6UCNkIzI85rBNnZOHOWZGC/4hmm7VZJ/d0gmwf+J63svXeRrz5/m5PFU0yVk
+8+/CoyKNceQ/v1TnAXmRreeTmofQAKJcxP9TZGmAYVEnxydLboKXpcrTR1nB+Peeoq6C7BB+e2F
vUVJqq2RZJ0mYhZyRkdur9/eWnk1wOoVoq8FeY3YrAuWDWpp4dr6rn/V+bczj0NPHCnj4pjlHODn
6pvwHEtxvXZD/JGhUR/6VFte9JO/6sr9Ey2Xwfi/noFeamqzrOAwgoKar9SEBaqmSAI7HlnrD7U9
l1Yn60dUBTksrDbxdFe/xt5n7afxw7/dKLM5zIdx70gcXb+FZ8CWGKaUP7tf4yJ0WxYBEI0LzsOM
DRKnIagzJurU5vTA65n/coav4X1GrwKMH/qr6aJZHvZOU6JdtpHGSJ59f0r2snavm8XnS0QXYcK0
mKEYJm5Ex+O4mGHvLDH3mpb+zZnNpnF3PmMkIy4nWYcBCAi1UwkxYVSZfHQeq2NXJDv7/cGRWKC2
tmUkIfvploDry3QCoxgwN++T0CqS8pUNx0JnRxHygcmB02vDLsyFHw/ghgzCULZrM0jZQIemjgF0
AtHExx0IvGADPPzd/f5GdHPHYO+oPYZ0yLq73LVZbHeIfu5l4El4nIBWU9Hx3iOYmD5aXekJfTco
2wFXcUIh1L1RGjwhPPuA8qJue/d/yuw+k6L3YkXFDRnrRO+XUiqKdLnYrBsfYe4YGwT+0fWOcKOM
hwYtXcQsBOK7tt+C4MQuYsYjC6lX3SXlYtCPLlGJLFMJ/PyM3b7S6PBzL3CrUdVg4u6nzCw0dz6r
6PKKdFQ3dIjnfmUSToqSEqmISFNxJArxu9q/WnJE/F4aKmzYkOBoCFmZMyuU96x15FB+bAImKKKI
Ks83UhC/Hn5RtRIAzKmjhch0P4zz8cBK8SGoyePHYzydSZEYVwonAYeZ2FjxNyNOzT2+Swk2BATz
UrCdw3PtjhqBvefN7n9LghnP5grzw3TgcF2k/7440sC1t4cTfi0NUr9rWrG/QaEasyCV5Nq5c8ZE
knNc+hZOvvhqWb8UMUKyx7/2RzldZnxHrzZQ6MJ670aDebV2ajEldgyj//jMXCTdmtXDHaSMCjmK
fJktjtKj31I6Yv8tfiNtf4JpWrblqd3f5Oa/cu2h9D/2gyo/Ioewe/eFahZ7iSpCZz5p0RcoB/Fm
Zd3sIzcOWAMKusoJjD7/Yn00ZwvTENOttfS0IwtMZEDvK5hd49uJQVynNx2T+yQ4Xv0SdGCLHJQD
Cnl+ZIneKPafIoG7L2DwDCoHVOgE9dfiBiCgI9xby5cy2zQ+sVRvS8zL7WdgIxXpGYwPDHqDZ9d5
GKtIveS9RpofzUIRiNNLLmSnqDwdqkyxq9SjCz/52BgMWqnCpm0tsFQlMOPmKKZ1jge50DZrp0Zp
tmOdg7nvDQxb9Y6CP0C+hnYV0N6A7XUM6BHibCP2+AqxWRVZ/tn5UojD90bcL54z+wCqmje8Y8AK
uSjOoSW5HZ5zMu+82owMBDQOd1hEMFNHqrenWlpvyVWgbu0QuunzlgUf2HIEVVXGPJh9FFOhrEk5
tvlHtca1p9o/dGB1/FfjmY5aKi7RVZZkGY5dorYUGIfhAhtGRA6cwhKc3yzTEcpOxSGULOwfAgb3
sp9cUuxczYOZ74YGNPR65IfHBcYlwZmNsmlN8XixTjIMl/CGKmaZbf29+xaKAQi8d3ofdu90L9cv
OFPtrQQIKcpnLLB8G9PYze+jEKTqLFzxbqRvVE33lhXb+YXB//cZ2oN5o/nANs5WBMxbPgTmg5/Z
65CMBV2JUJ6udoqcKd/wlPOWBhpZnc4D/9NlYeL8pfV80Y997xyNqshNfIZFbQwhel8OdKcfBfXC
vH2BIF1ByaVWfJoTemYowuiLDRp2kY5AKsNNYgxN0er0RtGLJhyYWNoaDk3Hx0oamNzmy7GnyL8U
XjRikn4tfyQIh4F9jlUEv705H3cN6PVQM8TEwPdVm2i9dKjLAC0sZ4oo0kto/lUrCtJdx6quvkMy
147GW2adRMit5kLYxLGOZrfhMAqGXweDDRDKTVlUDx/frz7DgA+pX5nWIU5hqTgltKKHAfpv7bSk
AX9BXbXq+cpkOYqYKqpyHhed6RAniM10v8zAAYhAkkdF1L7VLk6tOS8dk9No7+fZDeeRpNfFZ4x0
HB4bAwE31WSGI/S7Cvdov65+V30l7X1SniD8fRWHXwuolh/XCYqR/+u8OYNVuIrnZVIV+7WFxhwA
6hwBi53BFSyeLIq+F5fxz/SCwPpPDjWrQ2kT3pkWy6nD3ls1PeM/2OVttM/cwg7kPZcc+VdTaPsr
1TMD3d7xpZETAWNqz16vjhZPJ2fgNKtAQgsEMKI4DKc2cGUHkJ7hbTze9yFGptq6aRcAKjWSjgMX
koUvmX/a4fyNbuEu7cBJt8ObQ4vICGWuDNOOjQQVeiH0wZ3YOcXIgG+WGUjSSNyFWNW63gtyvjv5
BSTpwrdx0bkUfFpGe0Wkvmk4EGrwZPDQe0+HRjIs/2hwgjMZ+2wuk/0QOGnEgoINTje5zxSFrVfO
zQS9M+bs+nDxSXdtTxZ14Y79PF2VyCT//SLjKF/BrtW7cPxL4lWNGxgWP40tdFkIgqBXa4UbbDtA
+aGyC/AMA0MDexSSqN1TTUGW/4aU/CtQjj2MXQoSgy9QHpadnNoI+OLq0Mgq/HIQLvw8coAOcfUJ
FiXGmckD7V0PjzouXtkqhu2xTWF72xVvF+5BsmiIF8tevVTvnBn27N20Cw/Mliwca6xssfM79P1s
wceGnDmZFY0t3xYdDhIYb0dVartaHegjSvkaI/KsDvzbufTLBnh1zkbu9lXtSc5jj/X8zGULth5i
4IKBCSPyQeXuvQ/O+cqQA/F/SEG9Y4TDrqMfaMhNRYl3fN8xaENU+DdW6ff/yz0PAEweaCtLTIcP
qiOUFq+PXMB8MDYOktNP6VRlOoRkTTJ9DfUeCx+p7kSDryYBnFQneQa8PACTrCd5UMYuxTlttrf/
hkxY1DRspC5TL8DoTIampTKSaCrxAMnNFHYydcxohxt6WBFJ2XpQsyaRp2nX9zFbw7L2688FnRRa
aWI8zgtT5lJM1EAiPvQgLp/We4lcFEvRQiguR0bIJdReqYWnmmDNyPPTrLNyeRnx4bmExBjd2e5s
wSbGRiESnuiTmLcSnJVochQM3ST9rPundPql0B8b3ktTpBOQoMfkl9RMScHUzbg6zA0kQmFXlKvY
3ZZGNZSHF3whZv2N7zIGu0cfDWmRVE2sD5WcEE67e0O/5bJf8vDdaUnbN2gZ6n8bmi1UtzqqIA9x
BQJuYy2Z7ormN3Id/aMUGhMcqs3oBtIHvW8rSApdRd+9IwCgZbkmJFZTZ85xUzuRdViv50WOzbVL
U0z2Q/PBHrehs62fIXLMhAGTWkilIb51AcIDfK1rCUza49dIAwqhUNLcoxVBlIAHvE3NPzlzd0G4
/7lzvrgTkffplDQSMLbFV+RQxYHkdgGXqGrhZJtthmLB60EcfzwZH3dZsZ2zKnQd8dJjfE9y4C0x
sOcBvZ9LbgzrsyOsFcevCaaXqPVlCCyGsxugtkTbY59k+jNLY0cKrmoDom6wyqOrzHZq/K90Xx/C
TCWL2ZgEi0D/wv8VFjHE1C4Z31hCuH3mKVQdTc3ndgWpM9QV2L6CQW/bD5hdWzKAMKL/rd/oL+Cz
L4DGIMrcGSfGDxU66N52pk7VJ7+rEoL56onRw9FC7+Rm6Fb+iw/FenSSmlGsliTxRjTT/H0YEuXM
q0I2HE7xdwyd6qe7GtJM1bxr2RTbJFbRHZPDpP+HchNPcMVkn6AxlOzLwBHyNa3ujERJwpoby1oZ
SXn6BYTcsB74UFhiDGYg3D68CmWTC5IePltKsxpkFaW7NfxQNUIUSBFgcEGpKQHTz0l6pDqHKREf
uI77AUHi0zmo9IHC/ga6IqmxWWUwYOsugvNgHYcODEbpG4nqo1g7Fwk5Eg2CKuwYiqJv9gcNTyDf
zjNUzHDD5TRtkQDm6phkdeZWK1sof+9NdKSk0DemimqY0nnOVC0jhb+hTSqt5qhlUydHqQr1xSdH
YIYdPOK4peoENrzOf7I47Gh+IVX9BXHxITD6MSTGvdaM65g0MyJg859s55naj3tlzQGIlMyb0agP
EajeD0ad+Cpd3Fs2MWTcX65hyEyZ80+9zwfuazur9VURd0hvyURTEOAzMdaeyWCswqZ2QIZZU9di
iaLmC3cpjFXdIj2f4aTjScTSRXz0rM2tvhrUlyML0m5t31xy7cdzPzzYNVvIYMAtwFM8+1YCdwpc
iAquQlnVTVzVz5I1sAvQeqgWI2exMlA19d184ycPRHRnYtrMe8J4U1zEm1DgvZeo11whFmmfcsS5
TVbZiGdbPq4ZwFkbv2VXoQoRRygPKQHLl0ERVXV6TvcfvMpZueVHcanSfIsbz4e14BTTbxtgqYZ9
enIwyri3jZC8AqpUrpKi0nEVpZrkfyBFzrLg+iTazUQBrDEUo4TL9fQecfgmbtVllwqPLxgpKmu2
lif4KKXcuTxGRAnSKcWxqcUrQSnDRnb28l4t9oqGdLKfgSECQEsoos0OrBIGm/T8dD/adOBj+jHC
WtugaTYJbtXz4muhnNNKQdmuPqCKEmqRJlPqYCLwl5e5PJzw3G78UxjZWPmZlsfSTKpq1Q8cCzUZ
3WLAsZAqs9vP0SsRxmxEZ9l7Lb5OBGRPoDRU5EiYIcyYZvOv0qWmOO19xXDRwOu9PcDXYxnIgkXr
42LOmZcwllUaEK9G8q7tuIkDXBoKgseAXD0WDbfTXt1wC/2KjDBxgipowZpBWyuwnsF8Q4tgl0QO
rG1beyNzequBHPsSN61MoOWhyQVkfWEQPmuL2+Gdv/LbpwkM6tLihrlFurMUiCeEHNhJcKvcw+BS
KtbXLJqITD9G00kvh37KiexrFkhXQPUyu2do6GJLawluiaRy/H9R1+NkL7YEzBpuL71tnDTD9LOz
nIKqxxu3iEbJ2bn4mz0uJj9JtQVb7jLMOlpgeOaJPjynJ07EhwZ5V6aLQKtj3+Q8HXZOjLdYr8tq
A1coBxXpUrfp2BwAQq1LXKTCz3EjYm/+iCj/f3fWCpgy6I/eDTKkmzql0uWLMUPlY6o71e9aYKK7
HPmxL+oqvswoOu5C9k5ghRQkHEVTSeAyiuq+dSKVZy+iU2MWczcrEYElLyi75xv/tZxYHELMMmH+
18cx+8lOKpER5WDeDrWURAmrcOsKKo/KT6GhBrc2QyU9ZjEFUWy6DFkWaOHLLt71iw7D4boz8LO8
3OJnMOa4/3dAPXvp5WnDbysraHqHMJXbqQoU4aFurTXHhpiyzezb9K3cJZNmPdrvqe5E5CTo6+cO
oIMz/2TDYVE1oNSwm6UuqA10H5rAETc8nAkSg7vSIk4zjy0y2f/ys4OTKirNxN28ZjsxccI6FyVj
/z812GdKznlThuEMPoUwxPT2a+drA6X8kz8whtvyTHSsllF5oVWpfo3K0ie0VVfLHDMGmJArt1dh
xsmNOdk11gE//BcYQiW7cZ6qaX0IOPLU+W70X5vcp0T86Hp0F6nRoUxtusRO2yXF6MgLbbNst49S
d62gkLEMLVbc6zBpkv80LWOGNMwkLNlpXZ8UOwLQCSicQW0hOqqZ2cFcdKcUs2gTlbdtm96kkhL+
fki9jWJ2gPiSoILrNaoxBXBDYE2SKMohVUWFT5tGVTA6JQKPAJ7bh0oL1ozP9czCIPT9Amj0xfMn
CX9zHqa5NoQW3kwgPUKzIkEbGavUhh/JfXhUYJDEhHwORWLXCL6iC6/wQeiCr9A0dcLx8UWOGOXm
ds/XGEdDwtrRaBtDfdr0fDlWNooPDIywwWPAnXeWii2BJwKqY5gQxC9QfiRZDaQTBxN2ek2D2/1+
GoHAZhBOkDM/vcz4TQSDD8AnD8kTeUximoGjpxEMz8NPZGUQj2lF8FhjL16uqH4+Qj5UriLTPoR8
EGT/IKsdEW30npagZ6tIk4HtPv+4TD0MW7Uz3lvmskNTna2TL923K11iI0YDsE+anpfLRJQ1QUxS
57vfbCjwpOP7GXoRCtBntv+kkOBr9AEdg9d3EWOfsNYYswUpPOchLpsC4MFBUT79bjYIT7h97fUz
Ov5QYBrX2IU9NYTk+QMV5yC+3UNpKji4kGDYxqHIqHnAZ+03gapcBHEmz0gfUI8PYWGhJvt3rZwy
MypM+RBcAkrgfgs2tFkOsY8GUNTUo48c8mnfPAhkygFOVwV3o3EqCWSMGGRFIzUErbtkuVLTIQGL
Ru7seifMVea53L5f0GjbE5h5FMiGs/n2+NLQ1/9AKldyQVRbTu7AQ9TXqWdEMiLkr+TE6oBuVkkF
SwYLgzDQrJZwq+xTk6Jy1Yce5aydA9ofvpMXUB70QyuqzqItZkQq5uR5H82d8vAhzXTAazZwKhZN
12H+ZJBULRvm1KGvblUuNMoKLBifvmv7hNGijTxX6r6Eyc0QHLbPGSSYW4XMFYzZask9yy+bK8CM
/74HTcwwi1Z+PBIJB725vxg1b1OcbT9SB5fj6YbN5XMkvw6NiUQKHu6BBcUmU2TfPfClMlftpU4C
HjGBTOaMfzD+ijovTe6C78jwKaMweZZ6C0mLhV3ohmQ1w9VzBdhzFjR31GjOp4daPue9ugc0gqjq
BXWN7l0npsQs7YlFnO4KvLizNjD1HIusqvHeCg4le/EAk9sRaupxBPz/VZ19JXpM38Vk2kWWt3b3
huzmZhA7Xests3Ae5b28EquFspEMYZg8bJb0WdqLed5I8Qs3PxRfd+7f0mwH37kMXsZPQnJbXcA2
zjWMnVehCVbp70Hffatc8a4bKkaZsfa1opVypTnwiLd/dBEQ8dPKyp091rhKwOo6yr59KGvQ/9ns
nOB5n08iPMELlfvSzAtUq9UlJqmQLEU08wYiFmCXQoSr+7ITRUNlt3rzgUGZbtvZ8RKgIZb8Ciur
21tvuSzukxjqLCK6rY5YbXhMmcieT9s6s8qbzUWpILF3HmlLSd1XoGB94EWLDvmnR60kPzLZYT5f
60KdPClMMr7lQ+oKzKYhIVFi3mn4Qj5Lz5BdRp92L8piumEBNxAXGiKCv6eZ9Wrm34LBpAH/RQ/T
YztqvSIlRDi+9la5CcpND0kL3POziA5LC1Q/LnwR6UhaBsK5ncjC7gnhSNd0IujDYRxQNgcEDU0g
tuF+CqWGzg9CxzMYt4sOTFRxku+ZdUqns9EdgVlUaFVMTF+PwXl3BRp4FDDK+itQFEbOfCioM5Yq
5/zfbdRuvlPusUrvIvy21gAB3Q5XmaZ5Y4+h74tOMxqx1bK9sOlSl0kmPXFZviib7VR4MxvIzMNx
n1Z8/7QnbQf/8W0251KnPsk1DA0IKOt2wlOT16qGrPlPdk/B/2VJLi1j4sPlUJPNgVnIz8I4tO6b
TU8kjkPPe1P5hSDUWjm9uha8xZrcjDXcB3/+Xu42FO7BJ4vFSubQB0SDyEwPPB64kwB/gp9e5owd
ihY6oKxHfzTyfyD7Fy21/W4am6620Be/6/aocMOpZGjp9oG7Dy8utsfymxQB5NAE7uxelzNloDko
I/cZ5ATryAlyTgpk3b8VSMH1aElXgYzjZUpISLNhVnqY2rlIKOTqh3WQAos5yTHPR5+3OQPYTvY5
5FvqAh+u9R9CFxtNA/JyJ7dTA4lPBhPn3cPg0Xnsn4ey1qgRoJO5LLkHi0dsv6Ggxb8iBfrH0wUY
ptaVeEW8oEBH+5ionjUlQFwTJoxoefuL1j26RrXKiTn7VVDGCjbwd5VnuG+dL6h2IK0inpnAyKzC
klGikUNUp2qQSibju5vyaC2CJ943twVMSKi9qHzsw7Zze3vC4AcKjj5K2N1x8tBlqCeOtHpdHY8B
r2MklmeQlHkZe9tjA+v+GUSdWhmHdRteVFSFu+ffSODM1L0fzTS2P0s3n2WeRfnXzxBZ+jQxjXzt
1k92ctbXBcX0M4CucXTj4ovfPwnn3h4KN/Hbt7j2SkTWv1dS1WamLP44TL9NWCae6Krt7ZLyohEG
tuF7+aL84IKdkCrwy6jZMxQd13W3tD9ap6fUe9RtEYZ9NaBsG8/f58i9IoRuCq24X+OtDVR4lTAT
w8o6n7HYqTifjfDLqZ3xuXiDJSAndctbVTnD+byYdshmAOiKgU/aRB/cW0QDbpXgE+qFTqYQ/2U5
+i0wfj1apacaabsSZ8MjUycpczyvwFwJhRtk7gkDIPaUDPS8PNn4/dIAHf7l9flM3GYAr6BR7GE9
2wCiOfIAUhL0eNH7qoDd1Vv3zUQ+lOGyN3St1Q0pk0sBhmUho7xQo2S+Do+3xKeTDIEM+TTkTdMB
lCjn7ZQGktqtjMgXOkIj5JXvsUfcpu0MyBjDLoAVi9s7ZJ3pkL1htjn/UL/TFHhhkjHt+yvd7qXk
GC1W2PPnaXJ1PwCK65XJblcVQQFipL5JMpXCJMdW9OLDFwPgSyHPYfx8T5TTWWnMdo+ykfW0W7yV
d99rEKLyytOxvPXNlStgRiKVIZmLvRq1Pxc9+xlEbPqTuLzi9aK9j8AhZsphqX/KuBajV0nLPfXb
XF1s7zIvyhZ0ia0o4tbgQO/SGUEhMU6hm/rOH7+z7ouc+PLCynFp3ctwlzHf9G9yqjn9aONEOQ0Q
FLcSYVdw5/I8PkHPVmpt6G07vNoZYYBX2PpBt3lrb9q3WKUHkEUOLjixgXyvp0ppyPuuT3H1FyS0
kt56hdZ3m97kSPX+rfoAY+dszAYY/3LBLJUvsMJGBQLd/p0oEl67XjSZ6QoGeNAbsfkVKPNccnz+
rpydk2DptO47WO53dNglZeyQfu28C7FWoqywd7OTEu/8nnrRX8nvQQg6xw2BCwW35iiXxTyvuhb4
Coki1+8Z4/qwnoupiHXvn83eg4BLTD0TmbIiXKkDPjN/kOtudrU8HAhZ7AHKC13xop++ZuGi8AwX
tBVF9ETK1spSSIGywfLFbWve/9VtUvNYTpuzGwLDWeK7o17+jMkW2eJwjUzmwBbO9Vaotmv5BjvJ
8k3zV8qNjSV5VmjWH+15hajV5UjqtGuvgV+Ox5lxNPFRipN+GKwuUTNEKVydh0oeDSlbGNpWh0WY
2oPTCjgSqUiTxTaKqZ4zCqLr6LXWaQpXYxAFA3hr3yPXSRilZrhk04UH0kfe9Kb84UM9SFQZ7QXs
lK8iunsmiT2+cejNLN++AvXezoj7FbQ042g2r3J1k5W4B9LlwIpUhEV+Y+wqbFZKYbUjt41dO/vY
whcF7Tkf4n1EoS/cuNXw/aDCNu8Xizinv14JcYUtxP0cgbwL3MocWkyv2ZSsOmHVbU6pf/FGltRj
d3DcMRXZ/Hs1HKp2UhDVsAxyWbSQBMhvzkOLNjrVwy5LRfdxcKNNYh5VTOM0EsNwEuNxJxy3AJgr
PhEAHeq35TOOxjwNiMZXiJK24tbfY2laNr7ibIikv1nS1uvxB/1ivH/dKxVTIzAux3Qq2KnGl6pZ
3i4y1o+CPECJKDpL3N3ZZ8WO+Bx15FVKpWmpPPmMdUl1dCPJR6n+1ypCwkBotIDHx2tUnD+lKvSs
lSPFStWYkWXm8EbzNbGPwYe7QjDwgyxo5+CNgrYJ3COZS7pP2y4lQb9PP0HKDZu2R3tdmrlnGKi9
DEaG1TO1QicrnldVqyBo3EcBSmng7DVgalmGpffGub5/z8n9ZMuNfY4YWNuvZ71C+hXOw26HYk47
MQaBbLn6z5bbMkSJmBurCcWCxZAYJvSUumjWqJ+kXdk5rTQaOosaNgv69M2DsAkEfcIEagMYscMi
60zv+d4ECbRr1eAe9s6p3dw19XshZ04jr85wlMqIlBuOldcO5lMTcLCnO+yfhAnz6RtOPeDw4Pcq
AZN2TIyxeGYdJIbzh9uJ1FPajBSERTDfrYLRDiPJm7vlxJqN05PzZ5YkBQphc3FV5soJSkmStSds
0hIApfeToNAu9KcXazhTFDkHUn9Z4KFImEjP8PJEaOjQO2KoWzHiRP0XlYzh7gMAVEEw9Ir4C+Nb
arghc8P98sYD7i7PLxG6CTgf1M8AAZwEISvkObeSpvvjuGUgadUm1OstVI/5ySYb8MObWoBrGhME
fC50LSeJ39jt2D5AheoTDZgB+2i7BNzod9zahiwcYYeo3CWEvdGIT+YlncxanJcIOrHT2ezE1JPz
dZ3De/EATDz00ohmI7M64GCVVy7dT8Qu5gGSRTQsHDEm3HdW6eFlsi6D1LRztVmi68mT//7zPfAA
bCGfqmlijMnQ1gsODhUPlDTkDemBtBi4f6BARMjSxCzzH+0tQmTw11i6y+/ZnQRLhubWyKL/L39S
BJfT2nwa9JriemEHeZhLKnIyVfrA0a/tB9ezVSbjeUvukZO0pGVnNvsEhOvMMwN0/dXljKFdjYWM
RwsWSWB/2V5yiT/Jzca+nncUWP3Kt2/zd6WTTW8UMe7P9+h8VszhVpMMcWHdnY3SKFisLC8hSpet
BPjSMDiQRZ74Z8TEYA31R/9ZM6ih6JtASXl7m48lQs+hQzVvDk36tlQH4fv1r/Fsv9rVlcjCkAP/
yMi2b8rA+BXyGoNUx4r3ia6tA1B2BofOCQGgvQkXlUOxEcwyJmlEQlBPkARWx36vy/1xM7eOKAa9
CLCx4urSXS53ReOOy7fYJ61zNx1EaLf2Q2Zft6cmp1SrWPBFvsl/ppjNwyzwptYuROUAgZQ32uyz
+w1xPNPc5kaPWpSLYuXXceE2RQE+ovoSNzDVnkIA4oZ4hssQg4Ge4PQcZ6O+299Jj9H5MCyCcoQO
0oUfAZR/oS5PSmrFP+dBTb7LrtM6y+02zVnTJQCVAVeW2bZ86CEavUzvIOPFbkig2nx14ScWNEbg
ZgCpfJdrFaSTm2XCEs10lGEikuK+R7rb1Gm4As/TmpnaYKcXVIQvhAMGmUMs9HKZmPA4uU35QdAL
LsLXigcT8FYAsEEteffWXmc1WgRlcUMCAd7OkKkau8Os0jAmKyTUfW08er8FFvJ0FGa2MLQ2FuMp
qfZIrtATGXBEkUmSbU64kSDRMiVV8XiTB2qwZ5JZSQJV18FsBYAeESbPn08F1mwJNENzVboV/+Xh
5Pcv+aoSBlOSMayZPuXk8LpDzRctnyO4pzF9bBG24YjGF9QJfv0t8E23hYjBMDJ0WruFr2EYcWls
hErXUZm+YJmeebaXGz3huyUSjBMXNsA48ReBEQgEOR648wVTWY/wKKh2DEdS5ezqbvnOlsFYk17q
lKQr6IAnsx9gwdadwDL2zq1f8M674azJ7R+/e1h6rNQhGz4mzQ2/lVHYqH/TgM+R0lgDcKLSIWHX
sleFNGyllFfOwBxJ7vdNTBrHn4zwrnAZRLFMiQrQdy0e0XgSuoaAD5adrOH0LvOsn8PyZFLWhOYT
gIBqxBFNFViZVX1yWvvaZwHxu/UYxJQzwDgGh0UefJ21+ODUCXcrIAkUa5zJWGrnKIVPZ9DOBBO6
Iu0NDTE3hGrzGjvCIxCJeIGHaus6ROFZW4Qb+MSlM3+gDbNPGzSitTHD8NldQGyhXZzJt/j2x6bX
8/GEKsyStfXVf1+NVT4X/5eeJwTU+4yOGmk6VLwcvDvdrImL+nqp11jVLubizP8C3Ls3nKn7hDh0
o+i0XrF0zQiHiR2SBZ4bCXu6kYfiiCfcf07I3GbSQrN6ach7iIoAdpUUh0GDZxAxsTnmIo+rHQgP
CJsHBVkEi2XkVutCXdgVhNr1sW0/QWIAV7MJ5NcXwCp7BbXZwSCLNIaJd5ObMSpxVA+WUn8BuBem
wmvCuBomqbyeCma/uChITuFxnH/no38/+whX786Fj42THZ5m+Pcv7myqUJk4hoQS779EEBT7gexh
0ayI0XVrxBAf1ack6G5Kpxnvo/qkJWvph5+wiagxCcEbsHRxe1pEoRAO2Cd+avgOAaOTSy45Z9hV
QhMC1LSjwJljkLra6huj0AIfrdoEDHJXGf59JQdKlfIIj4NYx9JsYq4HnUZ1+Ctba2MR07M3dAVn
KlVWLobtY9opaOHcMeU7tifYSAyjXl5rqLFK/iaFE+seLFWiZimGVIUX/W1KK/rIfMULIp4WNVjo
F3ZUQLkkp1vwJ9QPWj+lI/HMQkYugR+GOWK4zvxoovFM9H6Tjc3ZVMe2NQNJW5bmiELDhRP09mwi
EzR5jW9KAsJXqdt3EGwMYXFjtgH+dVT3icEx9dy+a/SWkniwpG8O1rFowt7fA+LkacCNB7PH/zaZ
DgRw9oiD2NikCswB6AlJoVFjr/EPQpKWiW6fM0h1GYvTsxWZDPBzxTPbAT6nOBB6Qzt7b/uIusuA
cDcKzsN9Kuww0TZXpmVXp4bYGN95Py6ZkRL7k55pG41ZVEJgNEx1abILz3HiDTIWpp8A6l2dfJU5
ynyqVu073+RS/K7txPZ2ZACnsoVoKjZfgIkCEylKvwA8oBDlcVH7LR8al9NCmSPjxFQ8pJLtcntp
t1ueFY1zWNiKKTbXqM2ehImOedYLZgYhsA84mUtm/riHk4AwMl0eowzMVP+DvGCPAFq8pKrSDife
iFGZfk1fYPC//cqw+tNK8IWPmYVZ5VaQ2xN8AbkJBpvJAkVf4qC9YnUUwJWSaqSrq+mPagqxdRYY
UFeFeftIxh9Od9JWTH12N5MFampqM4nNcBrkDY9jhGpTD8XCuJoK2bpIfxfHZ7avlm5ZpKtXqY3O
/uYuZtpRdDJoilh3MFn3I6p9UtUPmAraEhRV0REAcQEeIeInNEJV7QJjAMafP8veOQKasELITvkV
iUspl5yvEKVu3tFVmKJIKrDjyKf2scNgNAT+eDLJEzDsSnEunPFQ/M+NpPAGjPrc5q4hqhHXgRPN
mVDVMT6j2BxyAiycNsFzJyRmpnkuYQx4KDVD0RgVy3p2vGYMUYFX+S0D/AJmMO/1yAAtEgBI9SVB
InnMbVnWrQRLslLBSdqVQaIvcM9Y2IwoIe9v/xk+gMqSlQxeu7WgYt/csEp1ntF4xwAjRH4sfxi3
12gOacbDuCCI3jx/DUJyeSD25ctY8NlVWZfCavsCT+8cSETGPlM4xuAPuPw64V2th0uUAlUvXwfZ
YMvAXk/ThB17bVTRpcVzlex3puKxjXCg5uoHa80IDGvT8glxzV/ZMdJFJDU4IcKN1gQLqJczvumq
oFcTLXBcHXUIOS0l2oNbLoJ+n1+BGQmtx/bBw3xtmJ6gEY5r1BoOcNWEIW2tK1wIBLNSjSwDyXrQ
mb8SiB+T+d7pUD9foTCo8PbzSH3fOUhIQ41GKbXvqURXbfqTfdAaWNRXqnRP81YASumaKhivcTvi
4r3wmZ9DS/LPsSMONp+iFZaJYw9wobBao6QQtuzTqMBV2lFNGxsWi8g1wjv5fxQeULnyQxnsLd+0
C5k5mkitDvuulgM1DFk0hMK5SgqGiktRpaRJo4WhF3JPBb321NgNZMrzZ4vctfkeG2vcGMqoNefd
Ko2nf4x7LdoGprnBuaxf2N50C6eIg5inVTCSysHlpH9wkvhF0GcWsYccF8t/yYpGANVhUX5UbO/g
zi1A+WtV95/ZYLbYcs/c7r4I2SGTgqvfpe7HdZX2LJZ/CvYSeqjT6/6Hq5vZDkutqraIC4UNKUjw
hgnCuGNrFRMvEhYnkjRsV51UEEOZIkvaD4P5dNu+NVciEsLXEmFwQvGUvrwX7Bcybte30mKMUBhF
f0l19kH+/DoyDw6dJNU0BqIfPoN9AOSJOvWuRPjd0WehIxZjHWn/6J9Q2Wkhur3w+XPgX+kO2W8Q
NIeNUWWiY7uvPu8OsUq7osd1LXVycPwTNybxvdsevk5EycCnPl6iMztF7TY0XtO7MJM/GPYU/kIu
nyD60YJ7Zc0vIQA7DY9WWuU9hOTuvKYYsmBDZSM2O/qfIlkWQ7fipouf1Y4TCJk/Jg/kWF72Aeli
fbi9E+zM7pd0f8yb6HXsbHL/Or1dc5hkOP/n/c/q7Aq+KtGIwKP7eSNixNzW8iP+fb2P6oLbxeuX
jV1igm+LXToEz3pJUdYhVREYHQKvTY0oiA2ko5PkTcSebPmTT/TVtUoCIebVdE47e0UOGipNbWyQ
6/PdlrSw7ZMpGhteozxNUb74FhFg/7klNTKKb8g9mISI2eUOy2ERwZ4k98kfK6eWn537JgOIoi2w
EH0Z/SsTSqzIBRXotKFgmxNXjZcnsByAhnujkBVARshd+OYjvepoaXcWn8libMP5g/Eoe0zDrXsv
rAx1CefcA1/LsIeCyRyR9gIylrIY6YU6ZxCQvlx5+Exs+6t/7ndMDL+b/YFrY5KiMfFPVbY7fhNg
BwQ6eVPn1LBcrmlm7l+HyPiliMu1sRjhOAEj6ep+kUAZE93LbZed2DRblmYtsrL6UbOTAikhlK0w
RCXZsG5/Ev5CvTwU9I2qrQsmpq+Mby4TEbJn06vGskKUIMk8B4lubwLILWIrynF/tjE+mbEDt/Ni
kU465xF71pQN41YesDJTtc0JQNbiuIHv732T6/be/VTeTeq6Gnmp5kcvbDwIPVBBxzWvw9G4bmo/
ws9R9RkTYCOLpobrpd+2TQ6fcm+VO1C6sajV4kvnKno1rmFzVU7zw3z2d/wlyIgQ8UAZkO6XhAxJ
UpbVZJtLvk3n8cjSCAEfqL1JZd+S16BLdEB7LnW8q5u836Y6jjRPrcFrE5dZZI1N0NZqAXFbK+Z4
hdg1st2pZ7KoTu7M9NgrzSIZ0Tg2TJmAX/6VuMfQc9BJ+JvDvv/syXgjdDltJXjr1DdxpFTEyBEG
ZFnN4LMxB96yi8bSKiqgT+KyDisULJq+k3joIydCCuX5RPG6DxU+/xYKWI70WemH6tPNaSoxWPbz
j0J7bYyPSlxdPmMLi4RpHIhnNckQ3xV3ffZZmgL3hzHWwzjnhPhdzV/ZqPRiuD6s2L/KKNxHOTpP
0mF1iyLzl6UFLJyb+xQmxL8yKKxfk/6i4pSV0HxrBPmW1eyYpAd0BlKzz6E/mtjICo8HP0CwXZBP
YOLEDIa3HB29X+xpGsXmp5MIWV+U1GuFOyeTCiwuga76cFgDQEMexEQEqmmk5sOae1cY9iegVRQ2
hhbHg/4I6yJ6aA2lDuoL3nJV297gXcHEfnaPvAU7TP6EzQSucTQG6pIOo2gCBscT36uotUEqSRm+
w05KzJ2b1FptUzk4+HT+R1PLSF1rcXzNTd/L0ZnDl1ZlY9CjwxIE3uvGlArqLFZaLg2r64LIP3oK
GVsaZzxds2Tcqw9mULmuipls4cUOile6ej66gwHCSr2ZG0YNkpSQggBVQKyMmsXFKo3CnewYnob4
ARJwu+sxZNg38sVs839Hgf8pX7aGDpJtRmzpd16aBeSUBDWavjXdaWCKBzZO6VYqqJK1ZXPjbt6o
nZfSsnTTdOyHujXT59AJmwm+iunSnJlZ7Tjy+MSRrzvtAibf6L6omkx0lRbhmZGSsflqXPYVPt3M
BWvqJ7X7r+A4TXOfwUSCTNxvc4zeZ2N5uVDK3W0+s0tmfX8dmaqfs6sBbvM0TDBiEvOQqC9rYRYV
E/SOhVhq6Uf+2enkaWq0a4Ym2iPI4JBcm8LsAPIJYyR+f2r0u1vTV9noGBct+eYgQSa48VJ023wU
y2bpzsBVzKjdmaZog8jYruz/ERIR9GNfneWsiZSXWmnVfFhU9qRlFKEM7/ojzW0dW11dUWybJWxI
wu9zczYtZglBkO4ZhoyhaXRPGUCTCRB4FDUfvNxJvlDcWqCkJcVpZzSf2dvfdqxnoHis0tMZd24K
29HUwKnHwtw2+QH29xhRecpbikYAanSe2f9FRKHNJSvSJ9eSTU9r7CJpKzFUCJgCZU42zQUtrTRp
0jXwA9qpfpGSGLLFYlR8h+sZVzkdYdSUtvOOcMAe+UunKApFufLa8kBxwtlBbXon9+pZ2giKgFz2
TV5f2GpdvDB3HnbDMp/uR5/FTi4XMvfQHkSRI6ULitIYXyj1N1KVJ4diQSMUJjTEkPgUvOjnPb1v
Mz8Aw1WNjFzi0esZKrp+wQsdO3X/72PuIBF2HHK8m74yCQUqJMbgFBStV32upacLge2gXXYSPP41
LOYG9u91ixC0WyaGfU9a9KdAybQUML9dzdS4glvLMvUuTYjhJxtKuk8hHViRioO8hK/wrT5xPW6Q
z7KaW/dL9sKsEfNkeKG4ACCtjPzOx8NWeN03TIOtu9ES452M1yKR2R7/fDWDTE4JXmO8U6WtHORU
mLo7i0IHILG5+RNEmo+5shfvHAPt9lyX/mDVYz6pJMx5kfdH6kIIBpHPkPJ3xlQ6Y8Udx0IYcyr8
phfX9I4rg8PidHHQxP9wctypQdy/LyVgSBecyFmZD/iIdxpfi8Opvnm6OBlbaeTi8YHT860Mr9Ho
9DHhgEsU5TAz+qoDUeihZg+qcFTL4MGQN6a8NANrU2dHKSdwiRL86wI3795aNhbEkZoaxUV93g0J
Q9160oCvjiXkzuS3krIoFFdoE3JP4D/1bm5J8YBqWs0ZKEfp5WB0ahLVLP8fv8Ddxn0sWxZLR8Yi
XeY2tVw9JMYXgU2GNyMzXExhhnsjlyBX4N1KtwOyjCFhhRVwMCIBiFO8YzQGS4/8Y5M01pGAiDM0
9iFUyv0ijbUPjdGTaIj7lUw+02qRypAsgadm36n0fajQ5XJQzzoTD63yxOf47ll6QbIcK7tTfiWb
Gjdyz8y3FDBPK791pfJQ8Y6Xau0DBDZB7YW3mDtrbw62JUQbQfeUYisWxpbd6jh7N6bTIxms7r/s
KFXlcSGfdxml90hXFLsFfYoQoPRiaDTDgn879K9Sepf+sxkrpt0O4RDlAyGLIY4IBwT8SeiOfzql
uXq2xS4utsq8pnK5yB5YyyKnkD179+ZI3PfvFqICQMxO5aYLsSB/kowSFw+xxgIDP1Bs08Pw7IpB
B1PaFPWbsxSLitdkLfy8BFDJsWTkJNg1J/ek/4dFLp7VX/tCeMCh0oA6hsni+zHoRGLJ3O7Jv+y2
4RW6m2v6nC+8WW/6srYrvrMLbzBprLeND69h1Hg/+o3M9XYtCzyStciMAi3xV6scjwcIr9laXOBk
jQWUkwZHkOIgMWMsmQK0+8VOpUfMJywzLS6A7pHrWfsmCKanJEMVFPEouklCAQmqZMMfzVdO6X+K
Rlj9EOhUbu/3iIrAy7DbH0QYbmfpRuwdYs3H/yo2YhDuz5EQn3YAfkUGjB0+aOq4YlnwbEBNkj9v
3XbP/IjKmaAefL784CsbPuh7lAWoCheyr0xHqdS3zizH7Yr86l3XzUjkVJuB7ugzhyNNHJ5fR17G
gTt1IsHdIg3thSFNP+JqkghZdT2hmQ+UmGiBYzWgZu7QO+xFssLeKS4wi9iPp2K1C1ZibWM72SUs
1+kBj67IcaNs0LHjcT3ckIe31QIpCdLA2adPreBBeFQfZGt8mMKZPZXWnaZU4GUJY8jRGweJecW5
1c4P20ciWuLbFJQdtEArbKEIC3FBNBqQjtQX5GZx4ngHS6jOcqrK6CbLeUA4mOThwRcjCvZJPoYB
ES/lra4QSKv3keg+vG06Y1hRP0Eqrv3ZcJtQRw/NaQiNIMorrmqT22vqSpqnMgZ4NIsMSO05k4lR
c0r+T6T6/OCfTa0gwfpEGO3pj3Bujv9PghQocAwV7NzwI1WuLCtTgWQA8kFuknonsEosrToIAtvq
Qnzg7cVU5+TVccmIP62tJw4kVJbvXmAQINFyeVH3x/tdXylXyzOcrnZOyYMLOQy/yNJHpT6IGfNf
6B4lIjdIzxkg3vNQ9f1rfPJHGcSoXzBM29ccwLZB8lbgzUyrDSid7Pv30VufKJbczV2SNVidLdWI
zb9cZa9eJS4I1HuNVFtRDwQv1YfAl+1w4ellO6GFdBDeBOhHOn2o9iyepKFcEmDkK7KFZS3hOjNH
g9LC9YStIEYHhEEXfV5u19cGA618u0Cbq8jeWJ4gM1/oGZh/nwtI16a3mDsv4KataFW9fUFpHzUg
OJdhz9DJoeoTti2mopeAN+3yD6BK/+DBU9Q0wah/62Aobs7zZyKJtqOFSO3WNLaumWE2PGAb3SyT
6B9rBwV+NNqmujL7gpHo5vIUQCi1Kg+p40H2Iz1UvqBtl65henPJa4s86vxqq5beczex6DLdTmOI
dOaEgMQA/S53sQwY9i+gfoi2sPai2BIia+gNTcOWl3zpx1YvcIMtJex9jo1McTtsMOW3grmbcNFb
QOX8yQHqhtP6fCCJsxxcZDTRkD2bU6yKW22xi4DKyOz0e4t9rr9CRvZN/Sh6+rRWNYR/qjNkXEkA
WCA0kWCU7A7RxuUd3gCLusvO6BDEkydvBr2CDymcFl0bUV7bRlovQI+kUVqf4aljoc8rHF+aKgPk
xcQBBDvLSpdJSNw9+8xTPDE2rVXheHavHU6ZFD408LIpigQKua1u+ZvoZhU5DjWAcy0X1C9KFP3x
LeqO3NOfAVhAXPmUpgc3yWXzyfYUYsHAhhdWDN7KKJXbJMITVkaJzqpCzkcba/iOWRr96na3VYbz
nOOmcmL2Xwy2Iib7awM53yJx/IrSFU9px2n2rqJLtX+XGYzuBvwUooFVWpij7GK+TuMcQfHE66nJ
Zs8fHITM9EvnltFT6uyAfnq3r5YJ/lKiBgQV627uYwQvnxldalzfq5QpFJNZwSZZOmNdg5eqUReK
wXpE7RK1y9XuWTxsU9ZzNLsmbp+7F3U5Jx04HjgOYSwPSVJxIM7FqNVUO8xrR4fc6JHZI+kBz75J
3c395h9kBGqGWYqad/twlpg0faFe/QV7UodiAq7afzlnYY8uMxidvqS9BZBpGBL7n3xhPodNEn0Q
eYKL2dvnqOhThzLSi1+eWCGyDDs22ytWcvsSEKxqteS5RYVQPauIlZDlUlon3rorrG4O1omQFHpQ
OcmkTDVTXZZs1Fr2nKc/yeL30mGmiLxyFdA+PAJdAqCZEqZvxFmNhmfnhZD2Jv8xDqKH4cwNOYjU
UA23IvrqzCMqD5p/yCeruBm5wgrXNi0mXgFbUQ1f5kxOhJouZB4bbtPDhvh/uxHshA0Hw00Wfyq2
PCq71mBItPGHTzoA4xYyVaTzvIcu/q57j9LJQBGtq4LgUJZJBOD1wn18UH+Z99H+/KxyMiVZuhCG
9sGrBDBAmPNjdzQT2zvgl93BBU+Vyb+ND5PGwRLcy8QxwPxwRaaS0I1wTCdEiets2yAAfSBl6ybX
TX4evyngaEichR7VS6IJ4BA1rZ9z5VicoXiyoIN3Dw+K6iQ9Jn1lR/CTKqACgNLT2JqZyfYkIm7a
yBLL+nxWwK/YO5gNQxkZj+hq+5ScXplV5hRExEMyw7EPXGKFlLAQ8Guu/akjXdWX+a74g6iCVltn
aFPGhjmLuWogyghyiuqc1gENradCGCUwG8nD+D2UdrK2wX2dYEgDE3RGK7BLZzQouDiv+ub67alK
0918LjaaF4Rf/f3xkBtB+x7eZfEJhG8SSccGCrrUbhI4fkkwCYG7ErNBDl3R7uWikOtAwhRK1txq
v4GkAi8yF//1F7YolY4gBmvWE728KCA6FUawVigB5Vmg0V+5v4BJskyhXNngvp6ShAIXe00vJ8MD
wlwbW0grEzZszAUkAhTyQ3cRoIzVEoI6clnuCsI9SnSqaXsU2CseMK9rrUM7pX0YU/rvWVHDljpe
Kzz7xhOXmHiiZMEJWmyWUGlvcc5kcyH3elmpfbp3nQQX2c+Q9OmtYZeW1iN9n5pGmVxtCWBCmNBK
d83GARK0YJcaTViNYEnvclFzymIBg331fACPurT2y1M+XpVzmlRknwtpqYYzJTSVy94eaMQF0mVU
Oki5WzR6ivmriXrnZxDeSeArbKMTOZNteHPtPxIYTG/8Z8puh69yGgMPtUkcQ9xQE1b+QH70CgeY
mj6A5LZyUnGvL54DuoOruKzwBfv8UqfLTxtcMpQo9ihsn1yjmrqGu3zqyqW5Y747vUVLepIYycab
wEi+rD6erS7KPmAng1QIAaKK6R1mLrMEGep/vRjfJ+GvMGbTuOSGvHfDtB3QFrx5CYJquOTJc9W8
HFJSaM6rp1CIXFWtHSpWcA207EQaUAKScExM3nLp/LMqdCpxC+9WuPZobnHLsj6bX5RmD/dfEmdi
eNlPugzH3fWeOV5+NK/jsQOy4akywrbil14MJwtxKMLGnFqE5wk0ZM2D0Vya/52/xVMauhftiNV9
KX0zRa9vz2xYA3cDSBQ/P5aUvRU3JxUwLwkXpPROIfKttwkQcEzZsmq4gnGnvYmqafH0rf+nBcfl
heOU8AMy26wj7u9aCEmVPulwuIu9jQ2TXiXG8PnsjK85cboRjAMrvyUiLhKRFSzMx8IMA60pzMl6
QK4R5g0oA0+KkY5NZczbTQFGmFn5HPANO7SpmiurZA8ZY2U5VMTDwZ39OUp0kKaYWJuvYyTT1MB6
YZHGUrKYFRIB9w3xboc7ylUZb2scAA3+7X+FWumfMf7bhQtWZKDb5pJLMpL4VtPR+83lWbSLoKBO
NfRtgpJKWffXZBNZv/YxFk1UQTs3hvfv+5Q6BfWzCr5r1mTbnHF1zi+BN05Dz06FcmEGft2n2SCX
qusBPU0vX4puPkAI4TE6C/XDyojkAb7aT6vgYCS3BaXFKUUYVojVxVC7uOSioLPPMzmPiXnsWpOR
VN+6P8TsQcytfK5P0L3/qfw/zPq7cJg/1F+2z4gWEXh+v+xebqVB51gIpX6Y9fR0O8PJKrul8UCC
/YkvuL9cRgbKNZP7tz/YYzf4DyCjDsjUyOX1llol8tzUsAw1Yiio3QhBxRHU3f2BznivbJ+2r4Jo
8rW5LexkQ11K7tukdQY72Np1lFiXGTAinbFSiVEaESM4bvdjVPDqvzQ7+f+xoHhY4vtJrkTZHMfC
cxBnwe9Aike9Ykp4OXkYKEh9XWy3L09Tc7jt+vG53vd3YG2HEyd5yBIm8ibZbgQeZ3v9kfZ2HTK5
hDbsQj1WcHnklx59R3G6IXKF7ZSpXNglnmmLuf49mIk7xC4KTtwDnrSc4FCp+WLMYUxVGmYGQhfx
fhe9rQzdfArHmz13OLoB2ekPePSajngEl2/BIxN2xXzqODDyLOdKaYTompX4A1pvxi+f88xiFCnR
Dcc82tUuz1jyjz1EFw+PlzlGsSNdq4e01cw03a7pNjtluqSJr6DxFYLq757zoX7xGDq51Brsa7qJ
Wg9n6p8wJf+iVNdGPxClz/G6ljyzLPg1OIVMKLG5bWrLnEWZOwzKVCjVMlfzeXhBaf2lq0RbAB0Y
8/1iSDBGs4PTouCGhbQkwF7nPhyxgr1ptOlzztpWNt68s0BdeyUP69D7krHeYq4ZpSSai72shbYL
AO76af2uHGven5Tiwkmiyx9SheHql92tj0a1fsa2g0f1gOA4rKey1DpXH0fposWgZ5pQZUomDBra
/DZEZ0nRayj7ZZF5i2qKUV+M4yBr4beGRW69s41FR5D/lrOzmIqvGlY8CjWGHL6Wa2qg5+MnlaY6
Ub7XVdeaAOIDopGOzp4m3NAqdtiIMDOYiTWINIuej47n1fOCJExlJHm8vR6kj3Smi+d6kPypuslw
IoaBMW3sW/V1KcfVw3yTLr0Pq4xjT22Csk935iFHxI/hsLtU38aMhm6zyILD64scpavW+Nyr7Gez
oVk9Y0k5hgsVM1hYCMC2mxoroApXpho3+d465T9mo69tSPLohoutKB0IYpKpPZLeHadsZz0BWg1t
0xMXRwB/097Y32gZEYvbeFXokAx0OLLES77FrICDqpOh02ciA3/Cw4vxL2fzadzv7pyYsjpe5plO
BbeBbShVS/pRJfWufJmqL2Gn23wZU3xtYrIY+HYyeCb7gG+DmKF7XCSdNOnBWArMEeQH3S1+dXVy
pIN6YFRhSCl+IrH25IgZ+LkHFd04Q+2mlosLvdizbK/I7REtwj/CTKGwNZrZvkIa8DxDwRIDzZV4
ocdOtLffI7lf/fxXIggT0JgDlIQDcr522heuNYq1AIMuj0aN2eNlK/L1pfWXzdabSsp0jVU0eVQ1
+G/oHLqJ65Tf4KJzwQ0aGy+7AVLsHj+cehHynHWm5STUDIZE2zHY+Nv1IIZ8F4CAIpwK3+rsIeeQ
pT77I+4LuRadhT/sKRPxESKwNMclu6GdASPdQPOKhuUQpJIkO8WmouUOnyRfERzbK9O2hq2bhlzL
atNFOv7knsVTcGO6VyBQ6vPZqMKL2fV44+XX2KM7+Y3K7/7QrCawN08o3L8EB9A391L7Z7jrH/3D
xgZdbi1kyyT2xn1onC27yulM39UNBOfBfDlJP8MgkXhP6mVvyIHl3L+lxdW5Onm6PAYKMjOKcvvX
CtYz4hEEnEqKELTHVMAxm7D3n/mveT1oykTMwcPMywa9LaPyBnlj9gwSCr07JeCpr3hx42Lx4eRg
/0jF/yYfTfiPRw47FINrr4jEdJ7DIove8J2/InJrqb/V1No1nQB5CaxzqHvEs/tY77Vz2chh+EeK
eIuE9altBfhRFIcLMG0fgpEYWm61ywXzgw/ZOyUftfJ3apQzAGpHoTgMuotrnnyy1354CIeN/JVb
u9WEfkzjksJL+XB6sLM51uXFmM5oeazyQlodv2IWYoB+tSTg9Nw7vYV5OI+EhhSrdIvAsgOVDR7E
BMy/siaG++kqgPCRySYWQv6qBCR/op6E6ddzcABBxNxON6yzUf6/wB/Sdt4R6l3b38RxxnaUN2Nx
wyMd+pi9hoLbNn1iQmYEZKxrCYIqbyw+JcgGCVSKr1wWybidHjZs8iu1dwHJOV3djOXKjpHAzKAA
zrHfhuSiEa+z6JsCm13KwXAFe/oqqEhOjddZahptWVW9R9dAEI6iJNfEoASLq9tq/6Vk8i/nl5Cj
0apzLTYKkinvuayoex0U0cRtSN6vEzTONPPbmdNjeBmtJakSGyt8S7yiE92/XoxAkU12EAcThxtn
SeQ1f/J04+puGWSVLo1k7rT+hr2hTwd8C6xFt827eT7iD1T2KFfZuKcFrMH+qhSnRIIJqwA5L1O3
NH8mdlRtzdaS0ldCjOGSsxZDh/J4jDcDw51qWrYbNIN74xRd1XrIfvhwUmtflAO6IQROl7687dt9
fS1YKWu3V2IE5CCWeQbL8m3CIaGkckzEeiOlZAaRvWQnfh9OIm3v9Iivx3wpkL/U01SA5Kh/KTdR
dN8eLkf5nDtR613/tJnmhN7SP7irYfK/k0SpYOob1zxcda0nmIQ1EE154tmJz510vNilclNyzrVd
hIAR/Y8A/YTdmEXZchJ2Kq1AMun4TLjjz8EJd1H7pDBp0aWHMv0eb6CxUDJfq9o+1Sea8yVo5QkR
kPTOivdrUrOy7UwlKXpYBYRShqKKM3sNxMbcCOMNeEIa0B/sMGvYA27oULqjdD1KZkixaBjRXJov
UhoFCsVp8YUB1aioSkoHWNwDaconYoe7Za1oChs0g/QfXFtljEQGmx35SP4j3KUcJ/VOv5Ikdqpg
EVBUL71EvWbPcSIgPBVWAFRTZcJOWhKGx6Z1et1eMQqbXz8zE96NZ+yeIJC6psIeTuX6WHiABUpG
en09nf+8mce/iBIYKF/EO6lndW7lVwhDXUNgvfvki4jfWaIOhJ6k4rdkOU/0iWZTRGwZ1/MK+q4L
jXpYkujZljM3O9FGm1nzpyapriFInRfKY2VI5l8Eh7DTl2wOQtLlfL1vDE94cZUmZY08VwJKuLBR
I1vpo0D4YyG/m8cKQQAHCf9nwjEMiTWO2lmeA7MG6ue3K8RkjpvqLtnW28CIx7m5bAQS9uYQlsMp
kPFQ7TYRcBZhVvMq+HXUHD/YhWd+PHoU9Ryvxd6H3vHYQ1wS8NGp9qbguKRhyMunDtJb/aBEqsy6
C20WdItvGtSZmzEyT+tGwEMKNBlBAw2w+qx/jRex53buKeucLD/+zmCsyZ53PiVyjYUoFnOjJYVi
1QncK8ZpuQcB8AHoiRg7g1yRVa/s7YQlDUNhewBH7lq/IJO8sFTGMKxl7VDK7BmUHdn1Wa3jvOVx
w2IuTspOucCHBMfOgmOP0+QLLdUop6Rkb/9lvTpWRiuZvYqSPf7xpeAanplB9rHHIgHAFREEycpm
lw4CTvkmZG1GUv3l5XFqg536f7rTNFy5APWXwKEBx8LSr2MJBG3Dqc9FFU3/48Dv938aA663M7nV
cIuy9pQ6P8nHp8UieW9eDvI6krPnt4c+Gup7n493WTV5fvv6PeeueSdl6hdC81oy4NB7FxN1x/G8
4hxYQqMV3ujpFQLp5GErgB8TLT3z5kRKfaNEks3PIVOG/N345anD5LC+NwEjUL0jpn7lAcjBtzv2
mbCQpPn0YXYJAFqGPZm6c+6OYi8N/+veVhzffUi99i9u0JiOK2Ms5+239oUtvzZ0/0QeHGlXMX00
qd6tqIJQO8ovMNP5nrf8v0hKvou9jD4Lwh7NEi/CvVHULYtvEhUxiX1NNoyANxPIxObjQMlQEKTq
DDZA8DLK99ZeQhyhm+7M7ps1oXt+QzTo1XW1ysFk8EWcMLCh4x/2+nYuXlGVaraM8Ddpw7ldNJNx
oYKFF6dYZcC4eYxnXGpQI4j74DiJAVwAwIJ4OIToIVPnuZKzzMeemwuuYP1xThLNWwa4hCd0jzxB
pBePS4II3xV3xDncDANJIOvaTP7Im2V0r41aOeZO8KWKXUWma6lSxXnEHyS/NMboE1z4Gvs55+o+
scCXUtv1spwlkmhucunk/AQW7T13G/4fNPSxhLrqYG+1rkzm0peup5hzDmFiCuF4VIIiVzE2UwC2
+CP0Gqe/vxerpxQpnB2rPMBL8PM0BkfSMDNyo1MfYQxNk+jyG3W5Hmx/QH5nm3gAEUvEReUkZkm1
6Qa0+XO73xsmzh4RAmi4ylDyQaKAtPx1/O1aFCXSktwz5EM75SrNtg/NY5mCJjIesOb8T2WD65Sd
w/YV6WI14a6SMAoCvjHINrZPyH/o/pWnv7ftWVZ1DNXR88JyQ+0GCLLCd30h5OpUSJojEIFf9eHy
doRVXNY4PygJXBJcDpmrGfx1lNUTSgOrKyadM7H8X8wHux+a7OR9LQ64eQfVf7NRIzS52nvaSpoK
zvsjA5BD5rdAFPAymDhwkofiViFeqjON693Dq1TGIDXc6Z7P7JMlIXJSEO4xNISrYKtzUviGaF2X
2VP6FCS5PUx69xICMGAyvr3JHEgEtb8ZaHBsshWUv4sX2Even9v1Kn34+KwFpIkwn3Y/6gnjw4kg
TSfTy+JsHMNHKvNSYHvBk4Vn29uEwcuLMj+geiP6gGzfvsjc1LNEfe1xaOHX0i69lB/nhMsv/O7b
/QzwUnfdiqn737G5PvYFKjg14uqMqXBFTbqHAADQWjBOhB3IC5OAuu1QKdvpkfnVVYL96DCHpHas
sdLLBeydxL5RwT22r48feH31N7XG4GUN3Zc9FJc82/eGj/pXTpi077X/bmw+kOikNxxDT+A2IJpr
Qcwmny+TG/mYLsDJDz0HJzFoyMCArJxHEmKZVd0zB5IHt6jvHc0riP0mxeC+A7yQ65lV/JZXHZn0
CahFWd9DLP4XahOmkyxNtfv4FWBvSQL5CJUCgCYyD08ihPHPLIgIDdBK3Jc+Gblj5YHaEtjmy6L/
fFaxDWsTEdx8qaMkC+9hS025EdxNDuMqRqzntNjvTYMcH3BChEgT14L3E67sjiO37AiDTvda15zF
57O0y2odRmsBSKrutD5ChYy8aU6L1UILBxm+RNwesRxd/ZDRlenXUSvnwf6QU/8BN+pzUhwGGfLu
gZTBu7YfOwlYi+L8h50Tp+0G/ZvFl0x0cakeH3VomPWhzKhl5JRwY5bVII6yn9xfJE1kkaFGNJYP
rl6uOVOHa8Euqnqt2Sgzj9bglDSRGdkPYED+WKgPmzUsJCDj9hvg4MP83TT4IVyCCA0umSyouulM
9C6keaEh7tKBnT0XXhjR2awf+gqUBSnKZ5PIsnEMf5i3KEEGOkFVvJ4QSYXqlGstkkwhCmwVkwjm
3aHuayatBKjDxem1rCREwQJQT0RJd2LRfyjelk6a7sB6scQaZL8U/0c0RkN6G9CPuQpQaGsvFt0k
w8FVDWipi+yukcu32AqS6mUwr3LZHV86vMuDQnGrOOpm6J+Vd2U6t48BV8vAt3Qpp5oiyE4WNfP6
DHWCb6cmPZyYb8zFwCMhx4YTW8xxah1Wp/W2aIM+HikxlBcqCDKThC6s9YKSn1FQmjIrr0GC9jSq
haPpJwkoyBmGKqAC7QUKgqoHgdIaGHlPIPU6MkarlkZi6KUtgAOvuKNwJYLWIcS/jfdPyBCUyGw2
F+mrPu8ojLKVwg4nrMtkk489HophGl0gnBY71BCBORW7XDy4qDMzoZtWmhJLIxZ+c83nuVZExRuj
gRsMDDrJGxfBdUsS+Phkn2hT4HWO6n48hILXvic8vB7IaQXeSTy+XyBtIjmS8lEwtPGbq5jmF1b+
u1nVTqr3+O3nkFyRJfud/Haerqy1aiH34Imxcf/+WIHXz29Knv8S8yBm6aWLkr9DryDq9L3zKo83
mh4LcAcMBY6GhI5E6bDAkyDVj0uOhhqMUYiU637arIVkYYBxPp0Psz/dMU37r0wR67QAvTnnv/l3
92k6H7m8w9CwOHSHvPQs4hibdonwvFJZSBEqMUQfQ0e3HHfOAPB6hzEOhbte8zMmfDICavCXGPuB
6NuD8eyTkP0/2uyv868do0XEkF0ic7oKGBoxWcHG+YSihM08+wDH7i6JUtuTZlZvxJRrccQ+UJ9L
DuUJs1Fvnelp2BQMw4czEhlnTch1k9izeOtSMwyvt4AomOlUZmpkZo11cFed9800Gm1gx8LIiWNL
MGW56r5RWQuVd8ZygWJmNo/ZHncQxHqN5xvYhrrlli2vMScRhdlW7ur82NaMnC3odz+2vbAn12qL
a/hgtrM62fnUPMYrACYjZxz8LpZje6RZxViFS1tk2yi5F3AnM9wIOfeEXvzlVGT/AB8yLSp2e8//
2kMcYhHAkX59lJL4zo99gYQzxpCcioSToYzrHjXQiooTsfM6iOAYZKHKODUI/SlZZS0wO8gqO9vv
hzYS/P3IeIhQ4tJ1Xj+sFRNy/gaHw5D7wP1UjsW2CuyRzTUzczWbleWk4FwTEOioj4rGyn0R5VA5
Qr9b2RhgQPvHciGFBDkhDZawafSllXWiRgujTRPWpFAmppGLiPT6/2E0LfhMT12uVS9bboLTDYW/
6oaO/U8zeUAurcuqTKu4qbFHS2l52Br/omMtTfdG4EMMJtq34mIgvRa13Qo7xuEWW9HelJdthipR
qvaciA7X4IFbXUcO4T9+VgE5T9c0WQazzQENMQP42egxRfPoa2ieXiXhhfHmruzGVceY1JSe07Oi
84ae7rQIb+N+JaFz48zZq/P7bv7sf4O5XXA9lK7anNlJmItq+nPc15A1jNzKfoiruClZG1uVkAAk
C418AA4di6e1HuLSSq9SeJh72T06vgHGt0mnOPrmTkDw0QsF9w+ZbJKQLXS4VIaLkOrCNAVyQJUH
WhkiajqeY+IdDvKxEkQKlltxUQYhJEc4TDIlZt29DsW3/sWXhaA/ASYLlEbDXJ7E0xe/E4rQ5DHf
JG8v4myXjXLWBTMBKTlNoEUogCI090HbMpnvattaZJkGWi4RTJKJfvOxWcpm24FcJmHHnK3heERF
gNv9ZJAyp3uLrotxLP0XcKgKudQLUvqAU76mq9Nqxotzh+CwaXJkwI7M2MQMPkYcIggaRndldeNZ
S87WUMt+BwUlZmFZndlbVvHwfCmqb+dBq41R7XXGDLgoGdIFQTdwOQZ6KN6AcfzL/3NT7uXMiITQ
+LzhPKmeIcczhMzSupuXxC2KtuhNIDNKBWs49cCdO9V9v+4Y8OZfgQveuyNVlfF+5zCttLf0ARr0
w3s5bVfLQT3d4PNg8ZCQPPSvA/BkKsUbjKiRS9zsHFaioxeCIS6tamubBrZKQu+4RAsK5aQpoTd7
C6ShWIBWQ9mLDiexTBzzZKawUDVYptiK/79Do/0AZvV9VRmVyIMemR5PtSfcVN+rRwW1aMGM3Xg7
k95YnuJKnY0mZ94njghpvK6SofjrwwGdGzpOKg4Tbt3lSp4/8tSWkO7tkmSfNeA63sPy9UqthgjU
BVtXcmfVwBo3x70rOccvbkOboxN6DmjgSwvdwOyiVEGcm7skUVqaTweAbYiJkJHh8JjWqtAPo68F
m+AdGqo5NJefmnBKo7aCrIHwoKefUJGefyIPCjk7OQ+KHkSZ3+0xrsoNfvnck0jHiZFqsjs2vn+J
4lky2RIXVWU8oE41Pa2smGkiSjLhVyLYIGM5bpCyVDYP+WVnFS77OYzQgXJhwVlaIGshhDBqOyZM
njosvfB8gf67EPqgPIj0wEQCDXvfv5vq4SbNyuHbhK726twnbrmIt1GA+e2aDBhqECOdWpDo4d9W
MEZZtMx2vrl+9ma6gLoVvCxv7p5xIAu9RFB5E3FJKDuKopvstEryO6iC1J4l7xBrv9a/rLfgcE0P
Y8LSIVeYsLcSg7UWkioicAl9P+xgV/O+mz1Tdqzv17k6zeabvrLqJxAU3wabavvRj8hK9hQVO5Cs
gHz2oB+Feb7bLLR7pTr1nEl8F6Up3qVTC3XXvdrzxfWenTWXm2UJ4yl1LYbfRSzXo6TbXC4gyOMA
lCybFCykqOgd2V0wScYkcNbVH+HEDampzA5lPGWgWqbTJYvNhjRTxWgUOueLUIV1JHvyQqcOyTTU
e7r+1yJ8y3ltaKapOAJCVub9Ue84c/bEgu06dN4O/YZx3FVK/Uxu8wDl9/ir7OvbIL6Rc/ao3+Ut
mNFrYooXY834Cz513e9ogqesqoou29t8SYUdirtLWJmrYJgEnL3ZHlGsS7nW+SZmZLCqlanv6vrm
aL3PeO94OBHgYiVVDm0q2twaTrjlgBgSA2qeMM3YGuDBXuKsSifg9Up/Ag3zH9605P0sCwfmjS/U
U7cgTlFs5olVleBvApWOGx3iN0BVjIJR6UJh+L3bOSfMl+fs7k4NKP9fJ1Y1miyvAnoSqYRd2Gql
CtsBGYepybYP/0nLL9noKCnu5Cqh4x0Yvo0zqs0Bazey+HycvYC3IC9TUfNjknF6gp45vVZFTpTA
U+2Ub34DjO+aU54f1sb4gQqnoGa48CdCFjOKV2ApLbmeWPP+FLvfPvouZxpLf51Vhx+WBzHWPq2C
DFP8d3bEQuEml3yidjSS73LJsseoSJqfKrRPVsrqKcuCskJ10I9zBpK01bb/TpIvucSlCi0vHMV0
DH8sA8eMCcuxK3+S0EFnl36+oNIYyZqEWx/veLHIfSbY2iJ+v7Vlso/gVXl+DXIl5YDoD89vg5yF
ofYBqeGwTUD3Kd/DQoCSZGGU3kNMkDzwFw/yU77aqr8Qq6+9jbI76v4MGRMc+ZHnQBfcofuZY4JS
9WKVJYLMgxfYlth6Nparq3vjpbvtMyUUV2Yxly+uxcgj+LoDvL+6Wn/LEAKijoxDxjEYd/L4zxlH
tMcnfKWWuJ6Cv7hFSt0OBC5th+mFM3a92vt2mhP4kZf7+O3u5Xt9a+UworxK8UJpyV1lJdt4kqw8
3xGkjd5+KXA4EYPO5gvwzv/2t1H8sOc4Uv7UqW70bZFETe7OOj36MQjUa6hIHhxo6hbuyJ0pZ19C
lPKpIOhUUCXc//BjvDCF7jcWCXm90gRwyKiw4BBUS1rwLj6sEgVyiExnghvy94HYt909GWMebikt
4UHty3AvX8Ilrmi+U5go9ihpdFNMIHfUufmBnpr0mrq/azqaFCKfVhXCu2DgpjWqnBlThKWs29qO
AoH5NJSXK4jnT87gbzz3UIFfg2EMJdSxzdHALj/Evkn+dBPuQMHTxJ5mXKaWcIi8ZAut6ndLavpU
7xkS6oNRCOyyXYcDvw8y5UwhHCfi+9iAFIPYS8pKoZLU86wVWt5PUalYbdOeV3jtGvYv5vx3tSI0
45UdunaqfUqgWKEAjhufBzNg8mYcbeB+nANvc9ZYVkzjRUSzo1082fy2wLGc7+voyOpRahQ4qo/C
e+PM5xnNp1FK6feF6TODxMEfeAqFfbpIEGJW++ESdZsGP2GvoLRz+BtGN5ppNiOf8OTZeA+EJj+I
0uMy0xr9PCzVvn9/LaI4nLpisjamd/GydNsR6Y396E4L0BrmmtolYxDlfxlxPBTjV+c9LTP9cFfC
isq67S36m/yPaz9I2+9cXNGG9q5BIfleSe+Pcj8dB+avL64ZB7VWGjGkc2+O1LKzJEpZ8hVj7LXY
eUzG/tNABnQp+E52cSK+VqpMJW9jjz55xutsocFii95IG6J+tmS5zSTVX9mbhH8aTekmaXdARIRs
VHuqn5eDMc/qjkf4gznHr+R/v4FUAous2YyI/NPzyeQEnniFPLRABFs7ohGi91VAMaqaeB4rS5yM
qvh70Mtv1ExyMMbwxkEUK4HBJQZxhd1D1c3MRgubTX6npkwoiks58MEFS8pG6ZPyGe6E2w3+YjPX
TtfVDj5FL+zviiSgLWUMJtRrxscb3MKlFtWBsY4V7iWE+0DDCUcjDY7dkD9+gh4C5AvJL6KCwVbk
ju413vQS10ctCsmsxxdAoXMBwtZcy0rnl9/7ylXn7pEXvX3SRFeaO1yDvvZ/qaXgJsuKuZpDDD9T
V0vV4HulWng7RIzW5u0X8q5Qh9cagJoNvuZFWOM42Dokp2TwZZeDi+wwRt06Xkfn2vxZktPzaS57
+AzaUQajNshzDIYEk88xvrSFCcJFdVbfb49lI2MOfzizulnd/mZdF1su6i3UCs7ZtK8KaMhC1Scn
erO/6FkFrDPoaRfVXowFgPTdP7Uxmp4epNkfM3eIsUsA6Ia2G3zGpL2RjNlOSpUlbdBBWjFBMaxC
tu3uLkSeMAjOoiRT6B0RBp9epKnam1vnJtWdOBAkMgZNV/oStsqPcOD4OrzUeuOBD4/00QVi29gJ
w1x4wXK58/Po8CSfeKbCwQp4GUwLgrlOoOYK7m34Sng51d66SvqUi5xBqMEOe87Y5rpsNvPzusCs
TS3rgq4fAYto+9PD6D97mMncR9X6j6sXpiTaZbjRXbvqbaHQzF0QWfFx2N6sdU6MCalGv1maHRU8
hKP40QAzLD8c3FeNV0qWCPMMZ/YrYygyqqGSG8IjxVX1h5DEmWNgUn6EC1vOmv9m8s77MVpu2Mjb
tF3nwyjpHwu5//zQmN0m16w7fIqsYY7Py5trmtJPU0J2DmXLu4Ju/Ru7JU3rtub5Hk0t0HWpjX5W
piSFE/1C/+z61MaCmeNoG10Azc0WEokFuDZB8lavb29nAkyvP+hbWvoerv5RV7dVJ6wQs6ShViYK
VBP1OZlo/GJ8QumGZ7phMXqd3lkU5sN+783kWVS8z50P1dFlF316yRFiQH3lQFpVXbQv+bgbEkRy
2jCbJFS3PspwPK51JaruJjs5HcE84pX/uorR3y0H7/OAcW1ck2urillzd6iPF0QmegbtfOfmSPCK
DgpfUTld/Gzy9bcC8rwzekjIJhOnl9FSpc7iJFO8nA3BmG+mKjHSxht0vDAM5lB5AT8DDyLRRyfk
M4DXJk2wrnY5UCDklo/yDBtyTbLA0PGS6Pc7qtRXXacInnvrS1SE2d+6aAyMD4w7Kqpf3/Ew3DWm
c1AqSWjVzgEBSk99zSFuplBFh5GKGkoDiN5UKoWlrNHiv7AfCNhJTOd9IBrX/Uv4+iJGb0ZEJjRv
RvhNFZvs/9wFUwe9luGmAYzddWfSjcaU9CtGXaZg4+Kj64/nZqf67fZmrNkLwHFo1xcUcjN/muRj
no0MZPVwD5DfLEWdvNWbOzphq+GqS/K+xNMBSXpxp3G5NWkMn+ymRLTRaMd/mTXVMo3n0xORUBJe
KvHVNLctsdxYO40ZcKyUHsmo+26gOEkbfiPPitzbik1BI0eXsoLBLPeCB0VL8+8b3SfwUfJzX6tK
/6Ny3hq0adWZXAi8J6ksUVdLuPhPVIZbNR1mcGmfZmJKjI3dWkJR/NItSEIqBFYTZHLcKbZd8NN0
1vBdR2sHMmFzxKl7EELSHaMfGR2Qjl3TMMmi1f4eLw9qW/wm2tGqJgQq645M0UnQxoTeHLDTeA6c
2we8+OatB8a1jyapsOElOnC5l7R/DhJT7+YpWLqPQuBgjkqLfwn7tY1v/hnM3ShzW+fIepnxs8kw
/mSRRmtsF/1GCS01LQ4LbLQOJ+y8pC4HPRuxthjy0j28zYvt5Bf9w9oSQOWGsb8j1Z1gA1nYJU1g
1/E7yn7ag8OqNLZaOG5Jkrvx+leqWn0q+VJsUdG8JAsxDjFuRBvUGVLJZy1RyFIHMYfl+T6nJKdV
2OwUgsV9JoJ50QDW47xsyiP5qTVwQOqxs1hG/iJLnZBEIWKlwtcfvl0760mBawmhq6TlDu+TQDVL
tdKBv0LIya5OE5O78jtqCUxb2IiPWfN3y8cFSQvPZl0w4yerOUTHUOBgv021xACdTn6U19vX8xTI
r3Wu3fpLlQpOTni2AGhPWjU9I/P86F/Xeo8A2m1XOzUPLY02w0tPc3JIpl8gdr2dAhL5l3EyPxl1
TtZ6pcVmLjdBnWncvEUgDoVW42t/01whb/bjL1BraroNJHhMeI0ButrexPUqm4NPLwc9UqBvX9ni
vMx6/sXT0soM3KkXsedYJvYkdHTGHFfqMrUbQxeDC1hBCjq0B6ptdQ7YuaaGraQRgOHNoYNMMhLO
FeNp5uVRFGvK3f/KBQhIiBo/f8dvaYURBqkKPii2rkhx4C8ru13uWz6mb1nF9sApu+InUGUDhvfo
Mj/QPQrjqcYRoTGUsVxRCEAsMa7vMZycIXAjhxLEq9VDCLa/WnCfEJvPm5kIfEOkmVncimVOZh0+
vEbuurhOWmov0H+VSAPCwdyBqjo+qjS5pxObQJBfGcWuX17wr2tltNA0JL9F0OoNaMHQueAfjrUl
IZBErYmIZ06uMhVjD7QY4lfUNqZgedvPBn7E7cO5dP/6mhO2KsyjN/LeeCVwOxmWblO1/iNewPQE
jLYYHHstwcw4RRJ3T5h9kBkF66mRb81S9V9Fu0/3VbFFIXMc5d1sx0JZJ0Jkpyi6yK2QvFuyJLPX
5I94AxrKeTpiFV5nvE5wZ2+Z6ZX/B7gZvkHE3bVEvdCHkmrV9XXi88nX90Eu4F5MfqkUMZc2WA1X
e7fowMTO4TKVP9a3tkccx902FHjZDbXsYFLXtYAE/hjeidwr7DoN+bgQ72gSOG/0RLijyI8zejnP
ccBDLe9B8lvrZ47txkhasii4/dc6pYzY8EsdfCB2fVvJlv9S7VVDP5N1izkpN/3p+t5HZzFSweCw
zeYwzhN2tbGSgRz+oa7KEmlrXbE3UxiDHh774YxI4mpuf3v4/S9Zhkw5boWeArU0l0EopsPbD7b/
IA6wOC5reIcVqiUaJ+EXTRrWGcOwrUeTIhTdt/EpC2o7Qs62yOirHcyzdC2BvY9Etyll3XyAmhfO
WMYNlmn4vNLJt16C/qBq+wx79vQTAcKlHAbEk+kigQOiqRrv/1vTUWp4RiheRypMRfzer1XcSI4E
lj5/JqrW7oZAlNuCup9ZzXs1dRBSt6IiX2T2GThGfH0BQRCBDNWbCD+7fZgbK41unOnirqjhc649
S3BmSjuUcKQXTwEnQvQhxLNb5g9IZHTcIsTaHW/GPI9gvulUBqAGboZavJPFJ8uAaAbvP1LNRBXl
+OdR4b1kuTXhbYMwjVMRGSyKzNEBLDLe+r+gnxl9ZUXWmDCUEUkRzZIatl0bkcS3XfQqsgvTPRMk
/GJZdCHdbuFHsPnRJsfv9XPbPCViKOSlWDsj6n5tGxE6rYJN6ZTFHjaXM+xtck+cuBTFw04JYjoF
p5NPzI4Tye52CQXZr/mAYw61qpThenlLDTsMhXvDF/wet/iPYFcRFKhgV8GoKxv7BEVadJ/zlryb
/6254YGk4F9xOyambQtVEmssfxcGQQUgTiWdwlH18UxifdPdfb3Icn+/IhKWlzuRko/GhhwP/gfz
zxeqHuVeGI2P5ElNjFxi9Xdp6u8+yW4k1w+yJzPaktr64rE9oVpQ+RWYFf8eu4kvfqmpvPo7Muii
2/NtPvbhd707NnKL58CBdt7gybMQBpJs6VJjX77KZAULskjFI5/eiVxMlug+CGE7UnDGuorDbxJ5
6pP3TopMxPCmm6LoFpZA1lcviHGGXAmHQiO2QO/pENs+SVysnpuEpCk9m/gSMYMo8PhVoaQJ4an7
DHzFuuVS2V3vaHFitNc/8xRYfvIcyGv6F/IAeG5EZeg/De1fuoSgWkkfPR3URt3z4d6sn5QePojh
68OJJBxwWO7TPwf0nnKv0z8gmgBn5Np5NTFMJ7OlFYn+E4WqWRB2HHlbXFlCIrVN5hRl0iwOWobX
PH5Kc6jUjSyMVmjc+PNBHpctJtUU1fFdZMt3QDqCY63Xf2/y141M6CT+eyYGgUnXGs07RQbaMblT
G23FuxAPF5wTHeWY2TJmbJ/MopWeqh34hKP069J3DCz25/139BHeaEsARybTUy/+odhoQmLq3yxl
/NJgGvnY7hqsv0O8PFfPwOcHT1NXaTa0htN3zHyhFuk6ZZlNQPMKA4BEE689XB//Fo6qTX80Yrvn
gkukOoDRxwXoAoz8Ky1LMPZDCELAqD4aHrxIBRc8VIri76rGwYek/Natw3y8HF6FylGzL86mloc3
XY39NW5vfB3GaDwYvoZeJgdtIkkrUe0EpOHbCw+nM2hQChTota59/AuxF6Ix8J7b1XxCt2W8u5K7
6iIjmB3cb9LQXunGasZoHPtB+0xtuzYKVJQKK4D5sSgVq8Bul2Ssan5SBOf5oIDiqMe5nj+fvvns
UAuACnoHTeNFwm+f1KE6d2ngEqXV4WUS6SxEBqZ7PfdfmOWYySMG51xDtahpS/Z7Y/WPmhego5Cl
sRo9BFDRLwfI3fTeHJBkLXsVKyWRs2xt96UQIqUoNJRS40+MNChqvJxSVZV+S5B0Qu76kTLIMEjd
TG1fH2N+Q5h62iSMeu11ZMiT2doPiMqbUsjT4A6wSzMUb+RwzzoSjujo6t0U4UezhcS/oZxzpuG5
LUgcW1cZgiOUNUBguTJ+PW0gdCwQfmo6/H4SD6PAQBbSCqyB7Jbl8mhDPFKvv6fkPmhat5m0+CE/
M0vMKYr3W8IfDc2pWBarXch6d//DrMKT14ADeNfuzXVe7685WqJYJisQvFygrmzr7PPTGDJzNvCw
oKQQ5Yh/HjBErQIAGiI0qpS+jXg60mWAxpaQYlGTbq5SGTc/2nllmipTjyXs9WwKOkD1Ev2cuvjW
hZ6bi+E5Y0DAU4q7Ry3naiOyNQJWwFMlQOLQnfiY9VTxwdQ885i4f5Dnn/ijxt8ElYD42Txtg5WA
RoA/3HgoiuGnkiWCdeYCpaT300gl+AYpvAbo9PGPbAdJ+DFZUh5VFVtPRGhB3jsLaT/fjTFegzDI
jGj9y1xsZPxSZL0VeWj/o9KMB9E+dOHGr9CDTnl1cS67qvTsbiifHfDyfI7OwBUhpPBmeybb5f8Q
917hoQMHgOBwEZMtSfD1Ve8mUJqkdTSCoTmf2AHVmUTUt+JqMI2LlgPMZ8E2xpjT263+umv+JD6j
r5FYmqS3CtDZ8CY7kGEyWoAfXfLRmbsMg6UMB51b5O7y5DjvEu8QcHea5kRKriC5DiwY15ghURxy
oLi+XTqBGettwWKiqtzmT3FGJBvoD+N/e3yd3BrnXYeFTi+HPeQW155ah5qZ7trajpENWAmXTXJC
9RjjohF29trlgM/lmFsu+qzss4OnAopAaRqKEuWsqex0GQG+vQtPsZXXA9sxFXQX72YT9eFgAfjR
4SgBKT/LgQJYiIicTNXGS+gEbZQXr1GN9OEgoTl+1GTie7R3J0YV7gepTGU9x7iAA4YYdUeEP8Y/
AZrf1E/DSESPg5CBwSpYAmRfVXgWZqYMNdBVy3d3t/UaWLQT6mA0tvaW+5S0IHZ6NvRc2GdZHvVv
ZqFoE5m9mwSO/5s811y4m7VGXMzfNF9oIN+xiicc3ZmhAneuVqzEXCkYkRqwmY8jvwuHl4CUPY2E
FxJGsdlgDN+KD3L3wMTMojeKRVi288LWC+UHQmgXZ4ySJkAHzdLFI5Bhj+r45SBAhLYdaejlNo1J
3ZYJFmpFe1Hl4IrBJThRxUksv8eK5cezFo2TYx6dNfcNMLa8Qe7MvKLWNhjJ7+aDGWqloQSz1GJO
qYncLcnHeb4D7FP6D1Y99ciacOaC+PX+Tb668ljs/3os93WL/gZiF57a3yvn8jVlRskyi5app3AP
Bf+AmeH7Kfn8gDQWFe7tSsKbYr+u7jX9aXsZEEzH9TfdYUT87XtYiR/uIxQHqHbEzzXwRZQjfxbk
UB9RTpxRLSoOdaEnz2OQQmkzrJyz8a3wq73suYwsgdMfvaGYNW2Eb+6SCMKKh6CkHy4nlG5lsRoF
VIcEfoYa/avSnexH1kqSmYc1gN6k8ygffgj66dozzwgurTsjFlaR3w8Hh3NEcdP9GLLBbyOmmLk3
1gAEJyPUgszoh0aFjR5WPW2MwwAS0xQ+mUynftRdQBbAJjp7K+aOdh2IfQN9hD8nClCG20AMpgFC
L6BGZKpHzTHSAG20GWdka1OIgZQnvZB7LXklEemlrh6geWyZeISQFSBCxDK1IksSlTQ+IK8FXwyc
GYBwPqX4cDNI8QDJ7FjIPe5wOs858PU5XRgYRsBKlvYIafNc1oqwvSQvfwhDsfoKoILwwZ0Aiu7W
LovWq8ej39c26y7y3MoSeZQBWhoRRYYuSCXVFPqnHp27cG0vTgbsi8/+THjMyvLydfnb3CCUxy79
4Kb6CUzy7McAib1UubyDCtZLsehq1pnhCuBXeyaM6q1ur1/ZtO1HESDMboBN+Su1QXWkfUwpKNo+
E9tVWfBM8u5/CTAhk4uf7zX3ZhA9nr+zUI1jKb8iC/eqb8Ruhlab+9q1/uqC1PADSVB4vvFmEwmx
Lu7Z6by97WI4WzAk33HMwiftf1VpZc3BqaK8fgGZU0YGBL2RplPggkkHHuUZmXIt0BBebVvpD9SK
XtyPSFOecDJ19qwdbIQcmF5EEYS6j0Mw1TiUq6OwMhPDlLYGsCREUaoeGj+mndPvYmWE2oapdx96
2wnec1CtBKg0LevpA91gsFm45NvR08w2uxZuGOxzysImOzsTH4Z8faRuf974elFELr1LYG2OTYie
B5n8lX727c51BH/SWd62x4pzUcUOrKHjdNPLiIMDtpvIvDmdBSP7pO0bIJ/t58LOb8u+kMZmAzKF
8eNVNz5NllLwyhbyEz2o0TIifXv0uv9CcSx8VIOV1fNSQOWsWztevt2Rw0EOEwspQEE3B6RnbO6E
coxC+6s54E69cmYxbdGA6QLyewZe6dlayDi29aIENxeWawaFvfVppfOregoxU67adLrOv1PJniBx
8u0cRRPoRWlwzadfK6+MrXW5uBPc/b6K+GQYavc8xL4qzoJtuFxHlbgSpxzBFIfHuiM9CGGAu4w+
ueXGnMZoK0ntaLBvdfSP3umLebzoeWR7AFDyCI1pszHJi/Eij3eVlaCqWUgfYI5QY5KPzo/9aT5s
rlpMsoUKAPlNyYU3YlOHlzr/uPKg9MboveApIVdh7Q0nVYhy7IyjUP7SRmFYQgUcc76sGp/6lSEW
tKG6emhLWlyme4k7OylBIMPeglIIsrdpC6c4omy5/bt7NTw9FbxQROpiuMyhwHlQHlH79GvJxlUz
fymcpXbc/HmfkCZmJ074BDu2S+czyEBDt2K5x7J8L4Est5cPx7x1axmZQjWbEyHqZM2C231E9tfc
x1OEludXKD4U4i9Rjcw+naqDKhjpnqUVQPA4BdqB82SIAkNuyBZlMmHs15a2YKPKiL3w1rQbzjXx
SqRezXghsOxVRBLKhBBSSaQM2mOmHKW4RAWggsO5ifoSDcFGdTAeDIlfPqpxppLwARw/frD0Zo4o
iNk+emezXNbMH/+xjoPQRkzUXJQo0CbcnrO5L93MmKUnLRwvIblvunCXCNu9A/v30YHiWw7qX2QI
YIPq3C8dKR31FWbQYVyiqVGamO4ktvfPclcz7b5U3icGhYt3HBFLR+JtVrTba3afkGRMiKqwXIhN
72L7ov/2L/UuAnI5pUdNWTNAoufyW6+9ofbeuS01DgFHhLLJQ+AsxfDCtV68R/aFkyafTo7WhF0K
MHP2kWYnwO7+bXYo8MFNJIcHeU+/f5GT7EBovQsEBqHzgZb2lACvf9R/avrsqfP9y6GqLKyBgYwC
Sl/gnc7tC9MrX7ZIefrVf0tXP7rJ0p9vMk8jpAR34X1nJ0hLZJy9rxywX35boFXmE1+jzB075BHV
sfOeE7WFeqNtwVfWAKtarOc2P0cP01bnDs1T9VfSNJzvNE/UHIUPDLIoi4aeHCI/kIu58Zpfkgrg
3uxb85P9PzYXsFMXH4IIiMy0JAvXpaE4q+sAvOejAH1gjWVLrQVwoQwVJD4gnfvMylOKWLKkUCfT
2MwoH34x97h2mT3EQJA+P3HvbUkAuDlapFChlTWoxRuBe3g4aq/PLKjfCGP1HRgKWRexDNTcCZkB
Z1N074gFAuMSz6R6MC+cId+sA4p2GogZayL/jhD4JaguSA2tVoAE6pbHyH35eb+xjCX3/CKXnupm
Akt7GZktUKG2SDTdM+DdKpEo8qnM+vv/4ljFvwzQ54fidc2mGISjEgd7gPMUhlbE5mk3w+2F6x6J
8M1esiuYNoJeBTgTzmUmMY/2bRqCsfRQc67cWLI+kkc9m/E9XzQZCBjVOkUAXwTDcdSxxqq7rULg
vmhuaNczVzVR6TUFb80mG9mYtZh0X+Lk1GgSsxwiMrJIdOmF7sIe29afWYxL3cHf+qCtf4KFzNN1
rUbBl1Tk4CfeWIrTw5DHFnRfwTd5g+lZidjdQTwr9JOl+jpVERfksrFvS1XfqIFfbhdgIjNc8wGL
oJX5JY0x35Axrkkce3RAeo/gCRRrNgwSlycq7HSGaF2sMdWwkAVGfSBiehVCu6yoOw9C9mvapAWI
iv0UGeIlJ+AW1JXWCP03yC64256Jd79Zyr//K2F2b7ih5RRFIXcUxVLZSwffFu+m3BKC49j+CVPq
enJN2SovolVX6zhQDng/U/KXmrtkYzq9kPjbdR6pmhMCld72fV/DG7m+XSNz5PcSlUUMHZzR0Iuw
YUb9QMn3yzxMOK00W0PyzlwK8X9YlS/D/CDtfshVQWGllYtTNCX83TzMCYvcz7YKMn0mgd6jjJP9
FJBplKWIFPhTW0LIm7JOx4pw7epdEy1x0OwfNi49786rHOOrD15VTUX5fw66sc2266dBbrpri/AF
6dKuNtfMDQTGXzAC9EmwNIuibdQN50VsQUK8Y5+ylSaeemsl4Lz+weHb2sQ4oLEoYMoWuBipkWXr
TiSrA9Wrvz/P8biPiE+GDD674o4EXA5ElyW4TqGTnBNh2NfslSK7Blf1T2nHP3xkeDDRE3qeT6Lo
yAuv4RZMNnyo5XnhBzyo9uzO3kvTUNoaiNHq3JisQ/+gqtDHEhhs/bD4kyHF88XK8qKq6sc2MXsu
tOyAvHnJNqxhJP7C1Kf1DBkEsLjzaPijC5YjtxxOALvrc84UdMJT/Xh6xLh32cn9LCJvzUeCDQmy
6Oc8XUbzq0lNRvLZ+EAsn1TCjAFybBvRvMBh7ofU2aTb83GPE4H+8AYTQLITuPAKjURaESAsZiWc
S4taafWHcFrS97cqt5GzorJmu3Ba1F4a9EXXH8P8qVblBryc+NKdQvjoR4pspWdntMV6HJfxPTDd
kOmRTB26U358/sUmQDIponvHE7y/ZyNZ4qEyrPdsqTU0ZOi2YaVmgj5VzLu3lNhDiWppsspQWPaF
ImTwbqI0+wkJMCDzr0OrbZX2DeGku3Rjsx0VjZKwF9HlkdAJiogXwNEKYw55J9dF8uJZqtJBIMVq
corPpW9jcxF3b2H+Ydpr7rFFi1EXxrvyLBLcC7hq00jlXHB9WAD+xT0qE+oPNkEtsGMY7o6DTW6R
CpV1QOymD23xBBIZvyXvMDmOQAPXTJxMJ+WmNb6SkfkZisWe5770CpMg17pesC+de4n7j7oYgkEd
yxm8+I0smPg0Ok8sK625V1dP9VHy5zM1VoOepvx/PxAjbfj60U6HxaifJbQ0spz5DNHsbLDihk/c
EYK/gRJr3AXPmXG2pR0qfVNC9QmWUX2o7XmWY2VCBevJ5sZ4PnqnQb4PHkRYk+YNIhS8OKvgijNp
fvm8KI8+zlAWv6ACDK2GXoa7maP+fqK0Woi2OQRYim7k4CBdXizeTyTONEJS7v98+eQV7GfxBDVs
YKuNhb+Q99tcp+0me5cQRvwlxrwxFlzc4kDVl89SBvkzOIcLJH0IJX+kidqDirGLqpKgU73odJS6
RCeBcwY35Bxi0yAo7bDYSYo+C6bLi5S8agE4uZI+Wclwh22lzHaau/YJG5NFrECQ7gE7XbNmf0P0
Tmirltjgojt9GY8/TdLalnYTk63cjk0N9jQ5Fs1jOdAOI9B2hu46ozBRTGEGA0/fbBK/OVZF10Z5
hVT1JuV/9aQiNTlRYgkG9rx4jPHkaIsfHPU2gK4Z+7diZizntIfLjdBOoFCiOkS7jA0GSlKRflIj
PmrKzm7i6XN23nrubGc22ivgxqFoYrxUWEKJyKllVN2vCC9ZhRzIDtvkwJ7hvH9DQNPzts/1i6FI
ixAK3C/sW3CGIPMUjldvtURA13jt9OvGWf1IA8Qs1z5i/aO/6WTmWtLJMrwgD8pwfJpNyEgDpGyx
Q0rXZyGLXfUIqUCTW2EHQMPU3aPVSWnKMThSgdpOeAOVg42VH1ye5MOOPjSs2VXX5oijUPrWRG9c
R6yWCjlT2POQJwnnu0U4eC8YwfVauVDoFNj1Eze4GmY94VCl+ZLgCbE/cz7xOwFsRQnEnqAc6qgP
iFLrazdXfx98qdBAjvJuAZkQYNLAH5vkrMrYDTVFvy0cP91nBADdw11hnjn/zMi6nYT+3Y+RstyF
0PgO9q+VcQJpgwF1Sts4pQRiS3hoyZvBKzHPsW4SLwMSRlOLvcNlB48LEGNaDov52XQ9VkSR9SaL
f2dSyfDTj3Ee1vpq1VuamsZmtP5L1YK/cdmHReQC5vCharOOl8I32GNpoYv3NuZTOJqEPMg1VTPQ
dKrnfZZOPv6ClxnjDy0mXV3CCZRT1t/lzJOotCqspG/M1WsAQy8oHz4NXGk286jdCh/aNNdRPKcH
z6ruaoytBSPHhMQIiyVY/o/mqT4Y5IIjprfFCMO/6zaFyP6PO66Bmihbd3kabgniGNjfQtgDJx/e
MTd0BkbWaob5bc97WfYudRwgBYlCKhWthvkNbtg+YcIzMmZm3+f+H2jYF/D/pew5IN4QiEd1P5to
ebrUkqOy81kXiwfDWvdRbog4wbhDEUf+4ivJ7ELr/nu2D6AC4PgMUWAfmNltycBS0K4TLpN51arx
rB51DiNSJf71m5WTnZJHRfLxVnuV6rhpkoLTvM9d3O4dI11PhhFkF1r4thjOho5D3M6gULfK8mhy
9jj0LX/J6pxAX2/KFvuaU1FMwBMPLpZov+sAhn8UxzgndyQvRAuS4a9Ft6fa0k0CkLrmyUEeMvzi
CWwkmtc4NVwlPHt4xRXTPl1MDHE1x6bMyZ/Towxe6oudn1j0MCjuGVmqh3aI2pOi5foIsR0DzV1N
rCCatnHPfVH/MQV9g/hXx2kXuWKHVQPbDbGxBDaT8zaE94gNjeixcPnKzI8jS3CqzfLQd8ykqMM5
ogkiFV0ugWGo4oq8TM3kpbvuE8OKwdWuwxzcqPoG5pX1vIZVqZqViQShWu6UwcNui0+Rm+dLBi4J
0pINj2Fwdl/OkbmHSQJZ+AOHOd9pCLMS0VM+fE5L9fMo6TDfGePRtb05JVSKOKUJiy5TJjtW3JMI
Cr1o+B6eH/IpVNvKlF5bD+89HlGGkQBl41iWivlDb4rezEZxasl4+4bQWQe3lUsEkHMszZiRBXYO
QHXU9dPjOfXV0Lcng3HU4cLtHN2oGcWfsljAgEbhzDUlrWqv8sY3NH7Ajnip84ASaqsCL7W5JhRM
gyDAJeOE9iyyBrhkNT6XylUmiQ51AELbBFp1vMPsLD9LmA1Aea2O0veTRFImWSfZMcvWUervSyT5
WRHdBPIGWSumcC3wUedjEdCe0mvkWr89NBYKEYehgtkTIjyTmb6uQnPoSWBlwtHTMUR1KrQPfwYp
TmZcSe6BxvlC/JIGLEDocCqZwBxMw3wIbhZsA2g3Z9K1dZZc1+N3Wb+Ic09nzLGH7AWhyL9BIBI1
QQD/22U+V62oq/kSOC7/jmqMqWsxbP2rFXfaTiPngu2qoMqB0bsqwLY3G11VQSnfjkwqoxQz8YiZ
VtFhZMO9DMb2Tq/2jUWu9fUtyyw1/tIjS0N1XjwVFXpHBHHDVjndSMvOLBBeFiX9tmkDVPZP+P8s
n93ChTcq5rYEDsWIWR1HOJdgSBdnsaDov9T/5Wgl814ziux2AGRcOuAkYr+Uc3uBunIIVirB6b6j
GKCc0mhN1ybmwjAJfPKwh4e5rBFuruNCzHK5IvJ5WWsBb5Gr+XZPh5+POWolpJtmbqbRDaqp68E+
2wfVuEeKhyUKs03nrRybr7t7WXq/jQawhK0Qpr/LzmjpCXxwPiAVZRxpb25Ph1VzdNIkrz6u8she
rg0PhF0JttPOolvm3lPKY5655iqizfDhVmNAXpShoioVmKFStb11EuHwdXepeDiIzKn8/WzA8ASK
PtUyOZTG57MA6MkWNzuEicxgAXOskBWNq2bg4QTHKHN7eAiWUWgfnF4LJW5JzY2zw6zHWL+xVRGH
YnSmYXE0OAYEhyEH5cJb3h042va4K48d+QTy1X0zhR+jWG0NbI7r5l6aaBTrGowku9b1kaq1Gcjq
JTPKr5pTjk1gN/AfjpV2iurIVfKifmKlgBCDCdNLDzmBP4eK8COFieXyGJIvJBEVu4/YzV/BwYSJ
IhTtsCQhJUlLGL/q3dLN35gqk7ESwsIO5Lrk2M7zV5LleSj/r2SbNzdHK1lmoRi8E8Y8j4tOFySO
7fGACuTxHqM8Dmd39AXmt2Y8zROkQgmwEHm0l5KEuJVzYrgFFA9W/Bp0g68Ehe3mXSp8wLReovP8
vOP5n/ed9NcB2qzv0aYQf/jSQrS6jEKdD/pB6dFVsaYCb7hPqLzlVGtnJFGnTzwqsVAfwHu109xp
onLro5S0rREjijZqkd0Pg5xx9gAhrJsqwK2ZRfPMdIi2rMf5OYSttNewf9pYnVZM8N+yk44wi3cc
LLZSfBq6XTgJFCDrUlIM7HYXDwUJ9ApA/kzr4OY4NcZcGYL5r3HK2Qz6hx/VJrOKYZvbVUDQBI5F
O3u45u/Ma0Iyr1oehSQfY7Si+lieNK8p1Su86UKTFmAdEeQbLcdsMevEzuh7p4dBd0b6LHLTkxNU
8wQCWZ0AmkPj2uIZrJDWawBghHN0l+Vhpo6Gs+y2gYQwlHcOjEMpclienOs7yBLhslrtcJW1Us7e
X/OScXOVu07atkBUsNI/v5oplAs6lAsqLpoMiNHI29tcRAGZYtg1bqr89Oulw/jDAWiEinyBno2z
MOunq+Eq96vH2CD941ehhrpMNro8E8k9PVM//VehSQPxeU2aBhknfwT8BCu/ShRx8G4kUmI4qbGD
2Lzo6IN2uQPokkNmLDQZclxzEYWVtiZCvcGuabVMj5O2KXmbY3ajt9VsCwa9++9X2jVbhE7Thtcg
d6Qka5zpJ/bJfvsDJOK/XO0enFE0kcDWiWpppvMvS97pmKipBO3qFSrZ4up97ngK3aBQS/Zl3zqX
3vKrDFbopFeCnfy5cVuZeN6Rwc/IWMCA/lKe+ryQ3qOAh8ugp8JJC1zLkVoRFDAaJIqSBDPAu0yw
eAaU4mQANrg8A/qkQdgDa/ei7AxEgMYWovD6DjAmvdnvHq4LGjpYcu58uGkIAqYG6rvflfjwet1i
A5iA+TPFOy3nxAN+v+gDLVaM6CBJljcZop0+7ANvb1rtpR7sW3y+2foKFozkF41lWEMJGFXI+Aa9
iBIMMaS+sTmeISOV12JsWs0rR0rIMqrNagMsGhBZlDOpjb71dB+5Z573BfEkmC+o1ANUzU9vdBVS
5Xg31lzxXaYg3PjvKj3pZlBPD3j/xif8jHPVEi5qsje9R2tqZme24yyUxUeckgtlnD9EICytW+w4
u2tu97S3aidRRMT2D3TcklQXQ6kT6DT9gvRCgRD93ja1hnHfW2aSIPXHHrOb9jn7+805Uz0PUDJG
iPfo3p1+2ECNyGHB8cR9Na0dfRp5+5H4yMP94azl6vVPf9M+khUsW+zZikPQsEdJwOQ1vXMLgAcC
BtMexEnwZfbB5WLhdM/rtmxYbqrOthkXRWxHNb6zKAPK0M757KlMBu5KdkhCBT3v0hlXFbSMqKD1
ufh0ivyreaBVoUKRS4QxNPXqb8FWPe7EzbsjQd2EIXKVqdbTloKynWjsM+avZd/YIvyMrlVkyAts
1dQiALHKGIVi9FIa8Yjy4aNOUF6Eg1BkLsQNqV6VLyyu+RYdYvQoAb9uXE97nPVokVsEP8DAew7G
GTbUtYHIAg1/ACkWURBqh/RcdQcb6/gg8a+0HVF0qr8IBfd/8LCBVhScz416yTMuJKpeVJvcBBMH
GVssjnZEnUVt8yKdiBnQTBQrsD6EKpbdazc2Ba/xQH6DcSdUsB22ngkH9h+x8w3fvcnrP7/Cnv6z
Ce2TmJamYn9+Ri460qE5JQ0hp/kKKQ0Sc3OrREEUq7rzeojIxeEg1+EYEvDExUEKaIUBPJm3lEHF
YcbFU2A79NYXi6G/iYX2kGu/WBZRkfLZpc13N/M9YMtgcYI7QVyrkQBVWsF/DSU1MhdPHbv4gAir
JALLrKTfsSqbtcomGvu9d1+/0ZKkgWdhLHk8y0ULl10uepzL4nqbVq8+ys1GrBga5VskJAclI/Zk
p3BeMfIneQcXdp0QAzz796yyUhBz0O4lFudWgnTgFXItgX/sE6YgrrLgzvKWsAKkMLqEAhXrm617
2oilkWdl9g9BUBUUfK0DcA+4/XFVv/uFtrIp+yy12lxIDYB7flM0ABzUp9orDNPis2yyLKNuMp8n
4WDYrhhDDtSAx5xVad+D9hg8SjfCDreJxzuytCHvYgacxJtxHkVg6b/m3/Anb05WzQ9c93VH4jzY
TJTgkZ+gG3o71cEmhvaS12CfrxVYtN6dLTXPAhxeM1bjBQBjpm0w5JZDYTTqSiXynYKsF7dpy/5e
zz5oTABAnNTLcV3URhbnHw6ayxT1tNKawbe3ZkODPMVQ6FAsrRnCeL1S7lcs2TjhN8TZ0skcuBUM
VSAfs9UI9ri60XiFcqR9yfsfHj/LybCmVYJ72E199E/dNZgSp4S2pRZnIS4SgpBFMij6Z7ghZ7C6
VtLrf8LfzOBQ/MjTsIpwiGQ4bqi8xq6SAHjaal3ePlqon1NWgznECSzTHIcdDcsRvRrFUPFajKbe
WJtktL7NGItrLcoMWdpYy2v9ttnhRtr77FXOKXWvWr04TRqX1/i46RjmbAUbzVNw7FhnBtXhBzJn
qt+FVctrujidjfbHuQ4jVvtoCa/GtvD/wAek+krrJheAMh7Si1wI5tfmGifHLi9TiYZBAmNVxaWf
SjpUd8Z7Gav7N1CWnl0WIChFONJujW18Cy1zTsRe+XR5YPNWUtrW3d7QFW8RiLqXWcQnVk/TCsdt
KS4CxKNXV9O/+yxGoMkGPoAxTGFS741w6hg2/qOPkhiNwFP+XZ1R+7OZRr30PCExangYUGx7kaou
amrTI7IWtPVffrqtEulTOnkECU9Rrz6pphxET8fCAptZYmKQzoUwCYQ7af17iY5ysANA2oyMhi3a
Xqma9EtURZkBF1qibGazCshm/6dlp0sA97FNHfEaO9nE2KD5VPZGcPBf8woHniQAcX31OEc+vfFF
W0ZeIOiDCrViDDTl1UV5MD6EBmj3/pAYQHiQU0zK+qO2psV9IUj91FFoBjgM6f3mg7h6ZW6gu4SO
XpnoL2Yvd+mrS8z01P/WswQ6E40s1CYTfHPA/j4upQBBmeueTXAOwNb598K5LwlUpPLYaSLG9tcW
L4z9PHoYsjMpXY7YpDiy7E9vnh0lofvGxYZ72EIqZNeBMvRLkUHc70YEZclhkDTCHuL+IUNLsxUc
MDBhPRf3EvM7fX79iC6Uy5bxURVVHNxMn8uePXvOgRNXFpQd2QLsywD2I2QjUlUdalgkN2XLsDyh
edUGvesKDxk06PTvrxFQxtmCeW9qAzHQliIieaKQqIXYmqWb2BBKKtB8P8UiQR8Js4pgwUvgkCi1
UV1QATlIxComNz3C8tp6uUbgN33j/7lDN7K0iU5m1yEZ6WDsEZAAz4FR6T56ShHcGCysRHgc7VZn
B53lVQiYdTlGonETBurhmzgARkuX90UK9BxbNHyuqzUgkn1sfC2krEtfqJs3GF8GmHLGilt8fcLh
5DQSFPe4UH/gt6ajxMRpR2nnMTfJDePZOkWLX0cqNd7WasWJ+BWRYXDeph4lZLs+z/Y1VJKNaITX
9qHrTkBFCPfAz3pwp0b1PV/QE1RMac31u5wun2GKreYb7X7nu/PaN+KFw0HpWhlVLd2Rg0RC8lGr
WePgOj0b5sD4K01IQ9lP75sD+6z4/zYdNZb4BYNwj9eNqjZUP+Y5YuYegRI9GxMNMhcVGp8XMy41
3YMiMM1AeJO8BpsSEKvxV+Okk3vAk3sXZDs537X9F8y95NRLgZKPxorheiTtUxoOHs3NcoTXvdTv
u4Z1w0lHC9isv4rwt3xr83IsV90J+H92ZkFzxCXzpMNSoq2QC9snTFxREXVId4Mfcg6FIKprVJU6
8zWBMvlyPzYMsjdBmigVF7OO+yZ6TQqSdv+AN0AvgiA0AcTdFyaq33+fcASmy192wrmVLjDFt194
xKS7llGVQEH8OqxXqU75DdxX+VH/RSWkM6JwLVYh/7p6EGL83zQX0acAgL5NZKLKQoW8NlwL8Xfr
+qoZbV34U39UaPE2WhhTqoy4BrvdTA0nxCxZcjplhCr5+HDCmudjcFX9dD4fHW6XpHrolW52/Bu9
RdGE85pVn0z+pNxecQO4NVt0KCA+w5utHZuadD5NkZ5YHzTrlwjJ4O7cbYIEx2E9HYXBo7mKSGsH
7Rx/iEmwjzUSTba5WBMrDXw3xf+XlUOWtR5MFQyQTPGuGSEcXKmxknW9DiRp2szkfkJJELJy1ZpA
cZoic3ws9ohDoa19raeRjpIkchK3UiPpB4QVSQ5b69vjV/hzB9Bk2d5RXP8P7HEvVGA85I0mh4lG
mviuP1O/4LxuxU6brhz8GInVCmVJ03XWuOZRWFjR299atLiZLNcnFiwLiEsMVWbt9U7PJapxI1nz
/ys/GDVld6xavqoK2Iuc2jCHNq7kJRMgqPp59o9zRfPdW2OWcM7bSooP7RrvaNlnQcNg+8Pztjbm
8lcvA+Xbu24T8lRrYhI0zEGQX+oWtRvUH3FKcqNsaNWBQvUkPz3IjeiEgbJOyYCBq/Hbu/cO9ZHp
qEQaMBqxo93qvd2MaAtG0GQJvu4xzaytmaZlLH1MR5/er9hZrpuyS4V11Qhp7SpFnh9SOnGhBLT4
zLoD6SRD5+PWlvUqp1Dlji1SkPOBBFuZ+zv8uaWVfGMvO7zB0zPVeRhoPRRwdJXpXpumrfH8h/oL
6S6GUuhdRlz3qb7KH78AhhrHwu0FPP6CegqAffdji4DVgnhljdWqVjhkmbOGPrI28TMAtcXHK1t1
o4VxJdiAol1VGMIDoktntsGM74nP92V06fASmzGyJ6zq5RUggQGq7+OuHwoiiSVIJKXeDQh4QvL9
5d56ZIpaSyFNsZGWkRZs6GWlRWnmgZ1zUmzDnNqfHOUNJDUDA1EX5k8/BuAeTewWWWECnqbEiKuC
j0nan6gwLbF72h3mxv6EZ4KlO+7ppgga1AJhtLBYDazZEdDbwg03jbtB9jKsC7uBDcQ/t2t/tksp
8c8B0JIy8A3dOxXxw40RRkrJbCZO2dfTpBevBeq6bgZM44vVDc1zlPU7W1dNimKlCOHBmCyPiCu1
0EppCVXoktjbSqV9QutuecXsSUxUts0bmHJ//IuBVdkQ6llXumK5uCcW66MjuMs9z1e5tA1NIRyM
ej8H1LM3T8cxA94XHyEniXwQlVpCWK13trGLTMO/O8j0Tm/FR3JzucThJRBDxmJO5Adak/Oi8EMX
SAqUJKtT/SLk57IS/PWFblDf4ViZX7S60Kg98iaaetGfVlsWJq7KQ6wEUrCEgGtOkw4rl0iFySy5
sFubaUzH09F0mKDFkgoSHh9NW8bVXlgN6L5pmmOA2xUO7T1fXxlUjQWdNoeCzmqAFeS6XCHXi2wG
79ruwTGYU+0DRf5x/wXdXXqie2YaVZkcQCbtDJqwShQCpbeyYhnrBe5cwSGGQWRpFX+V5r9aI6yR
WQ3WYhVj/9seqVFwVCTPX8GPLdKbTazSOkYHTLhxeRZRw8AxhDl1NR4j6o9scH3l8lvjAWyL8hl+
dmWoumxvi3GoFPgylA7BucD+nq2z81Qop+QiJhnwZo5kvz7623HbaZuhUsI1tKydv2zj//LLdfHU
VxF+CX4PR6hEWfBhcZR8wV+7gUdZ3I3peawcLmCHso5BWuHyB5QTIqLYZ3E7Bl96YZtBUqQIVL9z
WEh4JG4obotvPBNKgP9bg6rmlRo5YnoUMIiIbFPqT/ygUMTbpUQGlubDF8wtyzqVk9OCxq8EhiUT
WTUVQTIr9AaB73qQF+8Vw8GhLfsSa1MtWix4g2fxm8kzEZ+1mL9t33d3n3wMkiQgqhmxyYtfEMzm
4sXmQeFOS1j5zOn+3Amasp41YUwpSwWjjYjMm/Jq2PUbQZIioXmxH7vMzOt1esblMPTs2txh5k91
+pJf2E6bSIDNBQj0eiai+amYddZYj4Sav8EtkzyT8ted1vsOuyoqzsgvM9SCT6m9dQoD/QZEhGo8
3ApJYHLpFH6mNmw49zvxXxLSxZI7AtMgKrzi4vKiw5zz+sflXKt+WlD3I+vfosOmtG5o2GIqQ+kE
IixmgOM2lFHD2gF+P2eHsNx1B5bzGRy+n7AsSePBmZdf6kp3/79dscpDgQv1EU4+erRyISV4etnL
k7BmXUPhrMtTlBmAPx3ApneYnoLFa4AgOv/DgNfywZG2NLzCB70CzeB5RF45VCvk9zms14AY5AoV
OxO32n8DXScMJAbsU/hgSUDv6EhCnpNRC73aT9ZJGbwQ1FN6UZtokYpYly8QQch6R9IQ3Ec6nuNa
4/hEwxxv1voFgbf+7yfINX+h1PcjE2C9CM8JvAzYt55T9PzYAXHwAJ7kZtoUGtQeOuSBAyTKZ6/k
/npR18MNe0pc3kNkYTlnl0wC3PzPwuLi77Hccjblf9eB4fRE6rAGR2B4McuegIbyuB3Y2wqUiN0s
0IviivfvKmGnmwOxwQqxPIKkTqsYvK6dATWKMpQYg1AAw79FC1+tpcvAAJAcVsmJPcXw4i36Qu42
atMh9K8XlxdpqURZhDULMIB4x1DcgXpwAUugoiPrL7D3I+Ul1GjUv38ygzXF+ac6pg13ig68Z5rE
10XAmvSSOFNKApfXZBZ3A5VJLS8gIy4Bjgqur8S6Tn4HooNcJnvowX6pV8ZvUm8jdn4GhoESl9fJ
YsK1ps+mkMunoJ8XsIPx80PlWgrTVnmEEFZGFbnt/J1U6+AWyltJMt4mfLte7cl91bGSPEcy5Jow
JkKKX9+G9aexMXy0i+0g5yJpqa+bLgK/ahm97wAJp0/ADbmTpEeCziKA2iBWCIMKJFtE4j4XUgY+
6SlE/XXD3SQcAjUYubPL45cxofOKdLCcmgUfX70EKEvt7HgbcisNjirGDpuq8D6BVeNBwwBEWZrU
Hu4tPlJwVRzvuTtDcy5DN94rDGhdBHfn1ccHmhBEe8Es/6HB0GUlE3MwUMvn0S6zm4vGn5CrC9mw
slNFOgq0k/KJuu8lS6MlSTkphqEe43W2cfksRLo4R9UIJR9MKe5treBaXdbJu29m2UMbjGgSogo8
XJAhJ/z82mCWuWvYVbmWWDFrrCJrvh4vk0e8/OMq7JwLrlML0ZzaQnNtkV29VgWffIp4U3mtTpoX
0lzJc0/9/y/PG72YwcWOxx5NWubXwpT3hRKxuIhmZOipvLvWc79b3+Q2JoTN9opmlqFkUguOT4CA
28inXilB7yc6BMuhgHzz2l+79v/LMyz8bSPxSVOcxNzPhEF/jEWNZGQMxvWOdn+p+j8T32HkRZdc
H0lfcgwnHYM2w6vmMKKTzp/NMQ1Cslde/6/z9/BbO3fA9Mk6m61+oFGoOcxPs07NtglI3QC+1LPL
iX/8jg7kfAJLx3uGTpB695wLU9yWZE5iwGLnjDTnNNQodmy9yzCbKchsju0TxnlZ6iVRfOfp0edP
TMqBQEiNyy60gDHcI4+pQXFFK+KELa200nIZCzefWA9UzPKXryFbMUiiBROaa7QDnYrCCto7+oPE
VtSYcm86o9iu4gm5GISQ4HkrZRQIXUGh7epjQ2PabSwPMyE8OWT442lGMHvPVmfimCIpKeCrWn+p
uHyRqFkv5NzVPql17E67CnnCNGOBSEnZkv2Hhj2JCDtUQ7ItJKFjWhQH5EzBRHDW+Hi8p3XeljLP
aiDDn5KN+13z/pfsPoXVRucTxw/bWCEA5GS0I+iAwjzO0w3wDRrpgUOPAdUEDsp3iDkHynP+/eMP
kTZ0MqMsi5BfTjPcmYdtHIkX0a9XN/U/66Hqfqz92B/rp8bP9cVyrX/dRJWP/CPCvo52M170fJhD
jIi4pZkDcOVLeZl2gK/mlo31t0dwKb/bvlSJ6SNjQX9wtTQDMBPUpcd5BBFijlWV9BU9bKrbLKwT
YQEHg6QumjLKovBvR4fPqxIoUUG3YuXP/j54R36uel16vHutNvHIQ2Wt2KOkDyoU7cqvF3OTeJAS
IiY13d2qxIfDHSXOVAp9dzvs/NFAm1cuka3qHceEl2RugFku4/tl7Sn3rVZE9cPybm/bXoFfmiaN
ySbrH5kAapAoTb00cpJkgERhZ1VLNuBvqMzvTp2wnRbq5YwUWAQy8BksbGSmE1jsMmwatEgGZ3Y4
6+FxqFLIWNUqzUX49m9J9d948i3CcTGHe+PSK46q1oSWBq9T3JzYzhuLvpsOsPs/rO5KgaxNmfb5
8r+eEQgmdD1Wnk61mhfjck7/Luz491sCp41sJhQEXe8jQq7FG0RuCS2GbyMdmHoMUXOL4rfdhHDJ
I3G8pwbcyoOiCdXWPj38icwnec1s5Jk7gKqHRrvNEAvhuYR1Okrh34gmwjlKp+xnCWqCVbRemNAD
h1hfzBFu2jypqcweLqjB1f0g75/03gu8XqaEIUBNo9baWsbPUXYGZ4fhk2+hXJ4EJynaSpaP54yh
kRdWX+v0y53KR4NtGmdAShX6lVh01MrBUy+m0gzAenjZYKIcJ88hB1QYmS7oH8+vVuQysClv/tXy
k4t1UCbXhm1fbxOAEp3W6xzFrTKC5Rn3Im2LKteIwPFmrWtkxo4/yuktmY+eAu6e6YUGf/pq9ok2
PWUtLHOLwfge+nAeTmq4KXAeKVib23mNkhLwmsp5gLNb2fNKkYH1HkaJHwE9fHeQeyFgu8iV+sG0
gIIRe1J2aWvi6qE3Em7qlrbpnd/bnhQI1jvQjv5VcpcjAZu9Yd4NMWuGa8mC4tEKiNozGRttS4a0
kK1PMnTGYf7t3bG0DhUzAgKFznh+UDEbXF4em8RgP+HHfQwQ6/en8y48T7mo7EA/MsYu6QLG9nXu
hug0eVXoEl82PC42p06hKsu+huHI/PXt+jMDuVMLePOyRmfkCqGHwDIxJNLh00FJq/9kK+Kf4d+s
mCcFCHPscGbFZMx0YAsN1UagEWmrL87UX8H6lO8+U8c98jWR7WotYVtkb1tkxogZodXVIdQ4FMTH
i16U5LR1B4XRe41dOp7orwARkah0O+FXLay/dwHnQv6+Eru2bL5bwf54RQYe93NjVQzYHKasHg5J
S3QaiLprqVXZ6TdGO5G36UqwVFCM/jH6nP1OlUrYEFK+Rp2mRh99ChJ7iSmHq5nbz/KZqihnXCQI
pyMcGlMxc906mJ1k6x3plcwUOhuPeG+tTSbrLBzn3hdKLoi8ncqyyyM9zl7vQ8p83TPuKRAWTMsj
5lrpJKHMSP7NaJuL2Ho7HQTfAKI94BwK7XlVOk6/gEQJWDFO67UXcTWzxm+jNoPfJQC5V6gD0JgL
/pUZesaZzKFiKk0SLh1cQeWtpp7aVtzgl7TPjCfHT4eOB7EHg9yi9BUmwKZ0IYIgggHDvBjqql6t
1XhaTBEgEKW/r/5g8jYaXGEC3iiGVJ17EACuYF4PrKFs5m+9RPGYQOPnbK4BHOZxVcOcPX/BBx+F
wm+cz23LstMiSv9NLvj+kwVHfDGNW6t937beBfSr/HPCVCySvLzSazEBKDzIC/kIajfbQCTkma3e
5AwcTbocT6DgzDDYyC7bDwtKd4QnKM3fFKAjIVh2moWl5eTd0BCYp1vqXnxG63cOScYwemfssoFB
agsj7bfzYFfPxDabUOHAwPsKxfkH663wm/6b2s2PnZHAwOM+q377Ghsy9SyVvvxXXw6xCzvbS4J7
UEMudI0eaxyqtAaAxug5Fi/5hiOwftoFcM6flu10LpWJ5SN1yJZLez+rV2iq75HFKR4wAthhcUQ+
15GUQUM6zuF0HZ2lxTePIDs431Hz9W12VUOaihByaWG+yuTnQqi8w+stz3sz4br2q55r7buePLbV
isI6o4EpN0i7uuIbBcKG/IpUBcf6nGzECz9R24GRvNx0dqmtHHKx20fcRShUCxj2mG7PZOFeShmJ
bvnykoDynWfQrxAei+QdvAoqBKl93VG+2mQtYadJJuCnONoADT/PlT7WP1+hV6TweC3U8a8aJH89
ISuZihgPSds97hBVGZ4fMD1AYUbCqDXqSda1yXbFaB6DLo3ye0vLXzKs9Sr0Gv7JAf8Z1c10FDHn
pw5N0RKwbZMGCV8sCpuTuPiuGUfDQzWgETuHMliI1Vmp8eFowd+4N6sjTDEt8RAKStm5x2YpTW5/
zthJ6hF6kV3adda0prB+gn3/7U0h3gdX8ItHw6yJeygg4oHUH9mLGhZMA6gw1vwqixUk1nBqEz+M
AlOiOaqNVcsGvG1fQZydDac64HSCsR6zbZcICtrzJCmvoLW/b1SCAZSfwMJVbTNGNtefYuafgL8V
aEVvVkxCfpOpLhbJalwq/VtAuTqTKj249telQAr2rdKRAQ6TR9uYuRhijt/6Z2zoCXNvNLgG49wH
tocfmHnfKX0ft80nPCOxkeyPzAmvQve1sFGZHW/9EYPcHgByRlV8wNGGpqfp1eh3EA2kPFSLh6eo
c3bUxU2+wCLQaWGEdYTtA6e78EB9ikRv0dYidEfeYtG2SeEzaClwvvXywu04uur3cM6+uVlnXkqN
M3YGAezbV9gfcBP941LPPB4eT6iggTzd7mTX/fvvK5mb3U/Ihgp8iT5GAh5ffF3ynRLNzOhVsHYp
xvAx7PfPtcl2BmDr1k4W4dM9u6d+REJhCy7lpqRm3xhS1CCNKxWtSGY1Qxe50e4GmM4SUA2OAtAo
w7ZtnSrgAG7ff3KhoVOGFSWvez3iZuy5rPU/0E3I5yOr4YhGZ6wvYXj83RqpQrfnwEPeohaCIXsw
9CvtMo+bWd8G4hu06MUWYEuNS6d92mx5ihwP/659ix+e9v9dyoCwvumOXg27ic7q9ncYpiC5NOvW
mW0C65RJp3WOdVVuY75yN8nylgbodxMTb+wA7XyTwNZ3JSgrb0UCsAl8pWnCCDIgzB+Wckyv4lPV
lJXXBmeilOgYIxXBSIIpQTw7Pu0obaScR0YpHoq8B6f9b7Joro3e/p76SNAm9EkFzuHebtKB8yTe
kiLUrnK51cQDk4IB8fCdftekGKlEOxcPIgdT+VJnx2MkfjRovRhm6svTyQYmpdFraDlgGm8zgnSy
oL1bigEp5lnKPIuDZo3xDBW2SbUWdf7c3utxEtAXzDeazquMJKdD4JcPkASPVBjy5DNz8fw3tbII
HSz0xWxpRd5ElaLsVaTS7aTNYx8dYI9LE827UUv4G+nuwttGmv98WdpcnG3lGonjixsQSmS50ZP7
45DH1F0mxwmeBv0i7Lz62A3RXO3MLBAADodfL2tdP7/DY4QKh/BxDS+MuzPthDq4c5FpYUuTxUPT
AFuupYddIN3fKlnr+Z2ULkYQOCjSN9G1+MykfFdHa5ZHsj9HsuKbDuwSVwdye8r6Xfnzys6i6gER
1yY93aeg2vwcyet0Qs/G2qnMD5imuBCpkx6pGdeeE9UvhMGZ8sUv3YmyD4iR/Bo4ody2Qdx7/geR
jl7a4/09xLH+wwqmZCIlg9F6Wldc/fz6Wf1Hz/gvikM85nX9ObVnGcoG5maIqXAGiW0GFuCwTdl2
yG71Ni3Mxggc3B2Cmv2Qg/+YPgj/Sw4eyaFmumPf11hMtQsDvHlJDC1WzFJQh7qQ0mE+xTs1vipe
0qNNQ5Jv1j2d6Im8hi8glba8n34kB1re9typDRL3/WtIJZINenunLyza+LuvGMCeT73LDk+UzvMB
z4BIveooe1dWimCPIHkbcwZ8g66Osyz205KfAracrhKoLFtfLK3SZB5KbwEVOKIAS4Gj9TR7dkjl
CRs0CchR+48XbQG3hRMXtiYvwxQ/utkN/6VJnPWitRK15VvUhYUevEM0XA8spsLeU031TVfWh1VI
2NXyYILE302VdxeqzgLSckOrqIaJR84mjnGwT5rNIduvEoAWgIup+7HAhzfZvUm8RvI1ApeUycqu
+kdguzEo1qiE4h/qEYQd2X35X+p1lAaxPHoQ/hNdPpl9YB5Igbl+a6mSM9X2b+AtNIbAf87GA23n
vc6gFvo63cUZ/bXms3VCbV8c8y3In+ARqVpS5MrEtxkgDKYbXlbWv2Vyq6CxuxsJ4TOtXu9WF9/B
GhyGHGRkIx15ud1qGXRhiCaKhgLzPJhIq0ns9yOY3NtiVyxAzFA88ZYsuGYPRK8QIqscut4RG3eG
5bPEa1AvcuwqOGLiEPohuqJqnmKF/SctqXjzeAltY1bmX335TICtyTkrW/sp7cUTWrn7I/7hiozB
NVk8zD3F4vNP4Z5+7XcJ04PlkB9XxFTmZf+pFMWm3fAyFMht6TTTJVGKXKgDgIMT58xQSXgqZGoC
PfLpVj6NEGfssfGx66yktdsyUzjJFJbNd1NYDDD/d83D5MlY6YmrK/wzERfhfMlPReGx1RMc2MyX
pHyWwynA4UOWEihkZRCnIlLnp8ahpJ7LSES6uV6zMi+v8PJ1fxugkKXBF4PjIWqXCkM5zBTgOQ6k
fuHOBG5TNBk/MiD1Wn8EBmu9aaUMFHvXY0JImdlFHUfEXLWOMhOed0xbiIhyJdfAA5mS5Fk4BW5k
yE03tZZB7GhByDEM4fo5Jp0tGDR+/gFH2tecGINCb1Z2UIZifrfOIujuaukMLgdIRR90oC3/qWac
tduQG1rVydtLSHNjY1DIBmGoY1kCdByfYF/jfv9v3IJOw+hGeZr83nv8qJTVzuqzkLutLzvwmA3C
8RwX8r65AW+/QhvVi4AMxl1XOhvD43Q9YEeTl+hRD31MdoJnycdiK0nluot7HCY/KXO/IHnQROZc
mphzijVvVc0prPTrPZgZ/g1OBBaDtZzEYvFMBC7EL4Pi1uk+ERFi5zaWQxArbnUI/vTveimKaOue
r2i4rIwu+H6N5jvog/ZB08jRT0gT6aDuDW7Y2en6VStB6jFQNiZnoSx2DrOZtAjZG+hBO63t7PCn
c70BihqgePEiVNDqO3RHwDkNL3IsM38zR5ykkfFSFEEqx+cDWZ/ZfmqTMihlDqKo5qhyc/Oy5TlA
9eakSCTT+Z/t9fY0rf8T49SIUFe2hvYfsIlornO+rq4dqJYp9Mbcn8jpzYGXjbVD7RmBOG02KflA
6bhpmh4mt5jiyRXhuz6DXe3BG/uUkiePIjEMp0Rk9hWLB7jP5cKMyxfFNtdmoj5KGiHO5ejBIasr
IO+u4bt4GQX57kz6dW3048TFr8QXMywhhqxVS7t9J67jm20hn4va8Q8vW4Ibf4opuVk1C6CCOuu7
bsu5eFcFv3x+sRC6appIiqy8CQ0pI14DuSQUN88Xh+2Dfdh+lmkdBbDd4FVfqxEjfO3F+vMiZS2L
2Xr0FccXhD5WTpHY/7r2JsbLiTTDf/1qL6PyA1DYv/bjJjjGPtLaaXTerP9zMNuJqmyWInXD/SIA
pvhuhJ5CyZosDDsoUCxDkiCENo4/jL23wFaL84Cb9E4kG6grmSMlAQ+9X5I4kcHBXqt42KWHOlMC
p7UP1iX8c+9TNCozyVwMJ3mHWB5Ar04Cxsmf1v/WY4s0NU6903qer4zuS4qlCFrqU6NNpvRm3+eb
nJnAayCz430N5ANx+4h0gy4YD4ZPsvTuxw1NkT2a0ooKmqARwkttJaotz1M6n3wSy8km99CTiOCs
W2RJvIi1u0S2WMGCHx6/hvzCxjpu3hE1Zx+8AWBji9fB9HT8kdAOsSCfLqE2rbDyN9sr1E/CVcIr
urYBudvRpGMDL323fMPMXsUPwxw6DnfbuSuu9SgXb3yJX0wLtcBm7LK1x/08g6Vkfd4cCDBR0ews
peSzfrn+hA2AdtcnPiy4chwNuNKpaP9M46t8KodTno8N90DkmAnmhuAbwOS3WnlEcsm93ikzSDls
vlCK5U2z06zv5BCeNFMuwPw8iyptBa4MFCMa9mWtnadN/cmYsHgDyOMM19Rz2Uk7w6nObkSL8YVa
6re1XC5PeVmazH72dUbcj2XSUcAZRAxjdAQXku/9AAonY5UQzEKUrh5G6ELgmqkuTrvhj0glrddO
YKkw/MX3KJvk8lShrPE/7ZPIUoxe4/APl8XPBEzEXmXL65RO4PCAfTc/+2EmhEa5O4OhrFSU2DQ0
z1WZz1oa65HLiZiQ4/PKNxL8suYTRbUmBiQjXwNiGIXfTGefV1rBbtkuTQlk3sYlF3wI0sstQp4e
qhAgfzaq/XauZJKGnF9F3gS9vx5EC5ZG489mMRnLC6ksRJqUD/BiAW4g3DcPy+kalTZJ35l6Qap+
DbrHe0BlG/jNn8Y6hKAulXg9WH4gaRRTNsXodEcEAStaxHiEemL3F4Itvk6zakJx5z8HuhNNP1iU
yehg6NKkvGUKas5MXEP1z9gegdtXIeyEk+aPSNhfZC22gDgfyKKKq+qPjc2ehGCU4cDrg91/vEdp
zDUeY3ApNe/CIh/e+06lXEZfXj2SUUsVzvv8FfFhRy7FlMUWKGP0F4JyOtGG/ZVEIKbovm86L1sv
elkgX1K7RFD8q0jis3UGo1CVHqVO00rXLejT46V4w51amr172fG7RKFYxeMxxPEBxj6/fvnzB83I
zPzCQzbsX6Mqh8KBhyAbPJ1yzuZScD6E+al4dsMSosnaBxn492DBQ9jUPn3EMH5YIqsXTycxQ6xu
GYSeQyDhigMqVe4ERzuQoMV5KE8x+EBU4KkN9YPEl2SWstw/Pi4sbTzcpdQHQU+bfnmjmwUvnDQi
ZLd4L1W7UJEMbG57fKHRUo6zEvgDGX1WFMVCyVOa7pUYPE1McQzjSf9jSwGYK62NncuII7evb98r
g3Y9Yiq8z/OMMr4Fy+qPGi1Z+ujZyKyThRS98hWq5yoSe/osBM3FJ6wHSIon1qErgwBd16IleTLt
WaaNLG0W64ZJ6T/Xk2BK7MUVR/u+F8EbGc1JAegsLjvZ9IorDWKqym8rG3aaAmUASCnDhMOIyCfb
6EHTGKBQpUhH1yvZDHT/rvPgAYQ10ummg/8cgbXr5swq6Z5QG+mkA5GkDrRoKH45JecHIcf5WmYT
AjJj+5aKWeBfWF1bt3wqTvUGS757xb4+h1C1j36rtJB40s1TG9FpDyS4+JStO69gIe4UItI6eJ69
VlDaVaXdRsNcgKzWBXroLwSjfIKqDUF6+KNpYP2BE7rPjrf5Bj60NT5EAqBysGwT63PsMHjnV+Jd
8nfDKhelc19CQsqTJsumPeUyOIi6+05w84m98O9x0b7YXjt76ucAoZpMZeZnqlK5j6KVwZC3nxGZ
ky/rsjXAcrY8RbM2VWG+ylFAZqf8WTKdgF78lMq0zwHsXuTHlOgjY15p7uabyY3sU99ZQL0XrzHm
f9alyXNiZL20ZYMY+C3SVhbol/hxtaKqJ+DW+UNcc6H67szHIZO/NWqVpUHKICsZQ58Yf9xVrIKG
S3NedG93yq59NQFyKjfQ/tsP+iOZ6s1SxCCa33rMpIla93PNNSsMCnaR9lenwsTwwC2LLRq9l0C6
2Psk8BHoqlfpRc61s3jzC31/nP8hE93eD4EvYT2oM39lDi2JN1pLw2XDwtYhkNkZpXeyVs0hIXIh
0nMWCDb6igWs2eEVS/RlywcROOgiHk/1Ho2ndcI/7QY893WR2axbOW8uYNUuPyDaRjeCxvAIfXw9
eS2ODtfhohk7F3KWDUbtovwxqrJNXndMDf+EyL7Lm47CWzybgs05h65Axbx6PGqWd1FPY+mkm/Z4
LXs0ssuYhZ2aO0+0+onVwCdeKxjPlwkLnXU4JFMsuiTMfndFvJXu4pXb+5SYmDOcxMxDV7L/5apb
7qGgR5g8jImuV4LheB1+Gu3aaklV+b0aVYQ7SJSqqYogkERGzGLCSLjxWF4cHX3tQ/eTUKpepI/k
kOMLtoiy19FYKXaeAT3C7ozUZHNPi4Krb6gL+lPiXwlRrkcrGoN4FxsvjoscevhnZ/Zm3KwnuYk+
srlvuN2lNjowklofopdW6hvRQFziGh4hHD1iNbhoavJB84RN4TiNkdZq07fIjiCaIaqRX//+5BZP
1CvTTW1e68Os11dr5jvNXbav2n6iH1pgo7hqTa9jdcBkhaS26YwW3ivr4feXxvgy2EFCsSESGTJL
qMbQvAg/kEDEslO7r2iGNVmaWu6XoGvm31e9Q/l+oQTX2MKnHvfzuqRLjiWpvcfe5yA74Hjt+wJG
mcyfTQgSb0VsBYRoy/aWAuHx8wov4CEBZiN5FbqseQP/0OUetlbdyQE/mbpzNNQJrMXUhlB5hoO0
sOfbrVQ3uv28Vvqkj2+hiUeWadSflXo5F3C9hl91l395mCHnJ1KI4g/G/j968OAvb3A+U6k/1h0u
CIDWY6J8EELJEn4Wpk1TCDpAm7ilJ1vZrJdZti/kF1u/CA1PBebeaKO1U4oLB3kJphOynr7CldOD
3WMcHynyXAjAMlgnfnBd6HWqMxo53yHkj6aR5ITW9yantdvmpWVUmjjoIZBRojW/wz4vTH3wx14Q
F4DAEtHaSwGtdbbPGAZkhurA86K0n/thgW/ge5ZFmoW0X2N//6Nnzycs094k5mojc+NZhsmpOdLK
sDfyDjHT1AkSkQXBnPKcLOOU4jEZCUDbxJAmjJBRkNEctHuGYu1+gW0vs5o5OhngwbczPYlWn/9n
Ofm/07qYwRLcm3ytKBhIDkdH3jAJzLQwaWsD3FIZUaEFiiYXaJ9vR1Ip74jmwqwXjyqDRX4X7HcB
r0cRFB8JXMruIVO5YdZB5dlRpfuO9VD4WnRVYiUByNiZhqDGxjcWdPk7jYzzCMhXajbegE4Ayg0S
WKkV9kdVv2d59nyFV9i2mIHrgbG1FKgG13EC5onWkAcsdO+A0DKEDXRIlLMA5P+KAozcMo3B1NRz
VbxnvN5cjYdT8jhcBHOeThf5n5SBZwFmfntTogIcNPIpEHlbD0Op+gbqAO0k1OeeFRBKXvJPw4jC
fpxn+PM3i34QoR0QJLmIWB6ew1s+yVwJ9zqrtoikVTFtYHRCnUfk8U4CEFpQtu80U7R/bp8Iprj5
gqersP62zdJlqVwpS2W6oC4+Ltg9ZYuY76sZsF4BZwc6cWCQ80FwTChGV4h+da+7nKju4euaCYcN
oT3ooA6urhgZNgrl9GmAmmZ2I29gaLWCDiF9g1Jjh8PpR+fPgjZVRKh9+6y+pZqW8MP1GWo2fD/7
fMn/fVyr+PZULYfHCasANc5pBWDp8YVMvHpEaUiX9R2xKInJi8G5dNSOAWevjPmnavozGUKfYRfa
1bzenYJmPGA83jariW26yOa6shSNhkqMtKppGtkJIjQ/R7KZR0YTXTSsbSoMZUXgKclTco2g4Y/L
rXSX0hAQunebpD4KEQAqvnfKVyQtJzQOgNFDpVmM/mzOTO/BHf2rwB/BYcYfwFjiJOXTBcjF+KXG
TA2dujLlAaA7t1PZbYBejU7T8Mk78mWA5m1xzjfqNjEZCPQwDTM2VAMerXVlQBymzE28sZSJjzuO
2OL6d+AZDcMTGoEAD5GCPezqOiRUVFsIP76qV34Ug7inYa1F4fkEEs8jU6oCUiTPO4gJ5qAkzgy3
NYilL8AkHd3WzkEMp9THi8FqdocRMDLVZjUA3d5O1PLwmiyPhj4qTWwGm0kApnMoXasQDX+/uXFZ
iypTmnXxxLuDMn8q4y9SkV0kj0yKZK4jq1CwXp5gZAFIOPZ8cnqbLrSqWyPfvbg/jxUMDF6hRZro
BJCkVHTwYW6vWRgoR0cG6DABveJalZ/4GqAUfS/InYrpCgstzAYF47w0X7nyoqhqpjMxrYms+8KS
hw/XiKfYVoPs24GtAT7+c6puHkr6Fvun0cPKGg5NuzyIGwwH5FjmiHQAIrMZzghj9qBKrr6pkxsY
9vr33fRPudKLx1Typ2VgpMCbHAZRvVfd04ZuG9ctBf6aKvyITAuF5xr/I9oga2yPp3y3wwoxvPuS
WkLzYdbk0qv/f0w+yBd2JtShlfENZ2ovYgTCPK27w5GOzwmbngXFzWmZ7/ABpIk6W6tIXEj4KhhB
e3XoXCHBR41/Q/SKz0saDm1xusIyjDzTPqOOIuKuVHErN8rin72s4l0xP1qWmRPtMUVEv7cbMDdE
7TNWun8qO1GoTYmOcG/BZ1huZwyTKNWd5dYgKJU4ZBEZBZ2uWdYU0Pk431XfYOquVLkkZrq5NXeH
SPHMPPG+MfnNdVgbvqgicLmj8nSEHuj8mwbBucpxBk/tULct484qknKd6Zk1e5i+gvDX2nBDlV/M
Ki9ct4PUZOctG4xwAhf/0yrNwPdLwneZkdno5Nu2Gz1RdHYhdlV7FHNt/t6pcsoGR1a3HwoDllzT
EvJ8dBfQlawZZHdNWjPHcVYF2BrzTpIeUUsHnGd6cxUPhgBJ/73R0qMzTAQxZeMcmO7B/XKJ7LbJ
YkHKJHLNeA2zHZJcGWVihHyZ8GzTDRqafVNrST0IARhJra9CKAU8xgF2LI738VsH9/4LsPF9KdhG
oYZaWWSUpnSNbkt6ayQl7Sr/6YKtGoBaMEJlCv+zCgJGsZYWOCO5G/CALkzucy4wasPDeh1bfWjy
wxykRulOSnHytLAys1GyMQangTFNfxwtX1wrUR2lUKji4HWqgChghWCi7lJBBbSCQzxtHNEDrggj
qiYN4CUikBDLgpBbuWKvCaQMiFLRL6IJVeZE5+zGXoKhrJS/kRcX9O5I2E+N/Umi+g/29s/5N+bn
LEcD0nqPxG8Zy32MqqHN4/24uvzhTr4w1xWpPAj8ZLsLEGwv98je9rXfMF2lxlphGTrhqCcXqsED
U+X57WLHCmy/qiYCKJyUA2oVq9Npl6dFcqVCLa4iabFhemmMxaGZHsHuDchoTM2s180fIpROU520
Zho3UsOpYychGRaLVPD2xatpHui/CMr5dhxIh4+/nd0GVS+53UsXTbx37uTgWJrEtD2BV0pLRkM0
a+peII95fKStq84GuNQ0oUI0dXc9tw15T8EX3c0KgpQs+kmhTCsnhjU7GuIp3HTLekVq0viQKL0T
1s18jepQJ8sKr7H7d/4gMjE0VOodn5m6g+BWl6x6UO5Tha+L7blnMxsKN7zTZa3TtaxapupJGHoZ
MiAkF9lLgVve2LUkJXO6WHHaEx0Mtak79lEF+Ss0H71TCL2K7oZvhAlzXuFCOTmHP21X1Nd+Q36G
e7MpOfEslrYYP8Jq4LCXPCKpUKIco0LrYcvRETi6+XiaW2WLyTRUD9yQsITc2eDeIgfnrmCibaVq
pgbwPR/p/BKpzaYXzPkOmazAue4puZziQPKRGYfDuxXDTE1LlxYKxW628PXngEvQuiB4NBwzvmKy
Bpb+TsN92kZVJPVE16CmEseNl9T0vkwgZrUsPL0x95PkNUrExY8BsoEt5DL30ESRitwySmUucB5s
9Oo/9ulgiUT3ZWgST4nHrChqSjuP7S0qImbMiAmA5Ze5FyFLC4owurBHfXkyHBcOT6DUln248nVG
0WBnd3KGETtT4d9rEbRupCQJ95w/WONuiZotC61sEMWSReAJRjwSjwyHVfPO5L8HL0ze/HIsbcvr
sjkwtzI8Qn9pGQ7VywVWC2hfjHEDkudbRd2MBwtyHr7tD7Gt5PLEPKXK9lOUWoc+ClcjawXSw1MS
dAPiENPtQgH+3faiWYmmHKcPaAFLEuq00YR/zZoSNNkEUpKCEM0DTNfEC9kzznSOQuj8ABfsiPCV
dWdYyaGs1RfM4sWBO2tfR0UFy6eQna9SyUuk/3Jjp/H9MK7fx0s07HxkIXE3Lfv8vzsIvgUqa1wq
9nIRTSPnKwJ3J2tyF3yKiF32KzCSKkiK+LivtxeITXdJ3QNj2JVDtdKQ8NBqn0+rH7bXNqg7ZFs+
zaJ8Off+0WpbALAEzrR6oavDuLUkG8Um+ddIVcSS9HO8rC89BFMLZ/bqrz86eqgH7PDNYItLPvq0
6XReJTEPhnSOV0EHirLN2dFWPEycrQ5ePdxDwhDL9pJ4CMI8W1Bd+1cNh1xfChfRh630eHZr2d2g
amOQhLr/1oJq5Ou/stUjUiCxJO4J/0+Cxcu+tOqsYTGlP2i6fB0ur7FTF1wlYVwVATjPbdkM/jwq
/waGIjbbazP/9sLqgVH6lr0dfxVsHKFTGMyazMmAVkVPez9gkFgED5lezHw9evRGkELG2Oaqwuku
ZWbVvDgBXl2TozScA1DrJztXivuiY6aBP5MWUm98oikiJM0JD2jT5673MKWuO63oAYALXe44nMqz
9aMwsiMy2L1Z50ySZM73zJQa5vhn33r5/GulusZgCYnWs7r78nBY5NCgdWUmccgVANVFjCB1E1BA
BCxDRkXBcP1+pyHX9PqsOdS8KUOcx2NVrDxqAL0XTkFGZ4MGmcB1FrAXCunKgR3nyn+I40lKJfVU
l61NvyMinaM5KTpQarZThnvtYiUACmVYspsHM90DZLSaTyvlepsoFAd4i0PaXaRDyjrIzC/VqoLA
C8D+u2uIepecQvu14703Zc9KOrC9wAwYgAhHK4QbKoaSJmevUc9AESR1dYh4TP2CnRUesQaQ+kTZ
z1kQnqT77J4g84s4u/SNBE2tBGyYfXFzhQM5xvWrRRPSVpll2GKSVmIoAwdHWNW/mvfpZat5db0A
mD4N2XeR6uMBRY2XmdKEUojHaTPIZh+dZX7hBLKVYfqCeKHWc1g1WxaiYrfMTekVk1sl620npx9B
STfnX5yJ9DiK7n2PyJDZ6YtXKtQYEtJN2jl8HDMVMjQhz8j3Hi5omgk65XgZfsnmsh8xwK7yPev4
6VFNvaxZuFY2AtmXfJcAwsIKQU60P0iL1WGg2SxhBkv6Qx9c0rJ39xGgSdIdwjDMEGsdoEdNB0x8
uFCqvDeJQoSu/CdUYxrq3iRPmiBynx6iC5QUZMPBFv+9z/vYzCvgZkz3mHRuknZKrGgkMRGpk+tM
GMAcBKgVTonHq4MopcBHuUQFRxpbvttU4E1A7E4XwwJnaqtsx8fF+IwZS9K85iXfyuEQ6nbXdeRD
QqDJ8czNis4H09mTk/1owXlLzwoSL79Ht15+hBHbJQFa1brAGzZA4AzOVT/5B00cEmFt28BC8l/E
wpCYviO4fsQBA6AYy9ugR53+EXHq5gNI2jyAdjxbkbO4WmEFjNXHfiLW5E94YOLhWatIVKnrwkyh
5P5/RO+cp5blDnLZJfjls5bS+vct2pS0Am6TCQk057UxA2rFtIalFaQv3e8zhWaF2amP/HHPxpSo
hO/XOxWCME1tHB1BWZRsv3tm5dCS5kKm8IrRNJQn5nSpzY+7q+DT+Oe4i0p36VvDD9kj//32tk9u
IsonG+J2K9Dqh7o+eNUBnngTOox5qdRmWSLlblaWaF7Zf7DduCt291JkFi3ZxXgV/w78QzlFkWaD
WkOA9dKIhQGdLYJehdQmzVtWVTy/BnyfKMLfUFEi9RS3Ab756g/va0xDWZvfRz0T6DZh/v5c8kfZ
GH8yiUzrqlAGZJ3+Jm7t7RiQDFL+m4Y4eZNwOF+9b/wsLhOH7tDUjbTlnRGCtUXpEikwiGKVrVK4
EUH5rlEbQVTlSrdnZ+cSFeryEJ2gjYyJ/bcDWgExcFhMu8XeCvCRzYTECVuxTRu/atyJrPIIIox1
xpbfLw03FZmB6zelSNKRcH2aVj2RNDB67JFKFTIMVbGMRi5tZF+aYVGllQtsnTy4tUx9v76cxPsz
sQFyx63JXdk46LFVNW1RjnMdPhTDzVocG+yyU6zDCh4/ATj5NoeuqVH5fmPnE3rspgT1UNE5FPEf
4BTXnczZUhDJp5Y7XIoMhm1bXRdXt8gohHg1noSQMrvkgDNQB7s2IRkzzJJeGPm74ojTBQg2/v78
tnyek0s4UM82mMXhMrflmUpA7cNiI7SkwjPod8ivkLwpTyGNwWYpy02JemDpIN7UBYYOuM1Ydnu+
hs+8O/9sLZcIjH0FTRIEQgujPZvXCzMp0A0wQdF1hrO62eeRu5c8VS6IrEi6zXT/ySDGHDKHPvq+
s3V+Osqn4/QiXP5BuSIWTXrI96GDh78i03Yu4pMd/qYa4fcKVcvOPyczbdvNGx1dzuVDGpkvBgfD
/lT/C1Ed3jaKM/BUtRy832JW2mwqe4fZewPsG8ZkUEGNSZnF4DVcc7O8AXdwg71X+cU7LWDZ7GKX
vv2+9ggfDkKHdyUwu79T01Y2kIDbEvO1giqUcmO94WB7219m9yaxA8/Ls7TEOv+oXczBfJrV+sjv
N6v8bxa8ls3FB9SgmfzxEybt7Rw6tG2eBUmUEiVHaJkKN1jm5GMUwaXORFOw7UG0VY98U8vLAkg8
a9uB+5wxXWX+i2zEzq1lHzdUtPJrfzfe4lrvLV/+5c0fsJCK8/GaxvmF7+WeuV5KryyiFdD3hW2d
NM9oVp41gOgan/+mFbgVbD4MZlZzaURYM89spTGsMaMQpWk3Ay5ZS00Gop5hzsyQavK4OajOAObg
lUjovSv2bKiXwbrsUVVPFqD9WlevwLcTmGEmNwHotuq+eaCIGr+8IetJQXn4Ypo7MVzWa0Of3tga
g3PqjhVh4cE2ZTRVr8hpJBomepLvoTuLPXdSL8CcituXkv+Np46ZLkAuqwA4LZZKJYhvkHtSiR9g
HSpYrGPvYPHYVbNVQM5I8WVu0oqN+lt0ukybv4kRk2LKiWGJJhD8wHc56OIV4ra0zFFLNVSQAAbE
hawd4waETrgVUi0YwUgl1Cw1F4N3OHPWt+u0Q1bkvptIQob/OhxsbIHmkqXuYxi9X6qeb5g+8G+I
5wNY1r36eYeUK9sp+kxEhxSMSIkIgVPUEU2zlz6xQ7EFMcxMLSkqOqGFG26m86r3xgK5NAaMbzoh
ZEDFpPsmt8XPGctJ5SeyCd3Eb3Wg+dCbP0pvqdYAt6pRa085PzvSaxUbCeq7fuWq++ZzMYyS3y+r
VxwwcTh6i+WhTZ4fyU2pT7y0dhsEBgvmqn8vD5zfhYKCWXZMXm3Lrtx87fsfjhRkMPoDEaV0D7JT
3bK8duVaB1ojgSA3sFZ4ZPI69PnHwTCxCcla8ldGWg2hdTzDmNiOYUB8hTCdqP8OeMrFf6Y0XZex
xpML/Ty8pNx/q7mEWC10YhOQ+cxP6rxJXxfFDsPmQTRECD6+AFRURBe997BH0zp4D3O/7vQmbTjL
ESKbBkPBChPc5vXgJK8lxB46Mp/Fv/2Gkr6tgFOSW+MdjuDuBT4K6m/ORdZhWbvGtsaywyurkGzi
dnp83OeAnVctuaZEOOlO04v5t22rgwFOqvmP5qnZpjy6APtaZhXCfWHjuMSqOKy2nqRGtLuhQ/GY
gyc/CG0Zss4q1PQ1+t2zlXmQf6IMHCR0tEfxLn+ef9k/cEaQBbOLd7RUobO3SAWrXw4SNG8+/psl
0WSZJmrtIiaALfttmj+WYBe3PViAQ5H3gI+G6sBekEyhnV5j/uN3ETT7zZTVQY6qIavMBQsr58Lq
tj4noC3MMhWcSbnHalWGGUzRdVKjIHF0PvecHBRYmlmdCpsPKzgT36hR8NF/cPBc3fW2ehNzdpEK
7LsumvdwKSG0S6Zr1cO1Z3bXXcfWlpJyv6qf3UY/DDYLKpLAMp8W/8OavByV2tK6GgYEszKDVjO5
Dk477kR+krCOiJOCOieC+EdXfbMqHS3cFdXjBikOMFUy6ZfH2VXzLQRPOqkuYfWkgQAoi7KtENdf
4y7MDCii+KyPbLpVTXOtDwyCbRF0iChT0v0K4s7pOwCiIM1k9obELhKoIKsQADoGc7vZsF5fyxtP
XTy+uPQRRJGBwf1BZRMR7E1Q0WRCcE+o6bAvh0/aoW2hK8ua/l5Y5hFpBitKTV3qYB/e/rYj40tm
eyTxO8INnVDd3sTMpcOAuZnb3vyk89avIg5/+w6QEbdpTBTfpACdheiZUMDU/764EAGQq5WhGw4v
qNehl8PyxF4pUmyedNgN08ZaGnFgzjU2szLu1QWCCtE42rultBUZsQ5ArTMyan/w1M7yIt5xknH2
As0GbTl3quloGRC4w0fF9K26kXMiSIWSjBe5uChfP6EweB/EA/lRQ9Q/hvCAHa7poOf7tFbUpZAi
noHkNlg/oIkwNXD02kZ3r0U2WoAu+6Vq+JomfV1yzMZrFFuUSIKsnDtEcqxxwkl2xEb8qgZWyGVE
YRhT4tqdBluiwtTWwSgpW4ujRIP1gxbZTyaVfqDW0lk9QNNE+Af/wESvVr+Qylj7/DFzcEV313xM
G+hQhyFNQpSt71B7Z9ZuUKBOY9kqstm2rs5PesXiF32oX/05KDXYiGit66/GS4TZlX3PoT/KJf3j
M9U02KBYlPN0eivfWaU7ctRxdvMzeYSFoQ+jqVEMzMR8yOq3DgssfTT2KNWUkQNFYr1ljaWV8jGg
gSnb2OGgEc5GB2wm/KhBu9qG6EpFQHtE9JoYwVFqo39JwV7EpqP58SkWxjm5JkXOBKG7DlHJSpOv
YEsUsz5DQI1ONFayGYDzLawLvXyLwrSJtWxTinctMCzEdQVGLs/IpT7/znzAYXs99WaJJ/NHjcfB
t5+JOve7H+PQAw7JKQczYLGwCiKr3QGiiXcUNWk5ath/rhJlKWOWdlt+XMIYifUSWMQ+Hw+jLy/8
WgtLYdQ+M/QJr9JMAN0UO0nmkkSbF8tpMBI2weW9fRfCmzbk9UkdYUYKsWaIM9oY9oMK+i51f2Ri
UX9ch7DYVTmMfcLfMcwkA992Sb+Nyeu6w8GXT3U2X0BH8fHgTVvnai/DZydgV8oTWERzQsvq12Tf
kZ1Z6yfgC3vhKM9oG/Xr1ZG026AFEaJS0FVM+jeuhMA8vRogIGNNFKt6jWoTGfVtEzN0iF7vlCzE
eknIHtzzs9Qqjz5utL6vQGJdx48APL0+lawAj63B2LIpI3PqH/6wKIlvh4v8p4D3cVzFhLCZTkVJ
zcMvezA5haz9lac1J7CzviriJxHkdftHFky2WTam4wgKPI7klyst7xR5dAa7z7qksuqPyiTeWqe6
DFhVEqmiysKOZ6nh958yOYDuhCZskknNgT7eKyZoEuonyAblv/pRnKWEgWt7R/MQ3Fxg2d1OdDnp
gutcHYOC3w4woxGN1RvLJJPzuIoO66NfR0YOv+3xbODWR2XYr0DVxFF1LNJSBADtnZvXvUiQRo/W
sWC3dvXSO+TeSGPGLz6F3oQvnmp2VSGPeOPb7ACIuHynmEfyIkq284v/VviWv1lRjyMHajd3Bj5/
pgWW37uec7TD8mTXxqAKx39eg+LloyMfkks6VUMddQ2jemoOkH3oVQtOtHAAMsPbwZ9wlg6JOCh6
53aaivw8EQTMfAiFC2gnww/vuv0e9nkG4c621ikVSe0K1/c5ZojujpXRv/cNqDQ+iZ32LCSytrzm
VSWQIlkm6Rm8mTyi1WmkRJaWjxmyAbv8rsnE8TLTdSQs/FYO1REXP6ThmFIljzvSmyHozC6yMPqJ
UCq/xXtWK20Xxbk9sjd6qgR1O0BaEThsFa7g6auSvr5GMqin4gStAtGL7okZDF24Wm84Xh4auMV5
JBwinWRZOujAu1y46BkhvaywbTrpLluyR6KAa0z/pnFsbIxQz9Qj/Y4j2rAE+TpkVNWvby+tVI9u
qomRDgofa2mimSyxJWsCvr2ztXinyVbZ0HNTMYj3K+CRrC5yLIVgo39ksuqEiIH6x2UZJXq7NDxU
zRcoO3eNy4FBfvhNoPZ5FqeBPquhA2tYcb2Gubt2xRN+TfIQAxooNMaakcu4RtoTE3TbhpfAAiY0
RG00waJsaahy80gfLnRh/KMt91uK657pzhtftS11El42PqO5tOdWUkgUSDyHKSINy2ZnvOzqm9QG
JSxOGRub82Ec2c8GeczEGsmyfjecIlE28PJ48gzzA7FrkOTfNCEqWjYAea3br+BMWqzu4D6Nra09
L9ppCNGN+SY10XVvxI2zGieQJOAL5CSO3ye4CgySRbVoI2O8BCRKom+es7NXZ0DdAL58sP3JWOZY
NjhByQWBgJRWZKAO/6T5WlHKaMkgs0e0K8LuG+wxI/nC3CdN0BqlRDCaIdSwJAtb1W35Zx9Zn1Tw
V2Cgg3e2KlDpzCTDrDJuXdn2sOJijLE/yuBnpJYyJZHgwVuOzmlk3vz/rKCcest6gsoWTxw0TsU0
UmYLLoMe2wlng0Trdm3+aS+wgqIkXIVSxZf9t9MC/suvXrl/GiSD4Y07amYjohyZi6R5YwPX+FcE
Vy9f0Wg06gneu59lb2lKD5w6g+ePh9/4MrCoSmeMb69nOB6hYkr+kaqXWvW+/Z2fzqpmZVA2HgZo
NP/WQi5JdphjdaWJ4CnR3G/qE69jYPFRuTG75JB3WePzph2lUjvSsgEnQC41WR9zXi9SE/flQZui
dWDVsnN9lNoWc2WgYRk78Aun5nwaZRdmrxjkJR+hdKeZg+i1XAcIqnDjDE6OnBXW8tXOVqQp2TM6
e5xXnM4o5q5+BY2kEFM70FKe6hrFIkuArXiVSe5XqcBtL9C2Gm5VM9gg1ZA3era+88aNOA7qc/Q0
cqds6zUpaj3QfxLpwb2PbIeBPFkiCi4AiCIh6r06E3RiIceX7vo11T8trkxIeokRdYg/aYvzz/VH
Dz06xU0ZgK1VZmj1rFM+dKR8e0pZsWpNfc5AjyVSr8Sz62odUOCQsjlI+1Qlnmwf3fn4vx50N/1E
PeHgNJ8E+NRqv3v1blXOifsHMei8k6IA4jS/f5YSl/SBUYhhHscEnsSD/RHY+7qmXqMfRXY9jBRq
mCZcpfYiMGgwTYFKOiwYKevU3szQaEkm/60LNVv1LLVOkQKq4/RSCe3xUKLme1ZvJzPNVWxRb3S7
WIsI0EqToTrLO8KEHe4RoABh7tdE8couzdFhfqc3AWkuDy82cGtcYbaSw0acdSrDInkn0yJ3amaf
RawBBZ0QKrKWGl01+f0osRJIX6GpuZnbTtT1hOdkoxNQPnJ5BNfv1jMpx+ypvs9wa6blmnmJd0Q9
IesTjMt0XKD87iSX5G0vEhhPdU2PFqcQ7r13dpI09ZDn5omRx9g0Tfq+JUeFE/8aBfJQaR4mqOxj
kNR20+Ovt2rZKRZH7jnBJyGUKb5iGw/B9ug+/lREkIantmHqQzGpQ4/CLF4S2717IqKCAxDGXMm+
xY5Lyz7EGubX/37ejRHZlO3mZcRR/Bz//9iO+LTvI73eaIIuYJAgsYRtVCJW02FhAgt5SBbFWwao
j8q8IA4eI09iMFXAFzGwOAXBiXspN/O7hiO5uyAZqbJrMOx/LEnjxpdLz21fk0VJYzvwUrIRtyGF
75WuuBMvFDfG1stGjbhXlOnmSl6utlPEGqLFRUX7Ln1TBrQ07p3yCh8fmjqCkyLc1I+uqQQtqcgA
iC41n8n1Nw3lbSI8e1AX04q3AqiMbVXhJUR8U2j48iHLMaTAVOocyRtS4WOExNglDZgkjtExpjdN
c/V5xaw9l8FmwPRcV04GojLEylnKBrjv12jBy87SFUHQKQancZaenqeb9aKIyoheNmjqlraGDzta
Er1PDqN2n1/bVZl3jMxdOAcR9dbf03fYr11PBUUY0PTq+zeAfDZPHAPTdJBeVlhm1h/5/P2sVL7r
v6ORDXggePRzYXLAZJeONdauNe+CbpRwljhJcx/oOi4rRKQT72mxaUCLfWnAhB6sCEyOO7+aEm8Y
+vaH1ce6RzSPdPjwtnpC6ay/cu5GxiR+MiVIdECJx//xI4m+DQkoF4i3LuGqvvGGvv8u41//PuWw
6wrZLtLOCNKW0EYnKWtQVAb+9TzYI1NAp0FAW0WLLe3dXpDJhJb5z8FoqoVMb9iYeKtbO9MbafBc
N4DjrJzC2eS2ML9qiFWiGqNI0x2f/Quf09LXuTeapAzYelMTeTp9VmRw5wXojGNCbkopyx8X+Xid
vJ2Hv9qAWdquIv1VgNLL972OTNXAWhfmriHqnqi9qvsdQAyKJLtk6ntzBwiPO+gZA7YDYYaEJWjB
p0W+qAK447EsMtj9VHLYBIOPq9WiA9adtgV60ycBPJWf8fG5PldO0xkfC8j00SjJUE25GgOZ8O2C
cw4Ss4AKnMhLTSlA9JyrkT4KsfSdsVXMY5mfO6W11MPjj9YA3GMZdGquCA7GaxrdDJ3CUUgcYeo1
UGi2l9vt3u39s5OQ7ZVdWxD1dRDWD91cGi1Kc42ovNDWV3993kXwmDEokN03W2OY+u1OSu5SWuQ6
sWB8jxMgdUprRyR9Nexbq16XUK8ycTk2YcE7sOvSQZQAMC28mR2ZYb0zfrl009dFjJNi8OANrzzs
/oYTY1EUk6NF5PQ92f74NCtTtpJmdMzJS+gAXa9P/5+2UlIj4LCGEO8soA1Ouu47GQFGebbO9RCI
ijDZP1/6MOQGi5+mRm4QTVLHL2XmsM3pu00UOhACN70qKpduA4KBA89RGniQ+fUqTF7U6JcE67JQ
WybfrcWJZvZ8WEYpsMn58nhO3QYWGMfPbPN8TpdE3sJsPzNOIPHq9FEQCDqTMgtktxNDftYPPJ2q
W1HIKfVkmdiv4R3g8IxhiUWTPC4kkz/eU+g8ZzXSDKQwyrsikQIHq+ELKd2l5Kbvi+OtjpZkRdmj
8h/QRi/Lr6/MS9NCSic6Dst0+zXcLvHWmoucClJxuaynGA/LDyg4kbDoLTS4QiFq1uXjH7YF5+Bt
cfOXOE6fPhE8kjO7ovjwcUIGHS6wXgWm31v5kze78tyKGPGw6yN4vGUASS53Cm1ElIgH6S9mBiDB
W1ck5vjB1E2wX/88a0utqnwsP6b/BbUe25g4rQe5o8trP6LACFAjzvBsVfWjALgRheApfjzcac7H
NWjPouX9sOlr3b+q7EY/RlpFpS4JlUUJdmKaudjg4gOFZDIr47on2u0001TqBlmZgRNbd+NaBcCl
Ac5G05VNVpYd6nA72oBlo1ABA+ejxGxDv4nKtmJgfSegIgUjjfF4aGyBlttPnCq3a96xPIakbobt
ZZGszJb+++4QCEAZk7L1P4tfU1qu0+oXxCntgPqtoxnkrKuMgP2GIC/JHcaXubIBnzg1Gg6ri9ga
Atg/yPWYLNC3lYO+0a+3xHb3CX04rM8aangOOCwtGhDTFx4TQCx8NRiGUtiV4suVKrJHyf2wgLZc
LJtA1+tdTJbq7CtXFmQ8O5n46X+O8PXuOVFWGFLQQ9TlE3aKCEXxdXNllfxVb5SX4QtIXdbT7mW+
l5CsuZLQjmDq45OLyeiMP9LylviCBy5K/LXCxCx4+bILKaenUr+enu1WzMw3tOvy+MDvnG1f/Yb4
KR0t2yNax17s0S8GX/jYLav4fWXk1NhG5qyGnmNNTbyds7vhDbkp0OCzYKsEE50JdvLXWPPG6SsS
hle4cF+WsYaFrmUqA1uTNKSb/OhYtAUWk+DVPFX57qBh1swHrutE0JYEKmaEDTUWvPrpGDaYLf34
PQ/4pRGz2WkjpxSapEizl0S95i8CDgaQE/tVdLorTiFefs7Irj7reB0TnuGcPwkD3lmaX++71rKC
DDqeFOmP2fSsz+oo+P+MKgCAoKX2e3gD7wUNiOqwfI74HxgS8nnySGHmSHmqxoZyJPRQIwLEMFpb
vw3W2Upaa0z0kxm9L7A2NjqoyG/Mjnt2MgZlQtYKf5aKPKVnptdUKUbEA7yoOBYAzftCGQlFC2c8
2ScZxsI2OmwfYNBBwMWI88GsfXiB9kZYSdqDwA3+FYA04wunQuCysLs78gXRDkYyq0TCowx2MbNP
rqtYSYWR/qQJfSBi90lt3wibXUWq2Lfw34NTyvOSzGSCoVAv7yKGbATZqZHvcf//5W4v2BOzRNLe
dV4amqKp6V+i9ldCGgx2XHGrQJ4TmjyoXENgWJg1HsGeYb1eORWTWx/mFPCv75o54uZJuumA8p7O
EWXncjAPCdsQ7Kle3yoDFZ9LB4vdVHSWHQCartxSedqhDBCWqbVGgTFotpJJQpG+wbMgWT2+CqDF
FJ4/QBfvSm+675mLM5Kw0kLZ/L2H9VQwAmyzD7FLYJO1iS9BdeApDOcplUsCvMq+5KTZgOiiZ7u4
xcSoReBc9pGCluzZcPfuUx8l5XWFo8BpclkfQKoQgSennkAhiZN4WhrafOkCJ61m7cUPmTlTsJ72
XfEKHPcvXnd1pcHbcTXHlYzPuXv9Bvkes12wfHqxCatPSKQHj6bz170LUduQA5Dj46oeroZ5++V6
HkccCzvyjsOSsnaO6cq2mZA3GZtZ9vAFALr07hmjYh6sNENuJxTjlWk4s4fq3D//+0LCnZpWUFVb
jxMo02MIBzqJRQjIyl2hpQzADIJTPlXBUuPenaSbHlfbXn6wPFc5FvDThjd8a8pNOn++MZlLa0kf
vtSfHuZSORaGLbEbJoQsM6X789mRtsjJgYbcxRoE/2G68b0477k6apTx+3qhRezkMM4MgAIkqHPM
1NPo8p2KTBkraIOSh642XQ3H8dHhQNJNyOjlL+TbDdg4a70/aDkEDRV/3179e2gPHFrH8VvCCl0H
NB0G4D5ppXQitCFEogqOXXNAKUN1H9Bmg1ICzIdS01KVbb+Sa4pJarMfzjPykPoYR71Od1rIoNZo
gs5nk5KJLSmf89iMp2nB+2XTHDwMWI6/7+XyApq/n8V7kvuo4CYRl7L9dvrLDs9qDOP89zDBgTTx
lCJXapEOF/Cy/ipmQOBEBG9VxE9uTTbPJgouCB1yRRv+CNnGQTCdFB7p5UtxNiOrgXrW7xkh8IoY
8RPVbGbVJuBEmdVTn5MiDgB0/C/vJj9BMRz3X0/aZC23+dvbo6fegJY+07ez2452sQypZrcRwXus
4/I2hHk6q0vmhv/KvJInKLpqHvDXOT3qkVNAeDErgOhhgtr2p6cfl5LRKtCqLY1KOyU/fva6EXbu
+IOU3s4HknudojBnwGLK5x0SttLO184MnWgE+39l1pHXHz+xg3KachVHhSjORbY2gIYtBQlfAPk3
82y4ia5at9XYaranAxuaAAkFT0sYhKHkcw7bk5yrsocfkGSrwjj83PCDm5U1SzXDZ7lKvdUQlmpg
HJ2D6wpBCIE6DR0aI/n3rZ+HJNc1a2YH4chznblUJyly4hFnWruRvZKlvLaAXRWSkmxhG8mpKqJC
5YxTzTIvJ0d1BCf9AwhQd8sfEpaseVwuaW+2xur+MZIfvBlx6tn8BDrc/MtN8jI20vX8r9zHHqdp
Rfs72TY1zVGITwwC/OWic0Lsdx/Qe0mLSZfeQ96vqMW1mpYk/CRuNUXj9q8lRD2nexunWjo3U85W
92DyBbm1EmdNPK4DcRbBc7hwOp91QXS+d46gFSUQiBBCrt48AL4t1BpIRvUfVRTfUWb9rD9PD4jB
kO6cAvnxP0lBMjXWRBB8CtVc8dXczBi7LZDgcry8qFpdtbdK/6WJtgecBjUgtMPsD3Ph3qcU0gW7
d1LbsVYFmiSxRs2kq2ALuzoHjunXkCixG0IAOKU03ktd+bA4BNUUkRo4A6hqcaveM6oycShgnqB7
ThyTr7oMNHsC7KTfNLdu2YUCqywHOGXmbM60pq3ocANfPWMc8wEGWjg6PRlFqW3UDxl15yqbKIsm
C9bK7ETp3I/rQWrzZKnksHkr1gIXDuWkyiCwHaAhoTJe93NT/p3n2t63uUhonfhzuJ3uNEhAio8j
UJZK9s1c4EB0ZJNQLd/JjpNUnH79I0ZHZW9mkY9NhTxk3YLUJNtJ59m/V+xun3/FTjTiBpRj2scn
e2We0HCg2o9DPXrCx0ojwJxnUc0orznxXk/aet/k3fjLSZEP0KC8xNpeGormVKs4PoN5HAvwouDE
SEFRpm9Snj8h5RAqU0yIo/YqcRqZ0P9/IxDI6oWzEBLj0c3bv0cJDKDW2CXyc5xWSFqGPj3eawuj
uADta2nwSyXRsinkPwQPjCnyrJk79H0e4uYhrTc6bszTKjtIBIG8TLXp/Ngo86ys87jJDHkl0/WG
r2S5bmG5sseOc7d5ZQyLlFlW9HKATHTrB0nWuBqicIkAnJOZ1vnqDqnV6eBuQcguRvNEp5u/Ck2v
Uwgij3O/aX8jgH08SKm7ZHEh2uIdE/MugaiwXrlqbqOoLlLU0tbQO39fbPNmpzMP/JQ/4TV5ibrG
n7lqM5+xUb1QlsLCtfpLg2z59SCy03JMS5SHsFM3FDOWIhmWfKe+EK6ql8D3t/GfS67Pn3hhDs1b
8M4DD2gPAGmdUpzju9/Ov1phnJId9lomFuzfXxqEmke1g1CFKj+IRhk8I2X/kbdbqollJEfJ2pZg
aEdcAQElcej5JMTeY71o1SzuoGKbEC2y/Z51rz0fKyaoIseiUd07SPgARqLEbXhD8NJksmxcxfxg
QIBteVpbjJZ23WSazGuzDkqwU4pJf+jsdjKFf991YHhNu9jT5i31dk0tMFTHlKTSgDnK8umO1Yik
PGwbnquUx6d9Ql7VLfk7Sn6CmZiL5mrjSOrtDzoQ9n8qNYQS2phm6+BO6uGndGxNbwmkqj4NZ7Lv
WKH5ve2/NAl64Fdy0GC45sMfOTihIbnq4MEyPDVEP+7PA5S7Z4hY4Qm43+mbt3tZ79UAvB5MF98s
9OCMPYlmJN+LKvZ53UbuA6SMimNJrfS9Qkmr4oK+W9JroU+nmgsbaL8V0ObMg+QHooXy52qM4Lzh
BD5mwdiy4DPvD2g0TsQE/dsKV71ss97nv5G9qjVzIiAsNba+vTVRI3W0B67fkTw97pfTPirqs9ry
dv2HGetXYBmnSSVRNAt9FBINcRYLTOmvqOxHeUV9tDxEO7zsS0JXuJQ7PqEart2PegW6WH5nnLfa
eUtmK8l3IW6fSEoz8Z8i0+aN8ONA6SWElltm9scQo4ri5a5rdh1tVTKQs/sAHn/AqmtyoGoNOeFl
GXIiwEwuF+Z9pgNG6EtN7DJbkLtVtWK4W4f775bN7B97UCvAQsCkpsazEIiXYjou2WjMStXjz7qD
yegq9U6+Bjcrv/jmE4VPnsrG5W+gy2tFX7G+OcvqvNRi9YYalfvpqExumCTb2q5JQvgo3TQLcnYy
C/SvWDoXd+jLk7B7lozbhTXnUSBqZcSC4omxO7hAAzolQEEOykIVpuQ+FzM41a5KlQQT3UwmL4iY
4tkiwOQPCYZ7vkyGLOwg2J2xOc1BLIVd6KT/DhFMGA58n5pjQMbC/bGWxng4SO6YxJh0HtrdJCS7
0djvtFj7K+PyiIcDOMt93jk5S8NrG+XGj1IRy4bCRkiIFs3diYhzgurlLTHw5vmhHuh9+nyx+HNs
KwAE33lW1w8Rg5t3xo8Sw+MIFOxWoPTORwMh2VbUROowJUWM0irCCvqPnWL9FC+rLKa0e+G9yUR2
2nKawEd5gsaPA81jfDzVU+3GfZAf2lhicyyxF375bqokZUY8T71fzgeJJTqKJFXk6lo18JF2QCZ6
i4+zAmMdy+RhTkmC+pY8zARGtl3rRMbeQ9pwNippCkljrWBuj57RqHKAqMnzny6IpCwh3Xw1ABu5
o8lVWSUmFIo1tLtCbOyNiXSoUr4uqfJhOSmXcWRltvs9DlYvaF8eIlB0dPBTiy7YFE/aDDy3bc4N
o/lNVWcC3cSUipOHhUU9vhUdoTlw9qSzJVd6R39nUlYGwtAHXndADk7gLgcdbtur4vK5oS4zXsTG
c3kGRk9UzJN8CZgEM/QDUAJ4NDScSuDz0hegx9CKcDdKjBldP30AfkIBberpGzXwC6jfiV0r6+sJ
ZTqVQblZLPSGnmxuO+zdO2tMsGtgWbYx+Yjr70W/b2rHf8sj/y8HBqV9drdSpqaLqPDbPQHxrBNN
+jecQsNaXi1yoG67XRyIK75g+9HtLAB87McZGZKI5GPYtejAHEsRIsVldW3XHXtrGwCavAQBHBnx
Fxfk3ecwC4IBTnxqwHGiEl61gXIZ79txZd8jKgOtWFjZdoCwxA1nXxQ6WGMy4mbcPNs9V+5TWzFV
W0qnhl4t2gE2K9FfIr2fCd8CuKqOJYd6dpC/4t6d9SYDT6XxlmTZsG7ecPRdnX35+EvlOc/qBr28
xaNZ+jKnAewuvFEfKfsenXur0SJgqVQXsCLKtjtczNeK8WP9aKpKbyx+3vwBtk9nmIC3bpO8K8QO
+zn0vGcw2Vj5PL6malxw3QV2NylAODtY3pE0OSyGJB3C+umSE7l2mudSs9FbW5YV0+mbNAcvHHfN
US/RDBaS4pPUbJQs6NUOoD2HmhR/beR6Ak3X6JBAoKp+qdFIijgs9g69fTuZSEX5YOmEMG34O8cs
N3w82Yb/ZqhDBz4G2LHfwhW6pSYqXUzi7XLgPcfO++muVpektxDnNZ9lgxnOCNMtWvbQUxdekCbr
K0WSgcXaFJCytKddXBY7FwdIB5QAARLdEYqnmWA2BPbCgP/i4GEDjSA02IBgoHnRuvFTauOArX2Q
3L6YGze1iLQZ+1NpRHSvP5boYngqDG5N6PTdzw4lFv0wjLnq9FvhKySqIFgdJ5V2n1RLYSCj6Ii8
pfpg8tCKpmNsJ0LF6BIsv3FFqmOoaPryGIwmcenfxXRT2SIYTLr9ANnq3fozrmfzondiTykOcuD8
46cSEAy2ugbYZHLd94Jkg03uHr2IY+cgAo7QDJbPjat7lZfoUjSq9gmi9BHKyXH/K8nc8KaZQPfT
Or2RQYOQCfetbUJ+QYu8tSNE23TeYWOekzCBN3pA2RPlg/6A7qTWNS7ptxMn3H/ybLYOsafeCkip
BNP5d7PM2BrUIGhlRgb1oyH4Q+UbwL9LNLn62pyJgukZ4o/BNW8ZTFN5/iQ0bLn5vD2Fj2MX/EVl
hCp8huLR27qVdxGG31s5E4yyy+SeW7b4j2eD8ciL8l6XyYnuq5b9yMI8KMWumDHw9WlxDKobWOpz
o9MqhF2StrMT/kGnP6pNAGlw/G0ivynVYQALMcneQC758zI30qDGk6VTZHMUkNjR+NUQxcBoiau7
0PRXE9KutnOgrg8CgjXGAlxiZv1iuoVxLamKlosb6s3+L/liQvCE+4OBppH/NN7sw2CUmMn/OrDu
hEa8FpyorITUuRuxv8pXioC84uphO3VMT59/9DB/SM3BJu5ABKAuHU3UNI0EHTCh8b65JbeTL0XW
Bkg1tfrWzFzHOUIu9rESz0krREKLtr7OYhuUGZZnzHy44WcmTw636ffAuUCFw3rU39c5KJbRaL1H
wxBEOAOXiBNr9okOdZPsK+tRvKryI2HmvOk0QU3UMTgY+qITS0zS+s3m/Lnm0sXlWYu73Uruurhe
viIuTOX5ZZcZfvErSnYjtO7YoLYiJ4UkW3hPb1F9n1iHjpVTVgL8OJPm2HejP+E1kWkTjUwV3pLa
Y0KsPfxJVjJfEQiTZasGz3opfhkOo/P4yxKjwpvsUXeJllHyeOpTtrqNcNjFLojDwj3mrRYZ59a0
l5D60ej7898ri/ZDEWiMRiV/78rG+DS/ASO5XzNGq6tU17+ozsQEb3srRw8NdzQbyd5jsJWnTwHf
+6mqfykvdGp5Nza4t7UvMj8v6rV/22tKdupYy3K61RpFbky8F8PHzMabpI9PNgRd5i8fIHDCSUR7
hZyavWhqjD/qdLKO1pkUNev9J4cWEYEmW5+iJ2uhzZB6Q05tTHXhAewV36Iv5owcujpjiJuiDHpn
kdfWy4M3foi+hgoR19IjbNcM3RqQdy83PWiahZqcI/WnaLGg6ucZCynCEkdQ47LYx0E6IlzQr/rb
MhF0cYOzDZWPzjzukHBA0lbpTkhb/xAjIZqCubfS7+OtHNIJa9e17daCMX2r5Oy8TfEi4flYnbla
Tq4yrFvX2olNM0p/xCamDIXsdknmUmitlMvTqT7vHi3Wqg/Ml6GWTqHfc+eclcajjwy4x4A52NkJ
70g5PGOvKBEiwG2e2OwTiQTsxiB1tqKtbtUDMufN3+SxbSgGWXLIDljy2nrkCxb/JQUUy2873Otb
4/8hiMutj7p0VsIpWpmcbPWXqc7Q9WZZX3SiKK4UfMhWG3RcWuLfrtEaaFf8/FqAOAS92U721wNk
e81maeC3Q9dhEt+jfqaBQu7j+n1n7pucub0Yw9tr5gF9nzNVHx0kMUgtwSWMyB9RStK/Kf/oOLLk
L+dkn+FVMnEcnyQUC7YnHOPwES6IvYI2gb8IbyTFVLuKXHSRj6+inRPYzecnzyN9SlhH+MyYs22O
nH/Sy2kTJIUWUMjZ49ziMOvSriUHIlTM9iEMMjvMhPlsuxoBDhJmChvU1G7mT/NH22BmNftF/x+I
mG482vOqM1RoVCAmpz8eBIrvssdupqufmWwS7G9DYAhr/qvoWR3/laIvi3GhysLeFncjMkCJBIbV
Xjvb6sqDBHrAr3fAROCxbNWdBLiViycQ0/vPCYFAriPGhbk6sOucG00s4B1wScVKAY1DIczInHCo
YQklMG1kTQaQvBg8HicA0FNYx2a0cqDBoqykivs3n2ERJaDDsafjv4CKxJh8XxMiYlwNI7NpozOK
d2/0dLYAPfLknI9xb3xjueyl3SzHv8SUX/xD/ds/hU0F49rt0IbwOgpu+MK2ZlA1fg5OhUEdwteW
oB2OeRlToJKneCAYfeNaY5BwRj92EeruuUslpybNa0G+9HJ6is33rxow4V5mB7J/f96+HJvxwkNo
stccCxXx04o4iaaHxlgGjbjslWhG451VxL0YNcoqOCqww1hHTdfAoBMHAcfHKpp0okPMtOaVZVqV
a0/45kNRsWAa/xgb0/C5AVVD9u6w0DPDdjSmAizDataRJprr8xDFDfab7AL1Gtzqg14OARFrCX8Y
VzRgT7zPV92WN08bNI0So7Kt4U0MzM5cM7qB6ssVCEDuQjAHBwD3e5YzhzFTpIKjsJuRnHECldLP
MMkHIYssMj6/c1zS/BwgjmCojzzGdnTz4GD7kW53jt0yzDCnrM8wqDu2UPkBCfYtH9XKYbt5phSD
nzXhpBIZ/8PMDzr7PZm9+ZtXxQ6PADABq6t5riuugnCxuJGaJBFhxsdlID9zC4RTUJIkJfJcfLnu
kcmvgUGMe7yWsTeCAVmQe2CE6jnHtWNgwa9H2NoJEdOu8v4fT737GtOt0KFUkhCiWkaKHyHFWb24
16Xq+fXzrCP7uaEruJZw0BZPUb9m/M1reX6OwNQeN+9J/xQ//btDVbljNVpbevBtIa3e1mbuerS2
yYP16Qql4ANxJaBVoVjgSyQDf/Vk3etScpenv9B1jE9IizoTMuHp83TdKnKCxv9ONs2ShRkW0lxv
Kwi22k7kyCbUaByS7FQRWsPB8Xyvgbei2wXIW83YfzPu62MKPty+mTfppDgoFHpxzry3xMCnEM17
9Sf6E4SuCYwKsWL21vqWicuoaNGt+kfyXi2DZwttyFNWqsMr0ug30eLM0wfJIrFvpP7Oobmsf163
BVU6kCHvOFtFeabGQM5+1ekXsw9lqAPwZqxP880VhsfVw6W6B+em+Bcw6ZGXe2piKQd5uAdb3O8q
PptadIWkUq6zbrlq7iNA4SuoU0zy7KZthuwv9lPFMbfs101jxyBGFjT79LRezEIwjYWYDepxdwAc
EVNQ6Y91alqpXDtlzVQSeJy3dvnvN9BdgYUnqGX4AMA6a6RikKXrOQgwU1T7bTKsF3Wl9mQ0b6wP
fgrNbECKG41NuX8+WRFZVRJigygXgaCejU6B0/nbBG5xynfz6EY+ttoqYIgHp7GE59T3NgkSG2HL
flPleeYb1ybhBHlEsC/NZASazuLTeAoFg5aD0kXdGZLoqAqed4JiWorpH5oyetuFt6lw7Js47Gvo
BDiRMk+KYr2wdvr2Ius1Jl4yqrMTZqGgWDP8Q8Y9CY9lpVEvY8phjVIHdRAJz5AWc398mzPK57Bi
NBn9RdmV5jjHr3Bz1ouMHlqy+bFrE7Sr1ISqbZZpcgls1F/WuYY3wNURYjynS10c2tw346zPGRXw
9IlOx8EY/P/cV0c79XjzGTvKZyZFiYRdwR5dRXFUmazYWf/RmL5Sp+cB0prBFgoKga84v0XsHLPY
Rf/sweriRK21C1LNSg15tL1zbfp+rpjzhfo2Mbl9SiD+ZwwjiKzjBeRCsSTYt7wCYIIqoaSAcbG8
5/94Zn7mtxYMBM6LIh71zZuU9QLHVMopFC99uN/G9A833Ks58QHE9usJ/UyaF4BJrdj+J/A0DY6w
KKg6N4B+2Y34dvKPHNW/Jw/qsDqGqoCUiiL48TaoBnSCWLfxYTZ2QtnLQc2dQV3C+lCtuZxFL+d3
03Yt0z2X/m4wd53zJ2X+VbklROwRhPtcWobuI6O5ZuZ6u+d6kRKDJg7MlXk+O+6o4SWTwG3iYWtZ
67DgO+jLFXBcyPQsdOHr1WUeZIamA0sFfc1hPLZBw9VRazoxOzzF5omnwDisj8ALtfQ/gmwhLdJW
qYVSqM7RKQ4twtGl6iojjHdbHbof2CcDb8vCtfVS4OTf+OOgYwVqPPdZaQx4A3DODE+1lDFKu4Se
OdHCKx/4SLQgdCEpJY99fVF/8xZhBTqaMzZiET4x08s6qiwO6zBji0ezjku/VHAbjTsEx/wypvDf
iSD4cc2Z3gdT0lTgp0bVZz28ft+6PN2UjviZKLpwfsjvWi4jT71ECnfqwS9Vxbn9cmtX/WuEVDd9
iNqMKe+LPYdVUsmGQEDk1xLEjmB0zvjA0l8bpTQcvDgo6CA+DbKk8VN26r0yGtGaBK98kIMKOoG8
GLOAavN4OyowNuFGhcX2l6sgrdBxThWYiIxTL/GvGyXlr0qD70RaPTnvcuRm56JvUa8DnIdYKdKu
IJoAWB4kBCEtVbGoEfdCbatLGFpRgimDtkQhr+wW8XsuivDZUC63Rk0XSd52hvI1TkAGNq3wMoDx
gGruhI3R3SOAvdsNSV/hmphHjAvLbqjFHxk1EG8euryV2q0VaYDLaa/d/MKmuG0aXzhRzvfxD4jr
Q8Z4vP3dxHd8B9siVjAI9ckze8um8YBeh5q5YbzMwTs8hiRU1NvUs+gPtEkD7+fiVaJZ7zpxqVjw
NOXPLfmuXbbyJnmXvtBPDSbZtQYCVUeh+LxWJVOyK1XiGXdQhYW1GyfjBe7yDR0yoBRs/DEgeaqi
CfzcEFRAd9wFXs0U6bu4HfCPadgd+vjre1UBb2rhGN7vCAOhbPryGbhWTDzfRZXzx9jKwiSx0/sz
qUuvOUTvDiFaqEpeZ5wm62I8J/GRnGnFXapa2Pd4ZcH/DbWGJqMRjGYp3NyYdEXaU8OsRENKXlxk
d2+7Jo5Kqz+Mh+oDHMjdOJT4PrGffo38Tq7wAE4IqE+E4FbAp8vGDHiRs8BLfhM6MfO+BrpvgoBi
x7lgVNc3r1Kn+FnlZkJHMInjxL2Nxw9aPp0A3LfdjmDr+W/clW6m5dvFRA/PTwjDlk/U7On3FwhE
i6TcRPhxo2EiyVz/90PgpG242Wwf8Vta0o9nwI3QSDZd27iMr008tvDw4d/yJQMqKqp3yDv1/Ij5
Xglvvh38Qd2+vpLB4B4hYB55k/Ds+ED3Q3gMqpqt+WHpGZMdT/p7yYvflQW0eAv564V2s4ZlIm4L
HmKXZC2ZL4diHQfks6zhistXHm8tiKfVwYn4D9gW5IeirmCTjPQObvbJ1HjapxOAzkKypFABRk7i
g0/4YaZ7j6BUZKpcg43jjxV8cQWAHFPiKB6zTHO8q/GjgmZK8IJXDOYQ5BaLlxHmkrBnSWRjX4R3
p17CxZHouxJHZnXhMbAUK9T+GCRch+/XdPJV+etJuJyBW+OnnWG4N8rcPfNeJjAxXBpLGUj4Ro5W
sHRfQb9jMgGv0QIvII/3KKg4O+og9QPP5y7169dEGjopvQpnbR6Ut0FdSZSwbm5wXXoXgA7y7+gE
nAOiF3UbpbyFnxcjygvC06t3T/KaFwLtknyR0hFn7/xoQwNMmcU1MTUI03t1kmkdrGR+VoO55CYo
oF6JVg0Sg3UD1SJZzQ1tHRJRyXD+sdO0y9uARQ+5sJfFntwvdbqvgj5NI7lHISFrU96oC2KzFmEn
SDJdkgS62xhIB+f/bdH00BqK+VRakQm/8hEotfgUErgQfcVOsDtxZE8NzNuM//nHrJ4k6T6ML0lW
J5EilNsEZn2/WFzculRpZRjFvC6UBGYtr8zfULyosNIOmX2hhw575bF0k+QQ/5bChjJ6NaHK6GCl
m1aJnCFSc/H9ASxKWLC4BessqYr+vUNQKMHo/uWqRvdoxrYRZd1zi7ClnAjoiwoeujU6RksXEWAr
C88AHSXP5k4UWWtNWDImv0bv6gE7SMowobb0Q4TDiHXAcX/1YXM9xCC/Ex/bvmI/MGdXV4EPe1Z7
4BQ7SzAE0NpiQsOmFJHJwTFSRmFt/+AT3N9ttrrYbq63mYf60Nl3d3I5eARQcxMcYOd4bLuWY2qt
XZ8hhMKx7/veHBDoJpvOaN7fj3UKs2cG433Is4uO/LP2SmznIc0ip1d0iRS6yZTirHhifTe49BPX
8yqVTXt9Nsx7pFaKGr/N1Rl3fKLeMm816RfS/l5sNFnun87/MLmU2oVqdeCLf7ummAy/rNB4sOU5
EZBEi8hb1tPO5FLBBiQ47MF8aHy+3Qfpn0s/aou9Ay+0pVQCRCqZQo0VCkrbqlE2kZU7sNmW6Y2P
5Qai9X3oW3Ek0dmbn8q2GUIRe1Qw6US4crC/f8/Ha6Uvnf8/MDXWFX6/79Vwajsu4iVGvEnNjDg+
Xp8DMT1fpJminprDZ5zGy0nzy/J4IDbUcklgOFimHkd9vPHL+Llh9TP6ou2j+5bgYep8jfOYF1IT
s4VX9cVhLVB3VFrYZHO6Bj9gZh8iLemPfxCC3rA0n92Zj1l5mVovYMll0GukbbWBPqa25lwI//2J
RAQJd34Gup8hy6DTRALb5X++dzinkZNI4fX4Omspm4DCoMq52zZCac+HoZTGrNS4B7/jxA2jmr5t
DZGy9q8YUjCoOX3BUiyQBlW0cxh8ZP9hZAkiwKa7O3ZUQyrGCUHCMqzSiA0Mk7wT0VhltgJh4xSX
ZqTs+6orV9n089Cq51jW88cks4ES+tByi3sMJpFEOARBRB8IBW0tXvstAAJkDLxmI2qrdoqAcJKL
S0zQ6JpOzuuzVmessW8wWVyU+BT07J7nVCiizMp7GTgZc+mBCRxO/8b42wFEYPAsdnO+vb5AP5cM
hSPNGRuXuxSaJtXIz+wJPTzM3MIMfo/qW53sOr1a7bLEt5P/J1dZLZkEwl4KlsREirTOOTv+DmZl
KMJda62PlMAGUIdktaTrLOY+73T4iHvWbxU8qG6/i8xNwHuUacsP7P5YNY2Fri3Fsllcn/cLhDne
7+AjEIFTDrhuh6BQp/203Zb+aLVi1pMKoFWgpSdzOVtex6IP78aUHGarlnPS1VI9jGN3zhkl4yfs
bFsKsPxxSEoWQxco+vjZv1D8YN16uJbxSmod0zVk3zV1rys/CfpnqlKJfqEL1C8tY8+wrKC+bGR9
LMYMoyXOmXCdASF7ssy6xOQJU8YGt4GrZISLKBSN5kQEWTnOcDXuG5IyK58XgywKcFSb76xiI003
jHERXgyWVdP+kThcXDqk7lsiswzB1CmWj4Us8mvUGm/D0vLBG0B0gdcp8+0eg8UccRfJNPbqZQ2y
ZPFSKbZohYHV8ABfGhVDaWjB6z4oLfjwl3BgGvZTRcy5rz2Y3s9tRQiTS3EVVeYtgV6RvRd9PZJD
I+SlyZ0sns4ESzBb/zIofVTApy8792pB1k9fhgc3Ca0ZysDDukLFQ1pxMmlsQNMpJPXx9j37CNfp
tAzziV2T56mi7AsQtc2dNGtiqxcVN/FTx9VuOrhEing63oBeyU8XGrCJQRWi3e+wb4+32ms6bj74
10PWuYth818GJHlGiamT5sISdaUIsoXUyGqbSw8u5k/KDi45Nxsx5wrXNr67K2rmrs0Ggh/KS0h5
51MhfsgvZKojq6g1BLm+4TSZLwNh8beiasGqbXdqjnbH3AYZ+WS8qIMt1hOeBE4tMQK3yygqs+f+
IFSvSmTabrm+hn1UqFHyKN8E1xy5tbsGg0f9CAvkogDS9FoRyiKrcb4G5yVZKvUtDGYUsssgZ7dR
ummF96wBt/qEzFzDdSPrPSj9F8Insg9RskgWT+k3pqBnR/O3/c2w2NySX7OABPbxhWmkLoka+PKA
gdbcF2pk6HSXMr4An3Q59fLxfjyQ0RnkiOh+pQ5K9MVajBY//ncSefP7e0qaBvLKxOXqltI0ZDro
pDfokUpxAJYwDOT9+DGfAlC+5VhFRtdr32pvOcdqDBXYYGnzOv37lPW9BUeZrhuJ7MLq5GSKId3x
w4CCwy9q1vTBlziiaNCadZdvbR3NtKflgraebPU3L3JiooTCi1yMrSgsZzzPxS3JL7PRUmKVnhxD
CdAko0Ok1EC60ywOp+B2PtP2XNdnR2hknC1RHHEREDWPfoUn81u5DewlnkFr+2kC3mlzL1jRYf6X
XtZ5nFRx3251YJ3TBnjrslYTTqVzBe9IIFvCif1cJ8sbBJqHO8cjysiD7ICfDJf95QLzugsF5XY7
x+rCssG2x8VRNfeo50rv6VHhfE5azrewu0OsqVhaLZqJtr1Ya7eqEGwmSaIdwsAYM8P73lC8zOcZ
I6asAcjmvJ4xAByIE2ojQnvfCJ2AnW887O/r+JhBycHJ9KmnLU2r+uhr6DFJ7g4oLxqB4+wIA/bc
qL7vSWuaLzmh7gtx2JAw9A0MPN2hpGj/FGVaojmztl/ZnKMKMqCQR4L6DpZugbXWlcxKifiH+T8L
TUFyZULqFnzgLd7Ry+Lh5N4UWIc8uWflMKp50nOLqV9wIdYaMkUIMzbi63An/UVedscxgGScM7D6
/ECJerOwMo/mRNG46CbSL8L1ZO/USkuPt/FmFnIbzX7/uKYZGdnDoSSaKEEi3ec0H9WcbLngj8Er
8MPUd5fkZPUXdvGSGgG8fvRZB/TzvbIO0EoqO0Cr+wAOiI/B4J+Lj0Is5qpDOyYbun9XJGrentMO
FqRviugSeMqZjpoLv8oYfKqPVMqQC1JLyQmGE07FTms8h7UNau6joEok4lnhb+xVtU0KuOtZgAdU
4s/JpA9EpfAxEmqdVKexkENj6P+221ic79tLCITJsGTkjpPWWlx65pqba+vvD9gmGCx+8BsAKoN6
XnOBbaiZFsS5TyhptJATfEJa/m/COnvnNeRh+Wj9PGll0BI5BRTg45ROUtlociPb0VF3ct7/3f4A
e267IlwV3Y/qKa/50ftHynlQCaI+ZWZV6jt5UqVfOxZtXPWKKTqZQOZRH+eOkU7Ml15v6atBhqP3
cqXnPGsYv60jAepiTY4CdDNwObcST8QAJ9CZzYfG06qxeOhyJAkrGf1AiNLWeOxfu4prZ/ARTots
P+ZegWyDVYef4eu3u4FhNGjNBUXDUCGIOjbLE4rb559/mb6I4wIz7iq+5q4KS6WbtpnJRv/uMBd1
BSKAOwzf+cq0dyGn0DPZXRGHkVK9nBaKjr1LYgS/HMO27h2ht9DUa1bVFYaplq1i7rmgGnlBbToI
jrWbqdEkYhE5WSum1KUiI03jP/QELuAXpWIcJu9Arvog0W9njLJluMbDHTAx55L8S3CXRlQKW7h3
8PQce9ZpBboQDJ3cMpkW6Hv77/mdTnd/dNbBgpF4rdFrDQOmCzwUdAgWILjiZUT7t4NaAwuN+Pxt
xHhK6HXKNgEOuQnrPw88xvIec8t5+RShyjrBQG6dKGmoPMaW+3xmuC7mvwLHZq3LlwnDeG0LpN7V
NbAb7XIfoBIBDxoulkIjR5QuZiL6OcsVeWkiSoF/FyDZiF7NJr0OiBpnX4taW77LAmrkM6nGFl69
pqDb5ujFTWGYUpnVyoxe2SntMuNSKsKz56WiOEQg8I2JxzTaqRhsQvH54qYkJ2tQtmVMeaPqD+WZ
JMHcZS01BFHLRqf3M2cX5hCoMvGhh7+JMa2WWFI6dE2N0ZjEQS1K6It5/dW7ts6PyUl3bwox9KWh
cAtvt+nxWUva5C2qPjG0E91I4KOvtFWQnX1K8AJcW7t9xsKn2vUR0fAStyFjJwDUfY+rU+WXfoBT
I6cDOXI0nrVvH+AljK8xcrbJfnXcFX/njJkxdQ+hGdRWQXz3kwedvOY++N2/N4JOqwGYQHGKX2e6
vd90AF3HTYo4aYd90mkH5dp03/Ti+LC7gS/LF22/LnpVIysV4G4sdNAwpFH+hvTrNhDaZ/TY8F/8
+MBmhQBtmINT7XdoxHR3r/cDpXMkH+ZO75qdF/Yz0f0u33gDuBuinjRaoNRnUVnf+9mJNSH7tcjj
tlY5dWnGHIVNuZmfBeDF0RyRVDuHipTdIqs5TAC9ZLOeJuta4cTm9yxAkymMRMnWdC8dtw4AeOd6
rfPipXRnZ7XM8/V+PRmYjY9/QGbaCjVHRDANlRqUk+v/aFA+SN+q/4Ok9iPQpVCBRj7aBf5CG6OM
nCYL/yYKd8S/y9ZOFSX7xd3u6RY69gOjL1Jpn5g3Y/FU4vj9ynYPkyF20ue5+1Y+W35YJswebyup
WWgiuJOk29fzJ/1lBdsej4rRH0aMoePFYnbAwzoTup2HX2PSXuB+4aExovb2caHxzRSVw235W/wW
6WHSRnUuMP5fjVocfazMZWVYjysfzCCh38q5qA3nTprMQhWiV3QOy0cE/eeGdXFKiMbcwu0kOYcK
OGtx61ZVzVfqpYnDCMw4Ac/ZuNpDbKJeQHb5swwQpOzxFaAnYpe+R5uyLFMVEgc8xBxo21w2IDjT
LXRpXKxFrpAC2MfJyabZ/29/5eE0XKLPtaJLs/2750M7smzeFaV4AnlDYYb6JX+OE9U7VKSQbUtk
vNUPQMBCoCQds4OT7sbJQhQdvkJiGc3IEooutoEjrbLLe5WdngPGr/hMwdi++rkrkv9ikhog2S8f
IQnMiRZUBFe5irS2wEbydEgIvjdNuJKE6i0cESLg7Hd4Nb30uNc9oOuGjM5RwL4uv+Zjpg22Qj/N
pUVnMznlOl7DzULBNRJsyTxrrcwdE5nhPzYhpYImjKCyvABfrEWNruHgesFqVBcGimkbrPgQhuHj
h+/oraIrZpuIXwW0r+Am8ry0uYVrZL5cApBqZTukjieqn4c81rPW+gLpUhEmtWDQasEb5csmaKzv
BwlLWy6TA1JASnTPT9E/vrPrBXRuxVuLnyxYnVtOJf6fe0LtS2/wirVprVdzHFEYnG0iudNzKzfW
nWv803ONuefVOwyUzRpn341BW1BpSdv04uUyI3q40ghGRB33YF8LVXPTBlKqIFB1Q6sX3B7VBQYU
yfy2G1nni2t3atbib9R0wHoQK8qCxicKaBnF6wzESd0S8+nGFJJSlc/MugnBsxJB3L0kU+zRtJC2
aW4SZmUtVYy7Cb95yUgr9KkmesjYq7s84nQogIAL5Y2UMHu7TptukzWE81OMSdmiZFUvPW7bzT+j
38vQQijQC4MUE0bmOhoZzoAXDQGhY0B4HOpYXGgG27VWpCGZ7DpxewZlhYGcUJozARHlxMI2bOiy
lEqAXqVyLdaAFq/HljJYqNjr5yzg6h+xMs61Ulg0cvWSIayIo/4nrSL2fTJI544ATmUhmpDXKRbn
rJei3LQAIRrRzBQayXswV0e1JWtiYzQ8LXQBk/aTwu3MXChUlkaKLIy/CwooT25ShT25gT/MamMB
jb9MgdOUj8RmLLVXAzyQ3LQZr6wMtFrY5a4Wowayl/iWf13vxIOePdVX1u7YsqvGwYV19VnNZY65
/MQT6q549DqBSWpm+akoMowtqCz4avSoBuCkd/xNJlRlfL/fRpPC570NFNJlCbLl10kXQBdS/Q+x
GVlK6Tj8LnC8mR0jS5CVSYC+LZR2ghmECYSQbOXIb5HXrhk0nhwH/h2yD/j/KClYVPExO+VJnO7b
HhuR6nHm37VMDbkK14NQAx1eM23v1VoZgWnf4D5+sybeNfdkuZaOwnxZWLoazG+cdevGp2Iwec4d
fhPLFOZ15fqMXXlmfwvov/ZooUEG4cOG8Enqpm45+Upg6rJSbp84S+aUEOAESGXNAyDax2qw/bdg
BsKiA6SziUE10/A/kaTiFr4hTymltD5m8c9gsLFI6+Sdfl4FtBj3xPVVd+6FiWtx06Yck3c+Y0J4
IIHoImQjG3RqFg2zaxAxknj9wFCMCILHt8VCoBrx8gZ1Iauexjrfw7JEnd8CIHPiAm2sGElEv6dw
xq3VeqXHRQ9EE+ZRT6vEyfUC5ddnC8PXNYT42bcCfqniH5MSTzPqFIegVLyIJXeRzmt7K5QeKFXG
nx4zrNVyjLSOTpwdMKWL64WaljEjaOOoIm+nRv8S4oMZjmwgSiaL0ZgumxIGpLetZ6f3VF5ByxIT
/H1o9rLqA5GYtQMeTrrXrZg96gZ2UgHogrK5F//yy2K/NZlX6bFWXvapZpH8eG7oF1amdVbtTL3n
YgcdG07uflTNRT/0VZaxSuKgEWbY1HpUHaBan+5k6dAyK/GpDu+3MJkF52zoAO+9Svc4s2qx1TP3
jinH2YPBkArAyX2GN2VBgJAyKSIYKw3dEoufRdrhjpdd8E5gZVZSRhHfKSWrsIfmajQO0lpdEC46
d/uK4/Udk0xUU0y+5mogY8kcPfypCMPkU188szEPj/TWioBoAAn+Te6EeQNw2IjB0jgwyFJnf2GS
dPyP3Dz2jHPNXhF5A/v5K/rAsKXU4FYxRBO9CbDZD5ayLXbfPhRMPiSMPrwUH7V2PxJlWgWgiW8k
oyQ9Xlfg+uNCClPKZ+38VShhmzL+f0mwdgJriwHt+OWoW71RNAdhSrTJa4rUhNiYHRhE1hqrhaNc
9DXckO9z/SyI0xDgNFC5H2JTOCjcRbWy1+7YW0QTX+JKK39xSfMmwbGk/IwOMXajELvsfoFZ8HJ5
6nnTM5Nr6/zcCaEN/Nj60c3PArzqwf90LOMy0+nKlrL9bR3GIA24e6vQze+5PA2Bh3onV8Foijr2
JYr8XkfzUVfOdqEzRnnooXzIUAL+lcIIjnpmD0kHHR8jKDxsoBrKIjTPdsmm/pXaLGCszbCFms8L
/NaqGjGs4g5o9/mK76b3PUP0Ahg+vFoiPq3dFZ69M6GGcdvKHS4Lch9IxphSGOjUgnh0JJyxh1ya
lu2isUQ6944JwBqi9ubPF821TDcTlITUvu3SOKEkYnkCqoqIj/dFrgJ29Rh6d54L7YcOaOCeQynu
/es5Xe++I0n+jqMjZy9RrwbCjUhU0KPfj1FbOHmnEO9ggSyWm5pXiRxHNpGXd50jjmrjLF0FSntB
USLYJT0T66Z7Qp/AmM5lHJD6ehUFbFV0Fuy/2y+42Fgu+Or6Fshx1x0k+ZYcarCUEnkFMxziCkVo
afBLO763TnS1/ZhOmmWJziIrjFZBSgCVRJi9F5VujxA5w+1LqZv2SlUYCwV6nMZR9zhYc/F9pmxo
Pt6ILqoITSSWHpCLfzR9MQGXg14XtSj7EUyY1yOLJI6pWCapeaaJFrTf4n/FjSantRPZxyx5HA0c
rM+KqN94NyDMELv+hU4auoHulEpKbop0CsZcqLah+f/4YM5nz3OMoyT1LpWeBpe395NGGk5DuJY2
w6/7xom8xajvx/B1zrobmiXrvAl59pShx93pBFzRaQbGzpze4Z9TTP9iKfpHFTWRa+vm2nDvE5ut
PemgkPYIwAUBiTYhcXX6OOLFsxFHtTBwkjg4Jixjevhhiar6y9NdlDq7kqpe3F/0W02a07FzdhJL
/by/uHyBS1JQU1w1F1Y08jIUSDZJB2CJay8tTgsZOscm/os9YgIzw1zSckhOfdgypFABadHyeyre
+iku3k+J44Mwgrt/AtX44vrtaaEJ50YBW3rykbCPFsisUL4GndELQqn96+G01BDT32MMdewi99ma
hkkV/14n97FivAD3LWc1JBlPHPuArXDM3KotNBd3wws8m+NPyU83ZuvUoYOGhzSF48jtfibQpBtK
lA4PC7NdeWDVl4Xz5sYRukCpd7szWKioeCf8jGxuok1pXx8xS2WIqx2kyTVNEyW5rAl82Qnac/aD
p5I+RTH+vUmrq08lQgP7dhoIuAr0W/R6tHh/i3BkeMQ5JlMJEm9qeEUKW4PxwcH8xc+wZXreS/Ps
S1nSIDVam0YHy0auYDCYDPpW5Q7MMOWycay0Bk+QLYJ6URAlpV8qHyrcKIorBqCYHDRxU5exMoBz
iPr9SONtvlouuSv4c3btRSk8M8v5ZLDYGMN3s5uXASo0mgbRskPeYAON1hOXL+x0h5JIpAd6Rbta
+0X6DZCFKVcRvMHlegb2oS2i7pX/hNNhWjms+tIrzes0pngEhfUcF5v27V6VpCL+UtpmM91rShZB
J0XvIeXi0XwqLAEy7K1eugbjuhxrOIFaxZQiLMx+tq+4OuP9gQ3moszAUG4S9H1Uk0YGOCquO90W
POXXjyLkAcT/PqnoGnKbdo3JJfWL0HWn3v7DH8ewGAt5XS4rCEL3vn2ojOWCqs5yaeZcbxsJ70C7
RG/J3jphDGVV4EGlReP0X8RUsbHo5D1nTr9cbwJLBUgHA5/PBsZbOfwUCa8WUDtDqtqz4aXn4L60
dq08fb9T7Mbv7udVgANqKae8whDnLpTSWg0+hbUk86E+oBDlHra2VmUheCn9PAuwuvbwJoG9Up1r
V0bgxwd6KglnNYKjnC3NmymvwDXOhOGu4SgOzy5K+DFcYbw1S/sJUJC/0INFQcwOMEmVyQIrcaha
7o6qWEGgdYiAuInR/XYf9WLh4H/CtzGc+09qH7MkpBYJUtSOwZ3h6P/15fjgLqR7tMBABz7CysAb
dk5+B9jggofPYQu1ylSv7GquByPyvF2jb1Hm/7iTkjAacrw12CqinklTGxDDwOWGUDwVii9BoZ27
81JUmQRqNd/FSCkq40PRHmttMY70enmIFz77Rnn7zZ6IR5urdQNnb8FqTplgFDpQ0zh13gBG5n4X
WBjB+JP7DPOBr9DREYh09/3DskO2wyogH3NM/oWqffzVwbOnYoHYoUNA8gwG2PgaBQ8GGgU/W0cD
UhefwCvcS7uF1e5WxvU8hry3Xa9UImleR5qW+3U0qXroRyeQ0Ir8tD84AsSFSWeposgT+BFpDsgc
tdGrA26GDh8FNF372cPN5rBHJGnjeBq2WzoMWYnUFlF0s1MwDehjmV/jdMDueooPC4NQL9jmHLN1
7rZsvfc4wTxMGG5REO+vKNwkYMHUa/esGQQgqcCfcsYq+YdlpsUw1ed3syPIJ7e1e9IFr7phAYOU
bQrPg/FFyoJNKzaPSjmO35qiCSe2p+QjqPQ5srDp0mU+oerA6LUsj8zmxgmPTihovHhbaZlwIeh2
iV49FV028NX6eVDU77TNE4QnR+Wv1KwSjIM5Fj67ejkDRNJiqYLrGpWnmoYIYWA9bbUjGxbqWlSw
5mJwsBwjDby4UaJY7pLFNzLqD9LSk6hDMh43kg9zt5Q1KcwgeqnQChP3ahMzNc9Enqk5t5rdN6+L
+q5xedxoTRKOVJwiddLFOPvr7PHAtuwXuUWz1lhvxPuTfenQNDfZF4vWGM3WTA9jxvFjgaKKaeRo
JPPVgaDUDZb/wqR1xqdkbF199753xc/das0bIZlizZYmfTsIUR6q78jD4yI+s0B7Lz6kVmDpwZ1q
9heIcP856IfsKc6B8Y7TZkEH0CWLm4hQJgbZqSr4Kcxm27iqhYyqzuFe/nsPEtGdaFiTm1K1KDdF
tYNL0Ol7WYgEmelcdh6dgJwKQreCRcAh8rySSo9RvU17FiWBHhUfJRoRHcmxDLL1XTeaiQl0i3w+
PFbQ+kXYTuNRogulyifixA0kGGhvfs7/4MbfNbPM3uwP1Z01hqAfu2tqd3HvUnQp6vusGFRnZgb5
t+DkdrwIbZ+bpXb3PsO/IeIvzMept8CjDfEI1tbU7WW7ISfbD/9uYNMmQSkrKXqa1I/K+4692zxi
0l0eAGkqKTPVaBijqpDqcqVQs3TdW/fVvA+STelKTJts4vYjEYhz2/b6lGZrXkzXqcxYE0JMIglK
eQUm3V3BnOH/tKod5yCd/cgPJIHbhUQ/yDvWhjR3Dbtvk+r6gfBSrvebiD6jmsCFSzmkdSNlirMG
d7z4+K+KA4UwTX7CU7z8KgUAYLmriwYiqHLYEgkEi77ie/uoIFixTxUKh4xmHA7WXWlqLMv/FV+G
h+nTkxfjbRtZq7WxIsU0gja3ESa8xAVgIYspugoWokK14UGpmp1fP3cdUEgKIOlBv68xsrrccipi
XZAyLiawFBFZWAo7lmG9SNQU9htSpcJc/hir0oo0F8RiyPVCl4unhcJMGueuZuVH0M131T7Fg6H6
dp2XM9nkuZcUEtHq0rHREXz2K8POm694wfoMzpaEwn+h6KmbhbNe1QNtVrU3D5a3SjtNJNCO+GUc
2eCEjHGeSKoN/8mLqbU9R1ECo4+I8eJde4o+AOhpg6GBYvAWFjKU+Gd8w4nLpjl9aFX/367FdT5V
pwyoSV7QMOz5UXwJ4nXHFJHrAGgDVxFRJFrQ+5y86cEhJzvK1qCupa6pRJRhAJXZoSx8WQ4G0KuT
Fx/JMLmhhRcoErU0tmAlgQW4vRHEeHw4G4Gj0JJ2LA7MuCOity1vQFvrL6UiS+8U64YUc0Hxhan3
/PMe64I+BJ/g1/X3iauRgXi+YNPMvP1pqlBKpaSGicbJvZh7dekPGLmImhKFhWgwI6PzHweYRdxd
ncA1jnHwrAm0fg1Vlri+vUNVQ4KhAKuzvOOwSCetQQF/0Z8VfFZ7rjxv+7Fj1+1rRUB4cembAh7E
R/mTxGRd62pmSZ58vYLFEi/2tqIjiSYt+SluvhbVVgll5VGgvLYJwQr+Do4rQXcHomV9AHZI9avv
x5GCKKKGsg2VrSJq4ZHqDq6Q6tpfn685kx+9DJ9ryUdp6mU+ZbcyB2W/a5rGmYwnn09IBPPw6ZCn
8BEiHfxBpDGwhxUZal6OjZgWJKxmHlNJa6437dRYYbFb3y/ELWlENkIozyDPZpiWZVyHf8FkLT6d
HuI35gpY/cyurHKpDC+zTM7JInU155zlyl26Apz6PBpmw2BtlDqYYIcRQHxmbhXJEAc+NUe1+3qV
UZd4CLOQyCYS+H2NZZMhd3M9tIqTeZ807gZSc6CDfCwXGLNlmrJarM7r7LYZElJ2tWbWfsV4ArKF
bXcrdchrHm5tT+/9rD73iAilhnaQOwdXWLDhpXVyc8083knxMwkJsYRbC8Nvl+GoNzoj58pej6sq
Cgrw6OC7TPpn6XSasVcqO8JLm5GTuz5t/RlYWr7BgxKIIqIRj6oBrA8+xioqy8DIyTJPEnmWDQrj
zoP6D7YWj8heXwjMxmxxj2jYQ5rCxsIF8fyfDGpJjdH5GkkA0aQZZO5bY2ulG9Lu//BOiYZjBKgm
QopBRlZ8aJ799P9gyVyKmXzemVkLl8E3ITaC3UHFtcHlfpOtqSP8A9gERlEOq0fAsNjNP2BDBOLt
+ClYKQO0FUj/+naAjBr0BBGi2Fqh7bpQKdCnLdYDrpbMbvNpcXpwXDtgmPkK14uV/0DHZhDtg6V/
mg/4gXjbDpD7ZcB+E+GB3wjbCi+S5NY6Ga0wD+XFcQD/1oDtd9t+k8Nwh5OQVF0NupDtXWJEh8A7
qyvBFLhTNfm0i5dL9C+i8y1NlDOmWELF3yCL1ruc+MBECf6AwU/CbeLpahBemiFy2j1LKYuzhHRW
AGZGZ+01wCAEqO1yKMQ7/vqqBzFzlwq7HnUBF40Hbonn/616Gptmx/+EHS5x31nPhZ7XzOjm8sc2
Aj1A2ms19+G799T3Nv0zqPv00hk9Kkrxto/qHSoQwzURY660F6doHPz1VuFsD3dDG0jn+s2Ii6mB
lMGE9h174h38aivtdCYjIBf3UrOhGZe/FBIHnC630HnCDz/Joh3GHjqi1MxRyP/p7CMMYAXwPV7l
y868doTM4Xai2G6G1rWxyZ1ynvUt9I42hsEee8OI+QbikIgoaZAqu/yac24qzQVTrFRGAQItTStS
4TH4KdvxVZxjg8TOY5yF79TSCJqfIX4LC10UJzBBWvVyxh2E9Tr0y6bzFgov209xDsfx3+Blapdh
zjsbhLkfVK6QIh8GWebCpNeLDKBnOXkoTP5Djo6E/9A7HNUt3xLRvfbZTf7j2MrE5NGfiIePROyz
Gv6U29umcHO/dZpGxEBwuj5n0kQTgnlH8/vRxIeV/htZc0um2eSBR6XvOIFqQNIR5EHPyjPBdLEh
LgxB9NQ3sM2AXBoIooDtJUPoYRqNoAr7ol+HvGAL5Xri+PNiXU56+F9/cecxz3x5d08hRWVdkvHN
TKyAwF23lN1Rxe843iuCqbwy5C7Nmuih5DxMXP98AsjBvsM1v+LBQZTSJlyhl0LxVujMfIXmlEZp
rPXUlo70oX4PFpQBBnPIXMJbZojjhDuNrXpBP7BMYpwqxtOsyamZoB58311d2movypiNlZs5xOyB
ZjNbytYpUqZY+09938zNtVl6k8hZywKRrZa2yNYS0FfRnnRHqxQcVp2DSoKBYGBefNz3zy8Y0Jv4
3p3khux4qHzrduK2ARPuX2R7umK4/YIKvbBr09eaizupCk2jQwNjbWowcHdHAepyJewt83Cxwbfa
zdam6IUxfcXsqYpVsxPlJHyo2kRQvWHYQYp6Dys0A4AWCjaz1npAS8a6g/MRqQW1TozIGjT+Ifv2
UpYjXb7+1h0Ek+2eRv+DC/Jr42OzwNetpi6JJdR4yWyx6VQceY4AxRPyhCYekYdXZ7fcQSwB79y8
pitycH3myR/f0X5KqOg3nOcvcw1DKpZAsWd7qX1t93JZKPycuqOfUGXLbHu2vPSqZPItJjixA7lY
aLirRRPkALP6wNMC7LCVMn8OtHM2FkSqUyKnNgfyZpDXvXwKiRGRVrku+K9A/MzQ2fZ5f3oUTLMf
pNRjxvJac1b3b8cClwiM4kjNHrhQ+KHY5L/UP5dTd7qeVeU8lhP7dtvkXUTMwPdYBiEvxeWpcWEc
D8/Zd8aX8pIg7fgUL5VclnrP3DKRyrLN0cKa/a04Oh1o1QNIYXR6ONzGvclQSOCjC0pnxbp3wN95
IWuGIlvKhgcwyOvZhTq9JPRYYGN3se4VsoUb/XQPM/OSCqZM5KICaMtiPG3BsBl57fRVKADTKrc7
RddoUdaLClgE2TjDJ6SQVDlYwksJoqAExtAYYpZOxCjqmRjdGPbdHlnaKBmCHCYtReK3EYVn+5j6
Uvh0wmKrNsmRkfCxhlEiQ40tHj9hvwUpoUc2qibbh0UPelD0/+dg+tLBhlUKP+M0jt6d2JsPkMBf
vBJsKaRYwBZ/g6GHfsg+PVp5oQzy79gPs01mcDhcL+fO5zoviDU2AscojP2c2kKG5yczBfy2wIau
G564HwBi8Q99QFkI9a36lc6OPbc2lkwknW/gocmEUMFPYb5B2PEZdJntrumueOF9HWYyGJ3GvcL8
ZEgW34oTW9f572wnYNs4BM4DghO8QDc8/xd/EvZ+UZ4666H+OEcBqfzt4ji7ZKZdwyebePHfFc9B
dUBFGLd0Gs17XaP0TRNgf105Qdqrd3KfHpn5OdLmYkiXdoxL8Swqrcj0/xeuzuQlDaG5S2exHTec
d/KIIYnGg4wpgnmbQAMeAVoLq92u8ViEBFx3BydIJobSBdVhThAtSEa7sFav8QOlPAqrsOWLiM3u
QLkU2tiKnaRvIjNzw3+HbhBupsiDBCeRWJf5HJt+XZz9QaMGavWNQpcLDurHYQk08pbWILdMGCO2
x7yg6QlHrowgguLLNndhH27rMPYx1QQ3aIrqWYokGlErzfBa2LcqliA3gAN0JlyAv0boLPy/YSKq
wgCjrHMIyKvDHsRbUabaW6Ra4M6rO5dQHUY1WkmKF8brRc5ojimSvEis/TQ6QeHUl1J7Pbg0pYKM
2XY1+o7qOMWtOuYJVk+ZptvX4vUs+/IRfRJKwV6saBSK2Uc7lfT+nJNHsza8USQWBeIG+TyDcYwL
tXoB7PtgHwgPDIzWmhgScqcEcjOAzGDeiQuskNUtQBbtY7AnQQ3FkDQg9LgCkVZ6Ru/UdFyYNI5h
ILVBuPCzt0YyIHQANiKTDWXP3gPbTpJ319eLWm3jilD/1bs86wAon2hf6qrufQaYZaz7qvxhgeJV
PygkPEE5JUq6YOqWj3r5ylr/BleLmYz8Fl94zNxxVWY/a93T+4a3D4RPN0oU/qpqhvIlfjGTXxxE
FkChmggCs54R1DUYbhcGHj7UDmi19xZJrDurWqJsbbfTnuqqLv5ySsxPVVEha4vkLEhekY7Db53d
bt9xhRJ/Lp2vFF8aIwk4hUXY2AepxRkuQElNgkDJERZYGmjK9Ermc+QNeW+zOmOX1Qcz0lq5GQPO
hNNkHjzqExui0M8RKoUTnjkbjVnNHJNOdE39MarBZvR6HeoDbYQPPG+I/wm4rQtWoRaKccuzZehm
hH7DufLHU49JltE3U+Yr84MDsoDoRdIGDHiqHHTxthG7Rg4lvFpXUOSm83TW6P3FCTdtHfqRk/LM
LDM7Utmqtd6XS4JILNWTQBdpeLrLMyOIrim/QqhyYbSnVmM7bgqxWNMUrfs509HaDB9QWgFVP9qy
lpq2HLHJy8qaMJNguM5LbwQ7sFzp8CUNVZxfYl4JTQPXx/JDCu2nJqWV9yFlv7zdxNCmSEzBKaJr
Md4nu3aP9Z5eYbelyOLc3l7tgfieWHTk6cs/LdDli7Nm+QdDGqpsxYPiyd4qUYB0LsJAkyn5PRU8
rH8M/jxkgfjWQNyNKUmJmVWEN1DbtRaj+cpFqoGTba7veFQFx5jDHq463B54yKnTDRuRUFX/bZTs
OgUWmJB0xRiFl+tGoCa2Nym1Mr/sw4Y63DT94hyCXaibQEf03rcKOplxTMruBESpC3vIEfhRHLdz
SdBlO41sHxmHabbsDWwtdq6/deye7IP59uFhxciyuVU7G58x+nO1GU3hUZlDzY6K5EIvOMJ19dov
xQ8/O25XY/Q9JSRbe+8tqwMO4aUck9YhSNHaLmeipz1JjQVMoDVrlcDGGRXLAMx95zc1gxT+aJ/l
vB4WNFy8HSI1odEShJS4E5wSYxQapoXJiUK8g7kExNKQ11VB6nzfbwb+zTSRltaL8HiRm6kM9AZw
RMj95wWvsVSrPt5xKPbJuCBUl72UIdsfiwFYUSFixyVF8FoApqRFp54iy/KoNaCS7E1M+zJW8zMQ
6tGRON9l0cYVtGMDjrIhCosWr5x98L5agWGyntI5uiiAvMc3fpfxCsoZeTtUFRHeaVy4a0wqHN3z
SQvOYoK3p1U8dsh9B0DRpchMW5RqTrKZ168AkNAddfQnrFus7Pg55VsbfHDyYKPj2JS2AhH1c7Bv
g3gs2Usb0BYvt4UW063jR3vZfFXm7C2ivBS7Q8nUortUX1a+qHdNoPPBw+aBsZ+SVAI8DqLTtMVm
b67F56gSvCywQjbCFU4gUSbfzPhIIg5UzzV+VihVu0oAfEg2qz4PzYL8ysrcFQ9qY4xRpToZWC5T
hzscyNn1/JQTd7U5r2LSBnom2gfksoeOKz7fRoaPNWz/6Cfgcrhvl1kOsCEH36yYvu0DSl+URTGJ
j/Hha/c0kFv0LPpSkNLR/GphFaPDCsg2c8zQjy1Vv1lUGw7PmncoZyXusu9rBCVHe1GXTWOuHJ/t
ahNKt20WYkSYVGPFuxx98kck5B6snt3kp+GzDEe8u37SVAhLA03BUIV9fAMP9RLvVRYYgl4WLwE+
3vnxAVbHBZ0CG6k98XKc4CSInDNYij/oVDnG3JNvtn2diCD497MnkhAOzWU5qvD6CkKV5cAuhvtH
kd25oFuYoz3hEe+0VhYrY4W1QBclH+tCXHy0lgziMrJGSonmbR2HDJNiIu0R1onhZZ0BoG0OZtGi
3DYT7EvyRScN+YbKolTnRTo7IH7tq5jVH8S/WhcclqKkPmpm4ZGkt3U3K+bzmv7Y509WiSTyDNDy
4BgEPIAoZuPcnTIxvZVSoDIS5OD6+J/MtNYey5PO6cyXe1NUcHJ+r5saoZGdO2Z0C+HVHNTR0dKh
/UlkTl38SygmLTGnQFjB0BEz/v3iZ30E/fVetSydGfvHNpuAVTJA6KKDzfd7PF67UFtE/GtkCUFj
oNnlCiBKlo9jEIatffv8S+i84ai/Qv6ZWKtMSdnITsXtfeFXUgp5akGrXf9+Q4TvstzbA7p/oA6+
aJEXiTeoCqS3KKYxkQBDTAaSmr51/iq9KkEmaENbH0sdhNkgKp1gcAfgbAu+N60JH3/woq0IHbjF
wAMkuymhkpDfmPfdKQW1uTETUT3c6XWe1iYtPP8Z4jn6fvin9DouZx3lVS30LapSK5O6z5R2B0M4
hQeGuwbhPoFo4RtdPkKpk0IIwbSaPZBdmO1UOAgTQWiKxjTK7wfWmOJJkwt2NR6J+lPAANE3VqEW
S5xgGpN7paterQX9iJORqpTw9s7OS7ifHPdeaPHAnQiovTq9TTBLxOsjUqG/IxbMNU0aqHq18lIO
JUYiEbXXFQIsT34rhCWVm1i/NW9x9KYnnIhey4h9SS3Fg4DW1O2FeYbFUJlqFVi13S+BzUlFepyq
rklhQLCL1vM3nemuwNjhMeDzLbk3miln18bULxGc+HfeLdeFPOh6SXSLa1/MGK9Se2cefLq9VS7u
mcYfAn8PXBSmasKEit7dmva+uV0US2jG6x8p7vgkVCGGjqzdW1soUZmVoB0/x3ZIP9bUqNWk/aUq
bFuHC1TbHMWNP71jloG3sdtCmq4m3jL+VxGwsr1TNkwyYvn/hMV8y9rCI2TAbYQXRfiSWxhuW37e
3Vu20wCGa8aEzoYAwUvLUbBLuZnY6oRSHkvNNR72QL5XNKapKi79t5L1yTVfiDRS5mxBbDD/S+TI
py+0XACTpNu55mYKskKGxJajtL+ITHbbeDbcI1gJt1B6HHyf0Mp7U92BUvbxjzm1dLfHsaZSH6M7
1yTxkf51s7lo7rMgC2dC9SMcD4okLOCF+0yrhVgeKYpLhVad9elv9McCRQLvUO879B29ckv/aQ74
jwP6/lNB5Uk0VfgY6JTLdPld1Gp4g7eFzxCFIQifOE6o3rXe3Lo8xBZc0+ag9i+B8rByg2QZGbvf
R7j8zLBxs0YhsYUsR4ixCbnuH4GMKjdvf9A/ikXaq8Sbq8QcO41BpmbaT4+Bwf47YBEMTfTBNn0B
SWAkyRKoF9Up1R627BIkLoBlb3BESb9eNep+/OAGHa9C7FVmIUjzs/o6+h5F4eXFAPFnCCak+jhx
VW/kfyP4P14KFUutmervXXFewxBHC1lpGHuNePNcD9t6ecs2iOdy9c44+nMZ3+u4vDOYj3BKDd/S
R20/FhIHwmgAD3PPXaYSWWSzkg8qVJ/GvJuDWfX3LI89V3EyJXAztJVmPP5MygF3mSDKNmTNMKrK
WrSUtCf98tC3Sc+xO6FLMS6C8w4Rtyo+2mNcjzNf+WYju+3qQQFRKBCTCp98+m374b64x4hkiCeK
JXFOFo8LVhMB6L06buklRZrdNsaiyZKYYvGFNWMiKRns7j7slhvFo7xKnjvqP0Pzvu9/QnfUWoSc
p6HRIXfbxch/I/+gHyN8dMaHOrZdbKQJT60Lx2VEdr5+9Jzx1H2PxX4X5CIBXsI4icIejxMl+hNN
Hnx4cuuhYfcYXLJ/1cY3T9d9SHtQx0SSqX1u0uTi2zgWLitsZyiGZi3uq6Ff/9/od6Mj6vuzzPq0
BTjfoZ3Vqs7SLQBcJImcXbdWQE+jxMlikBxNphOuo6XEwql4m9puHF1OEaRSU9AagnT84Elxu5MM
p9tqqui5wE3UNfc9iqkwbbiZAbMBrQkmZ2iTHE+E2exm6WVgInrHCt6RHAAPOA+02mRkZtqOnAHf
dCfvHuL9ZhoDl/8U2v8M0GWg3CTxHeiJLfsmLSVCUGlSMSxIv05e0zpKLSMEaZZAru6mJzdqIkOl
L+iIECBJ6bwhEQ3jljIB4Qsclx5Dd3tdQk3zkgQoAo9WPt6wnu4a8hGoUO0Tn2Xd8Mh+hdQsh3sP
7RUNePR6k60XGKhi9aeqLE/ru1g24oetAtnWdjRSHP5oEYgnqXx24HKmyX/4swsVCHQhHSjz9i1z
Z3wnE/6KbS6BAlGi0qi7cVvvYdYApC6Wd8mu5TqvQiSTUrv15RW0kGBMuMl0jLlT5q8iQf3/h4b6
+7j2PM6o7IuQ8i+sLi9KbQ7WN7Bnyf+rNjB4lU5kqabKTub2lSLWZAU+6x0oYS5aeV/QSkxST/49
FuSAAqeRFaRgB8lx/sVsupxJRMJ/XLUYjQnlQkRsmLXSg9P3r/ozgLYllTf4R3E0zLjD09DVb7kD
HAkmtSg0GPr2hElFvdZQXSwsKvSJbZsLUWU0SyrPysJ5wujcRnJK16FujsT0kTvletHprkgP1BND
wnNG5TZKOhAmW0PDviKsHKT7WgU922dMTbGkmHKoheXZsum8CqPO4bbAW98HDQwN1hJGLS6rvZJP
V3wvuv10/ovjGGrgr845SwND4HGPRd2YRS9ckKI5nhako7V5M1SJvMennmhvNfb4fS2RTERfxyLD
jAWl429QMc3ZzjBq22v99XW2paHfaFgPbllXC6SXUs2XyipA2lNAXgjzWiccN2p2rMM2nIWXmDDa
Wj9cdHhkbPKfFuERJx+ORCCkW8mnKfWoTTQ2hhbGrBPoxHg0bryFqt1cEkHycZ4ieOk+b4Vn8bvX
5ogvHTkm09TsUn8aAgAmZvf7f86LlzJBcWBqgifA2HUq/K2Ta2h/cYC4rPRZpEZVrIw48i3xeoHr
VenByMztFQ66rGtKo+fenyswoKVYeCr1gGV3clwYpdqHYAY2j4zpYm/618KNOBBpr6UYyqBOsSCZ
SiZYWqdWxFOfYhrkr51d23VEOTrdniC9qJRx3aahwmaOJYwg8K1LGg+lyq7r2jH0IDXER1+lE4Wb
qxMonjZkfygrmK9sNMd27NSOkx1aLYnTfVFkZLn4AIjCwsd5F9ZzBDuxRFZzBEjo97sNoeGe22bs
baY2glpnZsk5SIl+LETdwy1XMRuCmn5+HMoFdSAXaxioSpqBPKnqxPHzXn7zKlTTS2dRwn71wbYe
DLfYO4/b0aNy0QTl8reb3/bYYq1WkwSO/SnAOZVo7cRHcbkRM+AtS8MO848WRDqIWtBk92LPrwLs
G7Qyn22QNr20hyuSWPflDm8PTsKjLE5uOytyVKmW0lOy6IvWR5xRCiOa2JWwFO2Hypm7WMtk+99p
R6n+nJ4l6a8OvbVFKWM4COrSinfFwBiqXOpiY4W7x80iI7zGaTRf12Xx3keYynVij8yUVjFaaZg4
1eHN4D5FE7xBFK+Ve5DZVE7l6jyPtKpe6CrDseABYpfc4/pBZLy1va04OEvoKR5Do5lyDYeP4Yfq
g6+yuhdCQeMPa3QD87NNk85cF7VwMbI5vmp5G/yzmsTQnXqKA5TB9FA27HXiXbD+lI0ybX+RuXEp
RJofA5yk3fws3cIuIU1Zl71qdsLr0/SWsg0lTCxOFcRP5uR1Nz58NAUvKfw4v4sGylRY6qIrOPm9
u2FgXu76ECiJ+PPgud33/ir8SMybZfPe0xfGujDa61rfMVMp9uByC8WMyV1hktmjxAq4oWzc8MNw
px/AYMlH8UFDd+d8IB/a09V6XvZDFHhH2vCZnQsCCcwvKFAScuKdfgVMfRPoSnt3mQ9AP9eEPmPH
YtazwOpfm+b9KR1IX9NV1EMlO8DG8429mAPta7DY5VOV+My6AqT+8smE70OC+hAbvb39qIyRd3yA
4By1NXhSlptD37eKLvG2BI8HjN5Teve5NL7q3c1RwIsmGSTYa/J6gN6k4icuizfduB+ZtDaatU7G
BH8p+OnY2XBdiL+UFJwRFanMl139xSfqpki8sV2/KGT99hlgdliSHyFr1es6Oug/mfoOd8LFKnDG
hqGNuDs6mQcvWJD+skp2366mRXRRSvykNgnn93VU7vWVc2L+AxlKhuQsIVNk71c6YtHOtlgMenU4
ZUpu3oEbnhr/AyxvDXzUFrmdWMn4zgCSxDA297OnArAAHNsTqFdfGhmmb5s+OGHzFx5XGGcayHIO
tyZuHi4naLlv+yaELs8WgCJKy+rGEsXDQHAYYVQqwiO8iVB5X8S6a1GbHbfqIVMlCUpKotFjDAGQ
J6THu2H1e1TFjMoFluh6L+2vq8XuFHTD8ZQQtcDonMINiDrwqMs+P4IvWauv9hqh2xPO1mmHcOmn
q5PDgfO63Fe4U0f4c14v1q2B2U2pR8zicMakws3zMnjptizNwhlB7eb+cjQHPibU1r9BCdcUOzym
O/vgeS1TrehN2TY5Tv8LUAJ35YTTN4j7FjZ/wBF4XUXSAdKFNAa8t57HAgNKSV3pEFJgEgDt0sSP
CvJnEsAsLMCBWn3XKojR8+o0zIvXtffMo/kR6pLdCcWnXvDe8tBf1gG7+VzZZW5iHfw7OGSH/dNv
jOJB3ype0SLjSpuY7A67TGDqeTMMQbFvC5QlMiIB4fwICpa8/VR2+3rLA5EXX2XNI+kN9QlhIw4I
66cXs3xTKvvot2qoW7I0p5Vx43mX6tfJg5z9KUZqj82qAO9i0y8tVLixbQFkb2k+bQIARotBqaJp
lx/g/qAEdwHy7NJ6uE2xV+vBkRuK4Q1aIhjLrgjLT3XK1Hg8565eQEiTdVux5l1ejmI4bbNlR0k2
50vqZ/dYIj+lFysjUEGRD8tqSeUA9+kVXgHQ/mVI8fzGKjjFNShxp4jPLCdeo58UwIC/RKJhnRFD
sGt0q62P1WpzMKd7QBWCGzeuGwYDjfwffjL3ZBIDGkl8NRhuwaFdHQRAs/3mmIKK/6EKS1RAX7Bf
9BVN43GEJ+TXl/Q8WmMS8OgrNnirbPtEMYjjjanzz4XKMGsFfK51Sh6QBlm7lhxT+4LCXR1oKQIs
V6YBs4JnORW9uf1v6R6yLQGtvnclLuM7zGu/mOur/YFkr4yMP0MDyPxk+s93D3WdV0fK5W17YWOe
Tf5HWDSlpabgxrVZEcCgtva7bRzKM3iKzBUMd3sQXdzzCQP/vVg8WXx/dqpCBz3w75pvlnrA0ZBI
u+5abwpUVTVf9wN91FJFyG3AJdzvu2iqqAQ4UDuDF2EwXQ/1M0u9q3RHQOxJ4igu6O0YdBtWhIcv
BHIFT04YBtVpdRcaeWm2oirgrfAbbkNQKvBoUCg2WNwiV5DZxtaqwww/Hdj374vlOpZbwdh5dXWn
UCkMHQkNNyXIJwET/JoMhUtnaLkxKjY+djjIyAFSyHD7Sadm3nB2c8ELfUP7PA+LxagmtYWCyj3m
LyIuJ16rhaWTvEMNNie0peFh1Fu+SERBGv42AJ8g2Uo8kn++WeKyVe+JCAO4LXjF2gRAqJLFpz2J
nnSZn7azolmrsKREZttSg0Xy1WIeC/FZS1GnbG1Ki4lFD0+plW57yBsLuNHbFHoRdUePe+rODsAo
+cUhs8EDTeW4DQH183wAPBCGcWdLjvtLUwEMRLkPyGSo16fWDZKDTXFTWsj0/KBzn/0+Py/CX0JX
Ansq6aSQ9TDBTxK7u8CC/IZy2zAEYxc/Ow8MXU7oOaW2XOUTdBCoj3+8/kZVCq+ADllBHEHljKgg
RnTW+VtXphRfbBE3yPNL+qn2c5q+jl7xUUFwupRXLBVOZ1zFqyb0MeSekyjnalf/BpzkR6WsdpCH
JzgXRgyhiU3EWRqP8N7h/XvQtBZAbXC/nzoqcwzV1e07uzTTxdSvTAZTVlo7U6W384um7paMokYI
nzA2S7VYT2tmw0vJtuYjNker5zJA7nuOFHZZGdd14oYEdmhRw3BqNQ1Q8iPHK2RP8Iwg8skKcujh
FuAJR+xfsRJDwIKobDJXZg4RpBg6jRNQenaLJ4Z0qwpPbz6zdamcq20LbDYkvDPFp5Gwo+hd4539
9QdbzppVD9CVj6CzeMY9yREWyzycwKqOY7hFbJPCeht4TAbOly0tgUZCT2muxcMy0vb9OUjMJQZ5
XQM07PWgPCu6zTeFSthDh3Tnl6/P4fcZmdipDqRgp+n8mZj9Ug0s0XRU5fMrxLBqPNz7UHlMVdmA
aXcgusq+4p8Q9Iy+qxkT2bjUoxD6WhZbm/wwsUYhzzBcfSUwtmsmhyO7RJj5ByzNDl8SS0zl8baN
IhaAfLUuj+9Jd7NRCIhRqqINOZ9jzPkpP7Tl7fysCFn2XeYGDDL8GyfDeNjs6pRtfCcVhZjXW9WT
n1VXVWRFL6OB3ftMnOil95jmoUe33lZvQSNfWgEjrbyYJCNhx8IcKFxmO700YAtzHNIe07GLu9ap
UzExB4UgPeTbVgTLgT5LqNfQ5jN10HGgcnD1rlC771SJsCcCyJkHmdn0eGxZmCujRNH/7o7xadZ7
/1Lin+WaGPHUxcbWBAjAZwqua+YH9fteWlC7jRWKde4Kuh/MYSnD1lWlZTri/1GMiYpDm4O4FX7A
3fFH2HOGC8SyKk1AauBpw5OpZ9CUwfKBBVE8qU68r5iLE2F2RD9Bq+Y0LS1DKR4aasuStnQojRkR
DqmROSzbg69TDZReZc2WZCuCcy/COHtLssAQwKyMdIBkZolbvtLLQuO6/8TD7aYJP83xf92aQQLy
DLDKskKpsjdf9tjveo7tN9Cspg6qr6ElOgy4psvWzLcSQoZGTyUyU0btOmS9zJxj65HG8+ma4v7y
akFd8kDvA0BLDgDkNnSZgvfSR/GnjE273taEVrzk7SKNUoFUeADrJDCOFJDSL4vfLWlQMrAT8PkX
xUHc6zr6y10bcESaris83xkTtwfHR2Ash2C/PZAQuGW/L7jXs+gS7OGN6U4rrhoO4ckNH3p3vK3W
y2LENlgvxtz7pl6OkXrHHQw+zv1RjOgVKqXRoOosfAZtXbQbk7HYV9vcJIAeY2Od3nJVCp9IG4Yl
tal6fEnK+kdmwNiiRz9cfECYZCDZxk4VsnH0Hitks7qGZvHLzJvja3LM6aZF72JY+XcTLSwLd/pe
jpPtS9iq2drR3S6fi4fhZR9dYaIfbAJIrZfxad0jOE+3qu7xl7RpQ791UhfFQzDgCA7mKC7xh9wM
LukK9FqMrxaC6yo91+xmJ5aBCeH1zz1EakJXj/7Dx4QxDiRB3FXy85k1+bL2w95W6vZZoUihnCNF
q1t5+LVH3rMo4nF9al/JU06xP6g0kks1iYIWRqiLJ4dLG3FUKlbE+wx8NvOy+Ize6/dongxxLJFx
57xpcz95WSB3MDjjLOigdmGOW7bvDRcGJ6PQ0LKfH7wLgjHmJ8vqA/3RiYLCE396lqmin3v/nLE+
oDxU3ziK3hOxRl1CSBa4XKZ6k1GsdKbRX0DzJjJcEa9VMELp56yRVQaQwF3J1w/TqenkJsWSgxG6
hYpk5avykNJcc2fkvIXrFATrG4oY3syPt6qC8znq1eem1DOK7E5CKu8arq0fWV3AaPMAj8nd2avx
/750Qtosuts57epesatoG0PGvfTGysc1oVGsLoRAxst8Dz5TRuRVunaG5jPBz6Ru/SciXUvodRnc
3B+pYCkHP29pXsp7wKG+m/h17qAzCSXNhdNmUzgl538+CrPejGhftWaWktrh/BSxYCTvpUXa/BYa
HegeaRP157IRtQ9AX6LNq2BH0Wz8YU0AdZnNJ/LKRPCueEk+g3wdG4XD0RBp3JIOC59PcRUQ3hMQ
d/kpA3Kg8smvSI3pt5C569/sv65H75x6I3PhK+c760kj3rQHGtM3RSuKo1uQ72eYa+yxr7LyGpam
8w5DzXEGYhY/Aktn+QQTaGqeyRCRBBlmd9Xe/kbL0uQyL+cCp/2k438P7GZ3EwYYMcJCpudsfaOJ
9m49y0o7G0p4B9qNJc9QeC2fd7YEJ1Exz4TeBuEhjHJgV7C3JmQ8Czsd4oMj3zqbIzvwRU/wDLaK
4bSSCDrtLYOuNW4y0BDfraOYmu2QasiXSIBAs1EYmcPNIahAhoJI8C23yGYb3ey67KWM5AF5+xvf
nodzlWbHES1Cp6Zo7hFvcFHFwi9/5uYMTLZszc3Mmy6Ki41OVFLu3z96ISvQb5JrnYhNszObthE1
QB9epsLq/rziDdsil27+cc/upRIh3SWVfSat+Vjw+TKGPUh+H3sVfqYwEOSa29vFAY3osqh2TIf0
BY9F6b+mQFt2B0rG51+Vs552I3phEfV1JWjLgFdO6FqPUrxffLEkUg3N/Nq4JKhL6gY5bUoLgvJ+
plW92C8c+7DUxPamROqBiiJ6NQcrYH9ZLiVH2xUmqPXqh8ws3dT+XhsDS9ZYPBaQfGEKWxnkCvaG
zVoi6BxqzQl4zA4sdY4OmqUt5X6NPK2/RwgpTzNLOTcoutJUXpizVhTx/WKoW2N7kgENs1knksk3
BB5rwgDWmJOPJImjZSHfZkz/OtZhm64Pk+EcF3gCKs0nP07uXSqsQ5rK3n4zqObpl4mQMioVcPLC
A1RZXDnZgtGs7e9ZeO3tgkg8antDlsZE4asgYsMx6VjIkROn0bYFGvSRk9HB6L6LydZy1rGx4zeb
vMvWWNdLvMn/r2HOTn9RMRnrV7U9scXAazc0/wkRB+jCNvGhbgjdSX1jOSyH3ORr+MMcmYcgIISL
W1CU+EO/MYJeV6rpdDvzC/D2MqN4vK7BHNDOrkhv2MiuDcdvA0fYfdk+2NuQlAvWb51da+nbkgu3
hZr6d6TsHmLnPfH52DvaZqdoeqjg8jN0SY0H05+AyfouZObCIhovPjyVUkId4itca88MytJG0byG
d9EDN9CKb7RzICJZOACB+QgkoGA8XmgLCydeGkGo6eSxbkg5/epfsA38lChtiZaJveStWI4zEP8P
TYfbc2OtQk4clMZda2hUbFBRjAzIZhUW/G0x9oEG5NJ0ZgFFLk0L8LoLliS8Xr84idVllzFryKZU
qX7zB4M4CUGW7+HqivD3IoJOJgQ7OgOEiOE6rMteXGjZXBJ0G7ao+h2rQhHz++ntjC0oJeRx9Fj4
8wdpJcW/0u0yBZAyhjkusdeEFKbE3s4bG6Rdw8xw4xSmf3Jr++wAwd+t/NLqSC5ZGIAsT3v0SYji
3iy/eWVy0hA8Gph+ZCKAhW3fQ1hfDuKgLy6UzbaXOw7f4y5a2UQR3YfP8uodTqlUBHOtEjCTYGwJ
zFQtFZFtfSzoHACyWzpMKIu3/yd2UUGJi2/fXF9LnaglyIi6bhflo20KTj2SUF/udrFFb5ow0qlS
pS/eKth83vGLGQ2iboTKauQbjErK7Uk3hOyfSSp0SHJKexWzxejkgmYjPTWXyzT3dn/IPFvVr/mi
AnU67cz+V65f1iyb1mpd4yUowHTs/Ag3tXWtV3f7O2i+KWAzbyuOAcKYL0XY1azpgXgxcNBK02a1
C9sIa6OPEKfLOo8p3Mq76nrZxw3FsBMOdMzksNVL8RGZFTOaJTtDQ/k+W4yfyeOoyIwUBo03/uhA
OmP4sMOAvNEiG0yQsAQTx0p2WI5a3ZEmMRBnjQlOsyi4ca6SXxSndOtcmDgvD4rmP8bvaQfu05+/
FdCDpWYC60k/+7WTEOG7cW7IWYkVcR81wAJClhHMKYvXf3p84R9VPpnmAqrm7oXYMH3AN6oOGAae
Z3XlalOmEB5vnlbQaOslDI2ds13IRXqfWPVDQGFfB0i1/XMPkpXog29f4/dcS9x9kOz0oihEXrOX
8YtymjMKTZnpIRbE//Xm3XoiOMDjAkf9Ysj1DkC1OHDuD95Cd8U/Yog2ei0tauu3lkpM0uRL+78o
FNu+m/gVPuKNpNGsDysAUXPVulrMrhUMpvhZLohAX5dPpE2NaX8/hMwx8tDBEImW+327TzuskKzr
W9MW/kdBM0jX+SK5mXd5w2k7cWuEBo+5FNiO9odsi43S0VgtgzrHPNF6Ia3Btdq/BXrTDb7Oo8sX
sZb5BhmYuIYUkzk08hpsQ/bVrTWyYLrZ6+b96IsbKc9FW5oxze//cuRvW/t77+5d+aHG2EJYaMum
X5hMAalo6yjSfXI3NScUWf1cWKfFmyBCyJ/cEDASdW/Rx+BiLrxiDMmUnT3ZJesacyx8syzC3l58
RKkhF45sY99jVycXmeguvYEJqFbQG9hO8SeRE4wYve48XcN6glDewfB/JXVIQlGhtLWTApQuWfy4
cs3Eh48nal7vSNNHnCS6UUrGzluLbuQvlwFS5CyG1m6wvYqXhsyjyZpNwWU5dzpqUnBdKOKj/FKg
sZ/LUfLbZsLSo3h2vjxKLKYZ7PFUwsXDYn12gKkB90KdO+46BOzaPxaP5sjX84dGNOF6C+NAs2O9
fxRsTBLkYufjyfXMOH/RzyEfl+5Af3X+Ozeo4GITk4szWdufbZDJ9sI0rOpYsf7XLTT1X2mEUNDv
Pcwnf2DNhI2GlPjTczXDwxMjX7fp1aTQyoI4jrT/JOtPOIWhMwG4xOht5Sq87Kzrf1iYpli17njq
FZBPqErQvpAHmnWFjlepdt6kRW3bWtrStX1xS8yxHMtopr37IpCChKnpb3LzgOeH8pUrtWTrV4LC
TDuZqwHT2jmL51WNcgyb46bM6sf4irC2NWLHZbW705AT5nASVR5WLyLKfSMgC1b63bTlbeyIMlmA
NYRxarZ6hPKRPoOx+JFuHvzIoBxFcjSfV9IrP378kPkCTKtisaX8+JUd1/Juu3nuLryyNHX8iEQg
nODwq2WWWj6TxYRB/i4cILxBn/ITFu2FQt74QQWdQJp+1+xOHWb9ugIMLrlHt3m4f8Ox9AYn/RN7
v39EImndXqLmylhzsTvXQyfZIKLpJ95NUNT1mPUC1r3eglN78A5D8poW0XqNMp+hjOvw2gny5ZHf
b/8F6t4smZrrZRSqccNvmdWQvqueu0SVI5FJn4gSwh9Tejg19y/uVzMrA+3da6DwwV7qX4PV+BCL
J8XpN6rL7qAnRwDWsnGMsqHMNc7paNAcfJmBSdJrr/9CKLbM8o4NTx9/GVMnbhzyDiPZcS2TVxb4
ufJ9Xi8paQp2mbqXWMh2mJu00CSOG7OUH0ODweyzQnZ92JEK68kzXOrLJaTiqtrSNmdygMud7I/G
S4IyAChXYMBH35DFJyDMppBZMbDiB/+3FE1e+JEx11KznaOsQ3cAqFGHDXNeUp3R+WFI3ieNOmM5
3ZeDUWHPjzfW9iK+gMSMM+2JIHx+8GgHJtHSf8bgL4GwMMmNNAQINllV4XEknIyzSOlZMytGN40D
d+COGuNYwfev/1EQ6jvPyWi44x1bBxKQWXhnYIWWdGbmFX9Rla0DVG+MZRbznqgM1fu55Ite/Pqm
QG9naqxy+7ZiQ16gXLc0HYcvB++K+YWc3FwvMJ8ZomGvv4KmuQMsmfow56U44WMWV80URb2/8lh0
fJtG8PA5gDaT6+/EH7MI0oG536bdBH3yU53hC36Lh9tddFEe3fCubS8z+FmtA9Wkmlxg9BKwOPeG
FVGA4h5Ro34Jzutfq/fn60KhMOsiDO3irw4GHG2u+CG4947ewwqqWk37DCPHjmXIdto5tc5To/5c
HMed5gd+hG1Cg8GlnUP0qTCXbNkq/zeMU/BQO3OFX9fQggNK5K9omdm081RqEFFsD+hHXJIgvRyy
zK4idOnIf5m3peZT2j8bSjEYV5f7xEQu9tmF2A/kKpXkySmMXgTeF2Ge5jX2JOc6HOiTOe4qmNLZ
BehITL45WTkpQst7kvu8vsNzX8CFxkvSZEdK1dlGMkR+GthK1fIIF1Qimr1vI17Fs/fTeLNSAU92
/D8+829Qc8xOJXIjZbpqRFIYNu/FK8Byk/+giEk5pMiSuxxJcts90ert43bGJsP9Ohs23Ayoq54R
5X22MkW51zAiJxCIBAFuXzeweF2irrNF5MgsebnXvSF4egSLKz0wV9IGM7LJH/XH2gN1XIcx0ofy
w3OBH5D8vvTKqVheSZFh6A0QgIC5Pp6IkprnlV+9OIKwBiXx4jte3nDlYCXsA9OJSBn7WpA3wfbR
LHlQ3TWzeOpfF49eRNBGs+wJ7wjmNiWNE+/Kh1814GoJY2Hg8WefzIFxuAml07HuXanST66jkURC
rSXtEcBvV9lj44M1lxxZUWbTgbLEsXNoSlXPuNwtfo4MbMDbdDFXJbhFhoM22rysDJaHy27Onv/9
mTqIlgrJmeqC5qkdJh5fjv7vY+DZZp9wzHw9VvDGTi6mW3BPDitKo0xPYt3Fymfr63oWhF5NKkjd
Id3DDPE86UdlgsooSbceoAhTkfVHPDErjSIw777d9etu73zm5uNXNnz6j6ZUUPjxtJZOLiQzPM9O
nuuzKbMXZKYNg0vbcRdaV0PC2ch7Raon4EqJWxfMGAS4QWgObmibT4cv+S5d/alwgHd0VYnKUqnY
YHGKRNC7IMfIlMfbip+GKEPGu+ssQj++gRHi9Gd1x2lbT/RL/mOLCMw/qGKhujZH7LFI/2kz8Rtj
Mr90MEOgqAqyp/xnaFOn3JdcCxunRTFjAqPRcsbFBFnqEui8OLFPuFl9UcLWjFqvN6YyLFuPe7so
ygiRYjQU+M3mGERfVjcgp9W3Gmne1z3n/3M7hOQi3fzdARs9ELcU4mZiuyyhDAJyI0y1uPsXnWgW
Db2t4wkvwcXa0VtwNMyrn+uIDWejcZoFmp/WRoW0oz+vcWc2VstT7lnALRmtuhpnLyQEvUT7/iBO
esvFvVrIrpOP7pEtQdwEGEkMp13fXQ+6RXwSHTAg1rmNIVixF4Jzuez0tQEMkkPFKtfY+Oy+FQZe
/urb5wser9c2ZP2WszDbgdTl9jHKv5enB9heVIERQTOIhdLtOw1VYE2YzM5mf+yy+rKt93Mes+RW
MLzKavD5zP315GU3CAqmz9BtyVVMw0H/mpbA1SPzKTK/iBK/71BAQ3HCdmCMg+f5dCS6Wl4OwbVd
Y+gbI7zb64INNk3QqL98Y14qW/vKNxJwX71fOiI9Hds3gAhSycrhrtzlfptXjwl61AiQrT6UAB8k
8m0Qo+mP89NUUfkw4k/ln+IoVFGlGzZ61IUK3NOVxL3d/dojODaMFqX6DKN8+hTuRAS/gFF9iym1
9ms6lW9BumlSzcAGToxtrwVvU7YWS9LuOjepNlTPgZlucjw8GhfTf/EJZt04w7vigO6yOVkySj25
3vLZQt0su+5pEAVKdVN+lLnL/4Fx74kC5VwwkPLTtVnmmo2ngwo0yhRuUK41Y3xBOC3yIg5SqBXQ
PA7UVvYsxt1etvLM4ZBY9tjLkFbs8KYeIJFKqj3XjG3SWL28zp1TA6Nps+mYbTbL4tQ3x/aLfgU3
oFrwhJDKZkAuEJII5ecyU0QIXJot+gt4jmgz95V+3O+4gpyWPMut12jlH8dt8Zbh1fqqyDUsTUvQ
0IERvb8TWIaaEG1vEwxJiD64rrpSGN15M+VVvA7rAu1ijPAe8FNO9zGxWdEfdIGamd0lsdDdjP4n
3JY3r/SWiefyW8gkliqvVNfXYa2VsgyP6I/nNQJREavKhq6eWIj5rDR+hRDhN9Yqv7bHzlp0fYoK
FD5LVE/BXCaje1JW/XgMHLZWQcbnPDkRQFrP7egMOF1rfXwc78xr1590PpaF21Iq/l/bJsPKsVWN
hPued5K8wbST8OiJhWNbA98S+mR8n0Hqv8BHpjXI1aoX4jTrNpOeNKLWbu7pvIuYc0+YeeJduR79
YmVPwOjHmGF96OBuOJ4FnDNL+hdomJLLZJqqnwn2JIqa7qVDdJwM/1LQ72dGB+n8/aucM1Ct4U8h
gA5MBht6cHIc1VDQ3W24/cJ7Pb17Qju0kAs/LiaaqAxJnwpOMthAe819Jv7mu6L6FYhbaNY+FMWo
sQzcvw303a68IGP6FC+19lXRvAKy3VGpyTRqMRjnxi9dmJiSFL5WshS56jvDIJPfzkDUnr5BG+iV
4nFezRSWkxYgPcFtZjoWtviGDHOWxSsZ4s6gNmmA+Q+q/zfezqhbFyolu1ehV3AwIVCb6RUNaA9t
N9CRh3OY7jXLZ2vfKJdxMQ1my1D37CWGIPfQ11R54Ddh5ifpN0u0EfTC3wvJkna/nKUyH7/5EqwL
tJSoaEu+Wr0nCV0OqWhn/7ohBqPlPyNvb7lzNwLoSgnZiOg6rE8OYbfhgbxFvDyZF68CaVvzgQpc
UXEBpHCzEaEcWeP0J2RGjVDA4/AcIWdyBvrQ7qb0V3wcq3yzv/+moshmQx2lwf0YEDvYJqNWnIuX
eQgOgNqhQ7mzQufWsLPGg2G8WogMj783Buokr3v9eKzN0z4Vrh4bHnrNJHbmFuGT+kfqawKZF7hr
h+XMgcovg7LhjWY9NHvVFqKjjws+10AuacEQhEIV4x2SqK7fK+dVilht7nfipzIJXuKkRCgoa3rr
TF6xNuDsr5iIj3q/cx0aDbsO/lgE1Nz95kIZhzUKcDDbjuzzyTtB9AjPdkQlTzBKnNJlzJ+S/5TP
WPhXFDi0xwcQ9mbnrzTYxoR/T2QAxZQDwrL0yw82Eo4cQS55XIiTQ1r8Z9soN8SWr/TPVWmysaq9
4jpLt4IhXWdxR07XH65XzfGh+93r79e6PXDEB7dMHU3XC8t6xhJLsH6TaVyqRjGbz/QdmVd5EpuL
Jp1uV29Hw9i11BvvTFTVXdrQW+XCL+lDVsJMtMFgSxzmb/1FAXHVRYJahg2WTFFi/gN6oUXxdQUr
wNxLB6kKKW052+DLoTO0OEWfbQIiJ/y83rMLvsGy1YvGR+8OfRFuTW0jqDfFjGMk/z+xjw8yWJI8
pQkvx5mcZRzcEu4BSIM3KG4NzSSNiXT4qx1GwNlMlI4Jq/hODaRrJnkVzqZ/E9eJ0PhQ0K8xvAZk
l9PgwZpwRmlsKqcYAdehndhMqSk1dCr3U6LdGw8wvydjc9WGjg6M02pcxMahlWUiH6O2K79wXUE3
dOfZlUQgbD5UJgFZVcxH60e8jUFq5CXI3xOGIWct6vkE5kGZwfw56uFoMrubTWW6lEV8aKXPvBhi
FW+IOgodwEvz8yishRomdurb4ma4+nGzBv5Rd+5W3WYBjgsx9jXVs5Xg5RDbfaY/XaEM8OUZtzW9
FifG2IHEsqHo0GaQ05/yukuoxdQVnMpIW0imPMfvaxb2v0BHCiGb9rq7jpMSo/gNmxtCk7eDN5Ot
9X6ArBml7Rykdf2mE44WvwtPUZstBG9ic6rk3pD0CW3vwYynBKZkpdoiHTSVEbBvA5ulwrXh/ZQz
UyItb9TzjTdfqcjICR0MZgd55vTSkiPR52rLCDGxR3K2JLLvOM+JrhzfAYkIpJleeT2KArzejfBE
KNTWcVN8oS9dZ/SXL6xdXG00JrvhOYL71mIt8JnxtgnXYYZbvNEDOpDTjZXNqP8uT1VUrdK9H+oo
ftHmIr+KnyimL5CbA0oyudPMQq+U7q2EbofB3/9iPpvVla+QHsXXj6zvr9d9BAWZ534LjytnQhoe
X4MJ6faQH5KePqW2a081ylMHU8ZOiRrQNc8HlJ2qcbzHc8yaad+c60d/bq7L5s/kzIxa2dyADaU+
kmHqXM9t9Wpa0GWPqiRpt0Azt75hQbVcmcubWYbPOYrOAwaB5TUudYGLoXYr/eeGUhXDtLfUh8g5
L5Yo14EP32sM5PUwnczSnILTo23Rl3cbZbVlZhF5i0/7b1p3AtQRP0/cXIWWGPtJ7sAc3oHJWnYo
NxqPA861ZbbgEvsmxvcX1TTtZQghGvIRCDeY4oeXwTU9GHKBFM8iWNRsC0JD+eX9PXFkqthRhU4h
BMIKA5YtSnwkur3ZQpqjQeimKsvXvwYYBDct4ovXo0+f3jJ74Nj/Z7dOB+OJg315lwbu+RUrzHCy
myUSK8SkFPERWNh4b3nKsb3his7jV60vl3zVFWRDB6LS8P59ugFHBldJWdxeAjHYVR4+LajiUAHM
XIZnshMxDxWQ8MXZjlId8x8eA8E1+uR6jkjQJWrWZBGRrD0fkk2dT4imFE7bEyJZkIVRcuwW5Lmj
WuzixSjRhcX2zgZesdSsY0Ekp/aLsKq7xglUo2bbrc9Sk6BuX+PWmW8pK7mQm/Jusq+iF1JbVHEb
WvYKYrgwWLVu8A5+1eEFRsUJz4KOjPBJPzqwK2uw2cG2DzZbvKPUvobQBAKvc8+i5Oef5dTMxqJz
NpzSDH5M+j/clxZW2iMVnibDBfySj+SHjrdMTOy972SgAsYuuh/IDPZ7Pb0Vf1icEPe3fut7Rfq7
3NjXJhENM8tDKFJu/+7J8cWcg4+fTTno2ThAY7FdolNcP14fNRYNpE/YrHRXbkX/3jx8bHPknIOh
xhRoGHIxitRyvSn2fh8w+4qjdsZP5eUh41jtg8zpXqvmZGAE6oItXTBCJnab7In9Df9TJoqDpBpv
mJLiztSD320i4Vgfzv+l8zQGPMDTIOA1D9OvxMT5kmF5vbP3ZxMZa7Y4onLlpvAVLj6k1Ygy1ERl
Stgd0HCrkP5QEl9649RvdnIi3jQkhN8jxicOHmLwiQtgDSJ5f/Df05K0SHg9cnQzFuj7CXLAOFw+
4rmoMAoY62g6o5ld79EOwkvYtxBItCoWKBBoI0R3HlP9sMwVVHkrA556dmLVaLPd1yCeC7VzhUZH
HTmqHCsjs1HjxSgw9ciWQNq+whsje02sgxr8A4vM7AeKgc65/K+QbcDBbaxQpUEChl1bYGQ5q6VJ
ktTKlzLwu6roRFPodE1jF/TRrmsQ4/ygRkETgqcgWEBiGBalHCy0iES276kbvTPSmBmPB5wdxqrC
yZRy0fb7CZBAQshW0xFBw9OlEkirCyUey0z6F8czQ8OTxprKlGglaCvz0cJvNbwNL7mmogvxu0hJ
HaWRq5OQqJiLqR66rJ22xGf+f6Rg9kaH75UxEFiUjM/zkauM2SGj7IO+y81sWk8cAF9NbJ5bEr64
hyGSPSeWjz9Xtfkr6EJuyxIFCHnA5Jei/IjgZDTiXqnhKrd+MlADhaJHybbyis6t6GxIfGTzftid
Fv/u2m5bO1qQT1ycc7+3R1wBOEVoKqGFu9j9EReGRR6SEWuXbdDLB/ScV/NmG26EdStSPiV0ArAc
Zbk10s+W+5onpn392PWovsvBT/J6MRxJtuq9HW9h4eD14eV7dzX3Jr0PFmOJX4QGLrXKACqxX+ye
iw0sL3fY3/wFBSFvksO5eKq7fa8GTkNiH/SinwkY7cPbZZ9e1Ap80UFzfOD5wBD/QQTg7gJ/FQMr
kxW61lUT5vy8fMxlSx4TjKJSpbd6Cg79rc2Ubs8uqFwUfdUm7UfJNeUU7z9L8b5y8QphcVcVzwTd
bgcexTACTFokibCK8UTXHrri5OjAQwO2R0+T3qNkq9ZZ1Mn7vwJKF1wEsLRbMm1LMoOAI6lHRBcT
ybz9QRFVCICb0VgPZ5vd5DFof49tf3xAUkVX5WfDuHxMPExDerWaHWA4mIHbU5PnyOWLR+piTzZV
OMzjmzIsay70mqo+QOtoj8tEzvvwyTy7m+jj8yZ2vj+XB8xpNfRXCrGQMpeEG+ANn2iPmiQDMe+P
B6yix9oIX/ERgHqrd4/6fDZ272dK/VHQ9nBeW0pUtcDTsucLyWBZr4gbIsEjSSfTjkflUhlf8v5+
pPNknJzRTHNjRJhHRypVw8cInkxuaG7AdDBrTkFprn/Nf1MrRKFXfXgk436i+MkxoalAdxMUgam3
4jat29TH93yEQFMg2BEs1bMbNxEKlHM/nrOOyal1scqOnhM6N+mnYORaYyzUX5r7hrPgrW1/7nwv
Kg78eCQkjgkL/NpLqaCBWO3fuWQi0huj+3ljVcRk9KiFA98oi8TgqP2OJfmAUfVGHS/bCVaKRReL
76AGtCoKo93dHzepBMnAfJgwAQMiZbQaNOgP6rP6MdK1InenAnA6I70gvhunPHhT3/CsmNQZgkHF
O/t21wbyNe43VDpfKKgoaVUmfzRKgmQVuhynfzs8TDEK7aq0eZSSZn5oALxCzX1IoQ6j3sVvtrz+
GkALZSu6cW7XN05YboXGMk3iEX348SEjMu6krFjQEwvdbCvFKDUu6vnZSAKIKrOjK56EqC1fX7bH
lw0P4utnmWJBuaoZ3mSRhVKkhmbzQZlmDVDmGXkbdvOw4IBD94ALLT/gHo+5MYnwnZzArxaGGssm
nJqisHaxhP4eFYOarQv1aMcieUN1vCxwk0o1PoPxR3mSO2XJy0KnJtSSR1uJJLW352cuFg8d6WHp
eQnBSy55P/5Y+c1XS9jUaQRu9B3+Cilwb7+RaAF4N60l/6uYwt72609De8/uCIYuvvSnNFvTS2So
n+5wcv7iL37mQSmlufvSUZBoGDWRYci40KH9WYqPmybQ7EdYpmBfgPkDkffS5GjWkuTX9rVdjXBt
hFMsHNxqSr22pvplqJXWoOZsO51XytqvhEjPnACVj3B0VbA8s6BnRDhti68bChYl57OBuOlgdIHL
/ptbK7zZjwdLCTB6gVZJEgoBSmFy82IM8RV/KDf3dMnEBzz9F27uA+F5N8rFQGYS/aAZtuvzit+S
WkvvXB1EMCPpwCr9z4WzniqlX9v0Ew4Bo/p8+wWay18QEjfpa7qXMS8TCkt69UUI6q+ReLUpTWoT
rRzRyOQPUt/KjOdcqIMtN+MQXlXU15AvvlozMufOC1daXFrz3G1FlOVQrIM9eXFZRacpoKiHpCNh
ElJ0+pQcBIz7rC0HqEdyczNUjjvdgqrLZN7I+DpMYbrHLizwlwe6XbPSI/Jk7ZLBGWRnAivIyakc
/rx2nODd2IzIJed/hDbgE0qCizgopsryChq/SzZah8ZukDmEYCzUFUc+g+FiaOW+CE8pxQFDUI9L
IZLP69AnQK6xnZ02ICjTfrnHK3R8i78zaqojvYwNwfiSI7S+CKXvYkMbNtXRYnff9th11fUFkY3A
aB8FypjiqmcSDfk5h006zaLCn1afOV+v6kPfjLrIbPBPENTNZPlqwSlDng6VdPeOe7lGk1+iK6mS
zIaHWRe52A0rRtxR2FHWbSIyyQDK/EGZCT9KelnM4hi57fUDgW7e0Gptj/Nvv8IYSIpj0Isx1zBd
bm28dpBq3tsm0/9vM7/mYOM233SuvmGA+OUGcWZ2FGaDhm+cr2lifgs2YTzDeIH/Oqn8+xUBJHty
z81kfTHvAQvSolV5+h5kwx29qM5hs1WRoSY4hqFteFX5Kiadqzm7N0rN2XcKv9ElYxPC5PoPXZLQ
XfgvqqtnvQ/rUye4AnSYyWOR6+wjVLqulYB80bHG/yfp40Njtdwd3yvbLrDkWWdHI5f4XGBHW4zL
56g1/uZaNPvRtkQjjH3+gqJbnHAxQNuZXuhWYyKrlcekpSGP/9GhmI/IS0eAh859876DDPXnCTey
Ga7qg8LsF0x/AFD93UAgIm9+ySvZR99/SQz+PX87M7QtlNR5oqa5hQ8Pizuh5c6+reeIs7hh6ul3
k6rRKi0NPhWiES+cH8WQFJ4qTMV3McuIxT2z0tSIX9zfa2z3C1Kgo/6dMviyKvnhh7wW5IdahD+h
pvNWdss1I1mK0Qqs+ywEE/jlAo6YcUHryM7ewJH+j5voe+WsExdh0Z34vvjX8+orkqbIESiQux5w
6tBdh3ZmZDiYuMsHj0Iyix+y0Qs54c6s4E03N+SggzqVZHRrrIqitqV8kXse+VcR9n+wVI7kx86X
6qrQcnB1RPHuUYnyRo0J+D7imh7XBdXvdrWY0ZbBi7+bWWs+NJ7orYnxFjLVaq4vJKWNfiRbNCCV
lk4jyQAEMrPqoT5YezDxlcbebmJefQjq0M4hIx2zEHo9QnyfdDgvJnFQd1HChAzBtGaXRCK9JRM9
MveYoDIhZiPHeRo+w+Kv8ReycN02ipl7R6A6ki+z2VazLZ0+GmSxMRuDuYvazdRpLj4FBjEJxstr
PItjWR5W3pFvOuONzv9r4nOeHHur8V/Dz4oRS/CS+M1dzFrtZwoOoF+qIWCi+0TwFpHnMo7QU3Va
xQrAPaPjPyoF9AjqH3ERZXFdt1pXAb7KEDdtRYEE74JZ3kFHRUHXuUm4XwlRNHrndW8ptKUOfcWq
ofyi1iPvbN8CogAlq/flaWV0/sARB/6l7ZA4CdctqHbxEDjkYWvDlq8V/vV+AcB1LBXYiocqtoSi
CABkqL4RaSsDTFssXxTUN095CrA1mAxtHai2dfAJhyyjNmciyjc97CgRsebFD+laNzzxK/J5FMxF
9Yp4mJKxJtNu/1neZT8aUocDg22ejThwM60WaINySbt9JtdSBryYcXVUvc2NySPrbHfudfw4vB5o
kpHaIxtjqA3LCXcf714tpeURaPZ/RPwgLj2iIS0JIEPbrgTWIy1eDFiVpKICVTOzIMsDP8NhVWUe
lKNgw59Pfs26rbXNpnnG9AVTgMsr4RJWL9vijsCRJ/mAzIBLRqn7FPEuQde/9D+t0h6chKGcEz+X
dR5TfIcOGlmdrx1ICIH7kowVJorJtVhYEx2eUbX3c205EwdXP7+7mCu9ghnTHFbX+O4xZoJQw3ig
rcONC91XS8AU+ddB7ImutkbjOl11MmrHreSSBrS3HrIJP0Nl9NGSf2tpfdEFAEhbwQKlgHRR/d6p
X1vG6EK6pAayg9kweDqu+798MpTIE4kEtTD4BrxIKlup0afecCCUnLikOlcjfG9c1XPgNi29Bdjr
2txFVbnVpXO8PbBTIiCVNOPPlX3PzQRmI5uyn1CVscEngMCiakLrYbcUqvxgoYmfyRwL8N1T+Lm+
YFuNmpJ1D3ywG6CCwaWGJUJbZYBkl+fRligpG4dxtrO2zxWsvdQzeUAOqsbwTVT5l1OjCfDpfo9x
GGga7BwUK+hO6K9qPtkk79jrAI89dN+6m00hO4kABDRvX98c+wP0uybOua+yJvfSgDvbki7s7lRr
7A87W8Ob82f+WHLJERG9QXwf7EZd7PrrQODMzH8Xeigwi3pmwhu39HnIaidNYDOV2Sm0gEV3kP9/
DVFwmnk2WsB9qdWaETfuvMaXpMvTljuOIc1nLpks9MV5heWJQNvi8Z80gRTOtANdMbwLhllR1o+C
0/FtlyDi5NjNyvuUT01eICN080/1LelTdjKbvZX7uaF3pOYq2eM+tb6a+cnU0SBS5sImbkrAyV1K
4LO3auk7toxySWrezKK88wpj4qx6XzxngIrWOOaKvKiEpcc/VhK11M+kVRdsBc73uFk49AxhzNWx
OVltcl+HbBWWShU43v5sA3IdM/9l5nKh/mFfPeGNbRPWg/Bj5raPxAov2WxDAK0Z7XDPxVT8cPPs
rpufxk/QROs+fEk4Zjfbirab34sA4H8BqoyYIpbMDPVw3Rp33H7I+QzlDkfgbQzr0SOtnoUFH/Tp
+ZHx2DZPzCZrUorG0L4A6ZbUFhoXQmpBGaV3+LO9OnJQeHrXKsE5WYIqheuOcLO/nLTLNetwckPy
D1ZYSMp3TLBq1ER6JX5xU4Z94IVHSq/Tbf3Cv1UAEKjK37ayP07NGYMGwuGNwImPs25OpR9UqqIz
e5OyQPHQ3WNFIx1yKqdN52gkQg/ZGtAxGKvXoyiED8AmYhM1t9vNlLTylzolpaXKek4xfclCnTZl
LIoDRZuTWImlsF/fw5lbJDYMuPNMjwj+HYMNC5wYvwrmy47TNAFerR6jP6cWbMgqoH2RBpVmVQMq
X0s9qDL9PHAV0I+/viQAd3dSpc4JIgILLCqM7a9X+xUxMZd7nK2S1vYnCKp6qo9R5ZBUCQiqnG0w
AR5ztTeiGLNhLDHQ/EIQbt3Za89DwYpcIFza3ZwjxQfgQgTQTkBPX8O8pELbk1vlfrISG9YGQ5IE
Izc/6HSMmOALdecHylYkiouEPIowPak1akc8gC9jR+3FLwRtjn/jJ8Jo1sLuPyne006d0wpbEWhN
usrbwC++a4FsHlr+ao3OjcWHj0qsbSZOmRtzIfOdj43vbNnFyVfiJFAOn5bWF65G9U9VKD0xjFt6
OSTtZ+KKF8nBMF1KkJWI7OH2XqRKhumf6MLMQI9WNJCEjY5X+Exn4AYvlbOGHGzla54aJVPsaQ//
2rs0YjSaRE/TWLtfuqs0C3p11RM6eaNfUhfOBKSz8jgjhBKlRtAT6c4/wokgLeLUoeexkHRqAZld
PwAW/3W92FlaSEFW/Uw6+WTgNJA3GO+bNX2KJ/ahDilaeoSFyT+fkRLdNGXh8Cv0SGhnp41WjA53
V7fgAm4MTHtkChPSeN7E9pYgvakBTxsbH318BHdS6eF61MaCGD2vNWy873wf7TpQcVy/4MHJQAMB
/HUVXdRP1ulrE1OsQEEa7ZFAI7nQryav9pUJcPdR7iAWvouftXs22OKGz8e3kML7hX6kSqpoF1rK
SKARtH93qIBRsyYFjxR8PPGHSwLv7TCVuUadAdGohyXPXO+MA6bGBhSlq2GFh2N5g+J0sbWEcPXp
vaPXDX607wSRlTNf5QImemtG9OxagmFajh6+5OZBFljPBqlaoPU95o2PVicqGIKXm9QmzZmJhNTS
6lqTumOONkeO70SWK5tmTVLNTQazjXusV/yHSiLrz1pDA3RWcT2gRYGI1YtJsHXdDtvByxBONXXM
S8rGTFic6rTCceD226JGLLLR3YTrY7mREDMEFfE3YSA1626JsutXbpv7IDjfzEKCQ6J6fY4AwgpR
OoDgX1KCTyKUm1769edaquHK12ZJ5osQxQcXIBnoGw82Q8RoKcDoxyQ+6lyjVAfpinJ6f/6KWw3b
BVz4Pfk6jFVjJIetHdZwN53GHCGPepc5ScP6TFqRH7cIv1GUxaEWcQqrRMJTl04WywIcb/j4DVOZ
0vhMMwZ1O7ZUxvOKCP9z43kSCGOTds4AXVhU6sZXfkVhS6uiUIl7RN6AshKpA+FRVCAH9n1RfZEE
lN9lUrYsIeKJH0m2HenaSadZTJCH5nLgekUrN01eM71XwXq1CzqBk3W19fuWKefCiv9G1HPBjcDS
E4wwMwEyAlMnuHIEZyGm0kLux6/AB9/TfjKb6Jai78plfILZQeiKHPY97Y1j4bybFF/DBGiFgPQH
kTpkJJ/urqPRfFUaQ97MAVLjOvRHahzZOJtnDFtBM78iA/0KJ31KnoPEe2ihOGROv3ivo26S6tFW
R+H1nL1hqk3bEoV6mp3I6g4k0CM0Imak1EnpwNwXi7r1nBagk1MfnYEEdCVarB8oNfF8Y50q10io
vMevbs0cYKgiOQ+KMUBXeA984znRnvJUzcGTTVu77QNXAOHzRr21sAh3VteFuU3a5oVKqK5ZNQwS
Cwe9osBDE9310eTttSaqfufOxxv6UKY7yel2TP+tEi6XLhfDnNw4qjQkCD6g+UnPSorGTZ488cFA
Io72Q2OkD4gP0rTecWJKOGvjgMq8TWS+4Ibvq2GlgjdU4UXIOrDID3YEn8CZEMqxmW0W6bQkrOCp
zxAXPvbb1KzxZqgapNn34y1g7/xxfV1Clj5nbTOQq4Z1l9aJ3yR+Klo+/DFkT03DTub7aU9MpKpc
6TH+rePKvCpQ1GlITsERNonuaLrjX6fHIB+ZeYfSwG2ge3Xr+CUmiwWz5m+0dZhDtIwfAcn/XuRM
BUiU2G2kL/sl8TGICIj4DFs9sZ8aJPKknmYx/7YSlo2s31bLJ1s52WjhR/WWcp7Z1sY89LRV0Tpz
Bc7FiMrLsLf9dgjRUUT/1fIKF4hqGTg1XFtkyc/qOasFbeRq940g6Q0YCncihs+j6ocetgZRPQdC
m4TEyS1vGvHktgIT/qF9+l4Yd2OqPJG8KoI/GdmiH3X0c8O6Tc1dtP+oSaxhZC1Es9Teb/YUAoj9
947T0WXSaqExbrwJfI29SF2VQIpuSOjD8Vm2Xx+re/CAmQmKt85M9eniOP6DElrhltjIKFl5H2Ee
9X5OuhBL8biK/Pv1AtaASPxDL8Lol+ajUHIP35YQ4G8Df0XqR50SVLjdrtQ23NjgqeYfI51ePmZY
wTHn5urh5PDmAc6NDvViAap4CL/oGJoprlqwr8kfloc8rDGxS9IccztyStQhqmh3JhZ80ZB9u/rM
OO0JUgG7GQ5mRXTVRuepW4KyJxdtXCFwPpAUCrst2Xr90yNwautrp/xTgHYRvNxnPMvi/t4bZ1ts
dIbdu/lBus8QCR9Yvqqa9ozrxGtPmlFlgBV2IO9ApGV1WxYh0+iMUl66Sjn+6Yl5khfsfpHhiWd2
didEO6j5FWskL6hTNsvBZv5JG+4uYdvMzHkEpks17aKONqtGdh58ECWnkbyVLcxZdaNJMUoRRCQB
2uwuCX9CfLEziCZYZ3tnQs35UZYqcHA7Z5nkwKMDhpL9oC31tCDpCDOi0a3NQPhzPWa7IhmTUYox
cDviRGbS66PenIw1EyJPukDfsd1dujgqVKWtNSu3/Ex3nOYxQHtp7bd4bkDatNajutQAiGxqbYLq
AuaJ3EfXTiUWPsOPyzij0h2lmpjntgE7Bv47AqeV+bOjafmQIdzAil7tOXTViY8lDdHnFCr4YUL/
HG4wU7C4KjPKjmFHP6x88qKAC/nUVNrpdV1zxb3DHhzkWT9pLCDMOzD89kzeJ7MFfnkijxmqdxoq
MoiroAijw7TPmZW+/16KUSSuJsfR/3GJLIvFjccMtnNOwYhXWP4vM3fsuMZNjdtwQLNQ9aWYM3H+
g0GIvCKuRg0xKKOB4FvquvOWb1C5Q0HMmuL+Cux6iD6I6SXx0jQvSzq/+Rcez2lW45ry7HdrVUwk
LwoSsy2/LNg5DlikZonAtIOEZvO44zNJnpdWdO7fBej4IOXZAExmxhRRoPa+GaEwoRL5U4m+ZX3Q
bsQ23CZrJZZRHrIugj7+0W0W+DvapCY1HA5T/srMrPZcZkHhhzfm463+54m9gSr/hR7PjRMKXKwe
3tl7RRD+R5TJQY0F6EdLm1lK9dSj9f5XuqprQ+UpDVgp1kp7JxjxID7XPmJwEVuww7C68WG0vHLY
DWwJOXgovzTRT9PfNWGP+uSNT5KPubDOP7lKpb7wSdWPNV5lJU8OAx6KN9/P0m2MbvTUeCdjitRg
fE/nv8FfWe0rw/AvoeNPKGUP0C6wvk4R6lnv4z0IPsZCeauu2wVuZa+/TsfsiBjzZbnol7GoE2hR
qAG04evldqBn1zMI9Qe0jyWXEctIk8lzifexCwB94726/W228t83M8SHioejf8vjEIPuP7lZ3j7s
ii62otEzOnVDTvmiG0PbOuyit7T673uKIIAozxZ0QGEBBrGH8hVwr+oLNmJV9N6AKFibynrmTiic
4jJT2Bxt4U40CLevvtaLD0wgqWUdKE/FPiH+g+bqZp95pe+FdEn0jRSwCrsnTxEimQmCTd9ACdMX
hfPXVUqRQSWnbcZEKFUVMuXuukv7gBhqb74tBg+tFs8RhittYhRXNdedfdaExIkjq9CTGgy+YU8z
TTRCfFgAsXsGD5XDfAsViaUvEHvj+NfATJT725XpoRnNJLtv+itr95/G3RJ457qmCCFfAVk6ewJm
sS7sAGw61Qfw2uZObtJQ2GcGaZDcprmcLqYeAQajGr4Bnn60/Qaz1iDYrey02o4wsUdvqKv2xKPB
wDXUoft/UHCq1RNfXIIbcAHtdSJBfxQwtrYKlJHZzuoI49EKtHXDSwLgrUSDXrQLq5vKSFvglVCN
aKOoB1QjHJn+WR6CLo3MTN6dHlHkVSkz0lEvhymQft1mgYOp04ztckr0phUWpVUeFnykVA7xXfGj
vIquCDXjgGB070/9yjcHGqmF6gr5vxKwr+WGBSsjw1fy4BfenCSHLG740J3jZthJ5k8SwdqdIJb8
/GFpOL6LJbBhhlkK1jGVWPFwM2naEk/YN3o56jZq6TbkM93SJsf+p+4D/Npt8gGOhFVnsCMsUxom
jJkPVAdUBKqTmOn8s15NVs/VJVVNayCCou8VzQ8YXz4jFiXi4Qy3HOCwhOm0GKTWNWVtfdM6Ntba
nPa1OnV+kPKVlYTouH01FLSEk6/OJ+XE/oNMWzMjXMYhKH2Xj/MLrsCAx3RiAM0MEC8we5IOHZCg
2oARJlAu/t5GdSSJsaZhgiYwjqI5dzGD8hksaYzG4u0R2WwA0x63JzkggKqYzwmfWtiV3chYtrHn
GRFoXFFZhQHRrhGuo4Y+tnjQutYDur9aGXEhuiqVZS0jR4MSwJfpPiGXqrkUoFstHRufZkDwIS1B
d4JFbqhs+QmmtoJieJG1KjWM6EdK03UjDHn/orpBbLKLRIg9+YQ6A2wjdgm3p4PVMvCJyCDm0OMl
w7rfggyuYca67/4WMER8n6K7D6avahtPWjFZQ8hmrJoUN9QG8R4LB1PQKhHyMuhgtN8QFLjsBPM7
z7VCHjAV3sPJzM00hCjwZeWzkBDUtOuZ6PhJXj+1VEdeoHSnoVNmx7dnSWxdb/EbeC8sbZQsnDeK
KzuD96jNdYqkQOmz/oRSTP6BhnDXi1YoFqH/JYGye7yIKBBStSQmWLHf5GpBcgWMi/WzvKwv1GV3
cCoGcwd3Vsx0EfNQIQHnMej48ZcFl0/LaKn6zPwtBc7p5XIDf/DlQXFFoSa0DZCtiBuptVs5igXV
/O/G6+1UHnR0ZIRF+77hvXRvBlJQ5SAP66AmOwCML0kthR2uYkJJE7i2sbxPohk7FjUq3vRMzl+z
RjVQmiO3b/RLhsYVjQel9sMmKF4qFMX3UDTXy+RxfsdkEs0VpvRY62fJ1wFAC6EZNtC8RBh+6D5G
6eLtcfVjpaIyPMjfY3LvsVBch44kfmrHHo6yjQMF2YIri0PrAQlrOst61REKBSFkGN3ZiaMKRdfz
7hWysE9+/AQNLE6DEPZTEAVMc2sHh59reslUJdp7Y+lIh0L+nDQn0Hxc2OXnKFn60xWnV75pnGv2
GrTlakFiRxnxZevOpXRfteo0+JGVAutiOEkW32iql/Z+OGdXNItwolMJmYJ+GvyiqoA/pLsPlEPn
UXGXzspiqY5Yl0rq5G2ZcN3pkYtzzFWCwipz1WhMXlxQUkVbovWTOWptF6Xj+38JLmzHJo6OXk8J
eS9niM7jofga8kWU5f5bduJy/2ItFPX8oGUqZ71unlBN4dXtEdrkiunEB8saeZ/sXNri7Hie2NY4
h5pdSlf1Pm5So8XecASBgX6ht2/Mh9T4EHI59zd3NHqmQUXqjefVqr3fkzuEtIbla7XL/Nl+svDa
5xHZcPLurvV4wajIObcVrzEK2L16coMNVX/JWADbYk7CMsiP+rpM33EyIdj089jmlLodrmhCHLQp
Id+7wlVYJC0RQ/evGFccl6RhegBuoOD8Y/eZg0U5tKRRnV+a5CNotoTRRR/kPf/7klDeQThzz5ET
0PjcXGIWa07Com4m+XdfiTyUTGZpKw1NW0EIVm/eLrAfadd27fuAkxKAS8Ry9EO2k6eD5QzTrkcp
NO69IEIC5jZME44N2fk/yMY/DAcOtaITP+ZxKQrZVjbphxr7BnUe+vzaabXdubJVgePL/DRRkCW4
FT5aKHLzOg05chpCEqqVZDFTVNpgOxswUgeuLBphoHNyFFLBygKWaBsZ+QwTAovrsPYYNN7d38B7
fqYdLhO57h589Q5YMQ4p39Yu/tM3gaJAS9v3fpq1sk7sgpFbWXDpGB/znsk648owYHAddY+G3Oe+
gBxwlMqllgtO2R9+5APJ0M05GJ25MBONNbO/pjP0cOrnkMdHivAbwlDnpPUD80g7+WEFOfsomitB
8ySVpHuDsP5c8PBgJPtZ/sJ/rG6sUMHvsy9Jt7tDJ1iakl3m1rfeOfX7SlBk70T8fkjhS7OPnlEh
SH1J5YPaZzOaySwsOsykEJSZO6T0uo0aSw2Y3XOqWppHaFqXS9l3SecQihBQCZ9A33P/vsJTX+cu
IpxxF5HpurmNnIuGc/wLjuV2NI0Im4CZn1PeTXSK61/CRmhKgXjm1wgp26fm1ixxPEX7B6swEmmX
OvhmzjTBQlqcifFXClNow0It6px29P8LOAFuKUVAvQoreUpt+SLau2LvDpKc8p8iohtmUpBkQzOq
iddBrrlgNm1xp703mEQIWQo+zQk2lnrQ0dVmumVsaGk59CsjjZfix3u9kSLevDL6ZHAkuiVR76/H
fj+UECJNyptD8x2AU8iK2bgPWyU+Y4PAnVK9EZKM9kNixB6JbOedyAEHHsfsZIJz5G14jgzNotGA
2LpPp90YVoJnRc/TjTUcnzpIHUPqTA/wKefkOKZcochoww1+cB9qtfTbD4oj5H9uOhUEpKjnOqGI
lulnMWJ2HNg5dXtP4JPhTaawE3NoqpKEwr+Zd9RWiQ7IjhsNLBLXk/AdBA2AV06aSLA71f4K2/vd
PLvh8uMaEy5nktr9dN447A7bdtAcWZMReYEK73X/BxnNhqz42hsLVBWQgWaTqSfrv6hH1ZmVIOsz
CNIsLQeTMWWAhraIHeXsfImYzAEohZvRxVgAce/LuAkibaG2WZeIGrReCorQHWmhlUcGv6lgsk7j
kSLM+hF8zQRiy/c7ZRyE3Ku2Xb2wDTqlBVPnfpPDIR3swDEqntJUgLP3yTCY+3JggA5WqjDxIlL5
MJ4Xfy8JCZ8+XqLQi3PER3t/ZtGZgB66luSBo45Dn8mFN0cu/4QVCkoRpbTk9Dy9SSK6M4LBokUH
usq4+RMPxdpgejPSmd8Hvoq3M/GG1h5TPfNJBduoB2YaTT8VL0Z8FEheFqw7einBWKgRwSTjUjr6
ENKc10bdUsyHvCuCR734DOa6x1SZd17hIlg5OYkuICkCZatIv8AZGpBHb3y+Yg1nUt7PhVcsDyog
va88fdIBrBrOLCaDISN01Tztm1dRj8wfPfZmQi7jIOQS0E5ukK2EPS2w1Tb1Y4C/wTYBnca1Ziyl
u8lddMrjlcm8GlgGRzEEVq3MSPHVeC9yyzIVsVGgk+y6Ej9eKUFObyDYQYPE6w2t8yPiNFexgv1t
ywnzF1sDkmZWRbK0wqk4sn1Yhd3E+EK/D5OUu6jfnJJEyGKKhLDlAdEEUmbyS5MZrZgEOw0vSxNU
bV7Onoklo0G10xI5+7GSZcd58HDyPQHPLHfdrY6TdIHxeBcrttJ+OlWUg3y/T3KRJ17P0x3GX1PR
NnjoDoUu2fT8r42nr6/9ZYIl/h1SWTZERwiCOIWAS7pebIFpsMQ/oMxzzR/mnTGBNNkA7K86Jpk8
zyhqPJGlSBcfuxMdMpZc4LIx3tQvPgesif25NOQLXfD0hUu/7S/GYX4axETviGlgRTf7/oKCYXhH
EOvHbR82dDUX2kxOQibI+hFGr0dsTcuFuHHQx3i/LtBxWjQ14W6h8tdRrkHYnDd8KHHW7SWVBHza
vC+OzJeXe1+HUunjT9ov4Wfu93wxVlv4eoEKnr9DcO8JZ5rQsB+qprGTf1nZE1ajXDR8q07Mw7fw
RpN4NENoycFzB7/0pvCRwyjQ/c1sDgtcbzztAbHphgSI2anwrWkd+lIO6Nlvn1dIYeAxfuc3WFll
WolgbaGUzcIDTzoKYuZweYVVSuJukmYmm2xQbo4Sl4qOqCVCHmuxiiLmI9UO+MaA0ZP2t1cf18Ac
sgdOuPE0Mp+WNYx+IjWbTYzCb6MonWHj3pKb77SpeHJjUGLQ2jfgGUwPKrzIu6QZwFaxcqtepOHu
KIVPbj6lzbyCSVyOI/QzwguRPxAuusSi04XdzhQiWMtzNFe5CFYf+QnlGrodRR1bl86xBmbh68kO
zROvulmaHs9Z3PJNOPsLPJ4x8Zu9Dkp25mecqmE7iv6gpo3rbmebzBI+lJ9hENSG+Bev7uMkvBef
xqsBx6S/FuDsvjbsE/sb0MM8+J/6Ouoh9A3xgWaI9inEQGKL61D2vStxCfYH9jNdZNx1TGZVoOnu
LcNpBh1HxDn1So4vTG0dpW5iwcVyIRQ1w1EdW+QQU/uI65Kuo8nKp1Q38oQwb9es8RN2KLKRBLDz
YxzffcJEAOquzLh7s3XzjF6OGVnUgW4J9qilmSXgaNAzqeaI9SR7Lvgt3D2GetjKM7Eg6P70x5JI
hQ7mXMy4wAe/OXT10WPcMm07VaWP8Luqn0mymGaQk+mHIo14UTj3w5RD6JQ8yVZ5chMT7aQ6sTWt
oPCC8D18OjgLsY/s3rpPhiAkAyKkdwmpTNPS1WjvBYYdz4ZsaapaiznH+1HSKQHU6jkXdlCoIP0X
WANBysKbs9Qcw1Yhxq2OIPGCGHZlgAHLR3BF/P5OwYGxC++Gmp6+1PA4WGcMFJcXQ+/THCce38Ga
xOq9tymzIk3OKyaBDcW2/q8e3de9nykX9jekAEZObCT8NreFfYVyJgd7NiVNBN8Gy+ueUzO/lO/Q
+USxsS2QsGHBEwDGPXuyNyI6eOLIINavTQyYsL034n6Sgut4WIg4SHCNzjydumJboYAQEBTjU13I
G6GnPDhDEYNm7zqzH7e48sujhjoDDL8boCUXXBDhuhFlo9Qmw1qxJWIIoPhhl61mWJMx+yOoAWFW
dDU2kiAir3dQZLqsciu8uRlBJt97c3Kd/VqEATfemiUErquRbXFvh+SEHzogaXgIuXsVVMEipsfY
DLSpfFZPkqbglwc/0HRz8xuZyT4OZhHgMNd9hBbrF1FdkaqfMaYW+441EC2csnFcEaIrmhcsobjo
g6T1JCB6W0DdgJt4XMMFep5q/uVv+gNP6DbDMLu9+aXV2DN05fqkDKOQ4l8P0F3Lsg/ES/112vti
eda+Kdd4bFZ5X3BtLj3zn0K4YzCbOjhDnLbscHhzrMNxPHZ4bHePMMxZPDLbXsNQzyLQ+DoJKAD9
UqTUk/LdBL61iP2b5Nz/I8YQH7pCfi1l4NTwk+CC6NXaeBkN7voB7Wtd9lJqm8tPvgHDFMmiXe5s
JWq1CNabb6A28KnQVmGCGUjVZirxUGSGAPKJltrbH7Usup5NvXTMIa0QsBZCXL/1FWjkRui7wvIF
OzDVHv0kuYxLwBt307J0Lyb2AreYL4tKisvTA3A+WKl0n8dircwzs12LG706iZsw7FI/q4imvKYa
DxdKYJ++Jpk4gGFCOBLY45vmW5riDJ/NP/jj5gfUzlEHWOBphDOcVuBaGEPnDVPNmqiB5lh/IgVe
gpCWP/WW4aoUJQR9uPvBZ/pa0uWVapS3mKRjThOBQyP9+gnVLefKZmuSG+TdF8qmdPyohr2D39yF
zENgywkZ6pCyB19N6vwI6BoRIBLyhQdfunH8+vpuhA5gzkHZWCTmg+5YMAiW8yQsTbQ1x1FZRedr
ESgrKyBCP8kLUKtLKjlo9TOrsexu8dz9SFhtBAf8MsTsiSjikt1hZAmoIaIyRCLevSgOuviVHYGV
xbdDkvL/MbB7KiekejZqf/xwIMPVT0bfNlYxys+aGeJ3fQuPqeBh5xrjg6tSn0d1U/gJB043fJNw
wJX+lsuoyNQ/It2eRjue75KLbKhetVkKDZ2CSKSLnTIEIbPoBfeFaHLSGIzOS6g+zMg1Fspxm7zl
r9OT2PrK+fvHZF2tJYajkMeepV8Tkvs+W6SRlbnB0Joo7cN3hypYpxBogVJs8I1zrGYijMauhQvX
vS0bkLbjsY0XWG8EnbObKzN3xYJRBjaAyKottq/5c63hIDodBzdTKHnUw8JdfEJ3k02CVbRtP27G
yCIo+lqx+48UPyplJaJGQvR2QpS9tI3TyyYzRJ7C3V2Lnn2B/D5UDTGjTsM0eS2VGMBmlk8GAaup
DRR+LUd0dOZxvu8SM6fL4yjpl9Qh18/ZJLAF4PYopO2DD7wW7AzBX3cAmd5njFIe+egjXUjYZHIF
zvI3JECwiPS5azYePOt/Gh9Mqeq7iLnMazqdGPDyyitNspNm0p1iVn51cQh3xsk968qG67okMqgG
z8+LP6AlBp2L4gqA66RGOMQc0kumTHNuLjgYsUxuhr9STbkcoGlsGCcJXm7LSOlVO8wU4A6hlrSr
TnhhBEocEjGXCl7OIOSzNJWtLHHjUalBjX4H/9+YnunNYYk3IwTh2x7Ya3n4cYjeFtYp3LZDXvOl
46DhXEPv2cdSk4Zn2s3padq/Qt94ytTZk3cUCl9mdjbZNP/qkPPE/wXhlu1JAtMjbL7oxwNCi+Uh
iR47MRTyx5w/cWDfNSFoNB1sDSmeZ4CONNXXhJTFSnd1eEIalzh9YTQiNaigvPVr7Y6AAMfs40yw
dkua3l12vsladI+aXDttAwxxduGBhDkduV9Dgad6fQ9HCPk0yCQgsbu2QPmAwED/KClS9fCfoGac
Cd8cywTh66w1Ro1ndhxnd9d7bilk60e0VgcfLDu7f7fWR/3E+/QiObCaDa5ldkL8cqEQPv6a7HzM
RDVn7At0QLioRiwIImHyXfzL8/73xMu03rVnaQqFpzi8TuASPK3JIa6mv2N8/Jxp9merD8bsBEqs
oO6XuQGhFqcZYeiG9JcH+LWDl2kKR4QfcUXrRHzXbxJxUE9BBSyzxTZz/GqWSE2NnhV6b+qWWbqP
mQrQGu9EHkilfszLFTmkLuZqNjqmefD8jA5LuK3+FMVieYpeF2JfMCBW+RBa3dEk7h/uawLjgUF/
Npu1DYnr/onmN5VGTwLO7khS8kDXmKsdbfXgeegL07EeuIbuncUfhixQJxrJQhsp141VbSvxdUC1
m0KBHb9Hx2MghhpmLc8EO4eou2lIEO/qPa9CPc2123DxQVe06t7PLEhcahVJr32zOORvCJ1veSRc
dh5lh84SyMaF9c6QCJVEu0qAVrpwK++QjN2gryPx5mDrlmD5+p28ED3dy6TWco++ANFEbFka9Cal
LC5tbx9HsJRAGFR+6kGHbeXTWobI34V2zUD0mDodz6lTktnTMZCbj1ZkPiSE8la+AQ1IixBp8riB
Xx4LmO1BRhw5dCsxJjz88rGhghZBPyR3k3loLXf5DY0wsSOg9eqYOJKW3MvRdai0GxuNvpnVHAi+
7IGkGlaiookQNUnZ58R07WsKo/c0KvrkINRkGXKjAjVOh2oQZyhEz4spTB/odl0CaYZITR+81bJL
oal2DqU+AU9s2WMdgferk+8k1PsD67uccQrsAJN9CMT/N+YrfkQBBwm1yvI76SDjbhH+Wpcs1DBU
f/hHVjIPINMj2uY8P4qxIKRQA7vgJ+L/5m4brfq1YpF/oFPLNecg1/hH+JH18l1ikf6iTjKpP8MS
+N3/fnLfF1FVqTYs0QnPPfVkwaOmzI32gzScVFJ6W0A7UiwDyd7FESkGNcCQfTHXfcAiadp+2/G2
XNvEOJn/NNofrimupZ8nYT1aB+FxsmK3CeSSxSY1pnF3T5NNEGVbSmi8jTnXBxotDgI3jU3GXTAt
Xl5cGSvhjoQfvXlcEcCFwEg+gWpdGdNFGoNK/qaOxLO1d0mUFDKDm8Y43KzbthgK8+7kKQOZ5Psw
vNkUoLRxuNRtqIl5rAwCHiDH/P/UimUZ5a8/y47y0vTCWETFWq9qiyMT6QwVJ8CfoliEidgrSFvx
qO8ZD0I+q1lDDUbw5S5kRW7/AAINEb6KI6leG/BTd+QLjdhpfLLWB5h/DsgwMhflO/yF22CYiit4
8mIHM5WwJvyukkWroF3hSt3u7SYbKYUoxeIVcl+FTPshnDrFxcvLo1HR4k7nK6gWluXSpUge0dZ8
jJlMBmCYf0lcKx14HxuwooTuHiyyfQKZgxFNunzOQThN3mk1ZgeOzi1EWiKtlbCIV8YCDmlz7QmW
4off9giHgLDmui/P3eSvm2I7nKzikINdMBESYnnbZ/V71k/R6RVp9RzbpO4pb6k6od/RlJLzqxxo
Um4dAn/cpVfhqIl31xjgkjQM5v5CKMtH90MxpcH5VV8ksa+3Gf8OA+1u8qfxDEhPJ7EJAq5tLpQ/
SPayYk8g6TvbHiVUu1HDhPXh87kjyDHG2VKXPZYWkR8euN4Zq69UKlHZzUfMYBUJs91ngVSgTPCA
QediaAjGyK0mVHnLpxAIhKtNAf8U5JICoO+Mu5boCwjjVgflhgAPWzvOE5/AsG9ikHNN5Tc6Qb9w
52QAAoGFM1N9aCv1iXhjgGxd3oc+D4E2iYkcOQq6Lxhx+qL1+SiNRI9tDxefI6XZvq4AIVskeBxX
c/c3mjqyeL2GOydQubmu7dJHh6BopKk6aGJ1GzhvHrE9wFIyPNrd3DdP1RK/UAOhT1ynysLT2LYj
NybAZ7VdIzZtD0puiOKmAZTjJoICdbcdKtWMGnshg5ts3Bls8MsmSlebAXWiciWeY/j5TQcjKmH1
WWqGZXAOpT/ivOdb13nyKk94S2238xAV9BW8xlWVyH0qSxYy4TK/MbB14J1K+gssnEaAFvA4rZl9
4MQ23Yi5+rn8/SedJrQu09u6IYSk76y7ud5p9WudotSdFMUhs/SGeSVAxHlEimSVcstpLzsckG8V
LgA4KbqBeS1y7tOM++DY1ZAQdZLfSibA2xyZ00xvShfmEwYiS1oQHuCUdtUchDGOyBHOpPnuIBKq
gXM16+rqdJUsj40LlrE8mKJsV8JtE37i6ocDN1dQCZA46fRRjKHNdFYpoB6KhgAvSkdTJcgD++/J
f0nw8KgQul1z61UAyUWvGh2mSXJs38R488J5YgpszlOnn9aruGIGdFUGBEAQ44IX9TQYvEFxY/Li
W8wDfG6W+ZNFfx1SiaM67c4kmEaq71d6eBN2MfbLD1yNA9gGeaoct4zbBX8I1pTIvMMIM2BiyyS3
NhPjmIbziyZgPQwNSZndUGRUB9+VtOOAWpRPkQCm9ky+B5jDJj9qO1Qrq/e1WeG+BthsD66UOUX0
FPGG99dfF4SC9vGvBvOKFqR8aLZHvWMSOnV8o4FtNPEbUkBVzI+hklMVLNgaaNOsMvcGSY1WffR0
l4U9vhObu38oOyYzD5RNjdQMlQxN6LYA3VcDNASOvaM91YovHIoelWxPmDBA4OR0dVmWyRHaVegz
ISOG1B8FEQj17gYQyFN7DGg7QtJ4G/9FNXt6Q9+FV9N00I1i4WfD1HAK/miFb0YYWWofAKxQxClj
m/Zs2qGmXKw8MkuwrlASuJkfCTxWPVh0gJWDVeqwsF78eO92TF2kYzCYM4CQFyzAn0y5ctPOqOMF
ILZZ4qM+a7NKBMC37xW9K79KuQP7L3+j1FXp28r93J/JEz9y7UaN2AgDFZP/IYvnoPaeQlarUJ/a
rp4nEoVrib3VrxTrB/bq2xt671FoaffgNSsjOmpXPcvefRJOhQ5/qy7M0JBjCA6T07O6hd82cZOQ
I6SrIs5Uu2qMdL4QEgrNwul9FcTowMcCcKkDS2vy2ZgHz95N9zVnizxcgyru/KBcO0UFkaaWK13P
oe7/KdWKvO06PDFyhxp6qZ9DzKDVWoKBGBom1vZqYyVEWlkzN0orIeOO/PjXqNvo9wl7rR38zVaZ
2W/Zwm4RaYWl78n1NaJDTwiaUCImgxqxVYejvlIGNXFBksLjCkDDrLR/WNjj3RTo/ooG6v8AzbM0
l8TbCaR7QxFVH8RLOhiFpXLTxm4dU3okq8d1IBeogotDqYn3bk29fs4j1exUeHIBDgXpboOlHcWq
KlGpYnzBrvLPe6Mevc8gI9KvoDezM1znIUN4DPOEwvxUeLCT0nezi599Rc6KWNGDK5DGNtAuLHcT
az+qlkxxCkyJEcepKwPK/L66Q77FngW4cMxA7YaPFdKgmTXHUZadtAnYSifAjJRK0HQVyJPAHWuG
EDseZjFg3+8deGQKmqWrsQL2FBL27xHyDEkzcPj25pPuzlsTN6ulmHXvIX+O9zWL8f21gTRrrsc7
CGirCPf0ixeD0aqA6xcJ/i7cqouveDvOyDSSBFTOGNzjjlG2/AAisFCvp1f1g/i3KWIthVji55IP
Tov9AwrqtXTtMx40OrygiMUGDBYExaHHuotPiB9ysboPi6jGu3ACoTTrKIyWPbgTtomHln5lnT7Q
UA0tOcZyVZMMIKfjNSIS6qxn/bi4bLIzVzxTpid7cLisrZPoiL/eJX6917ZszlS/0wR4ljKvzZZc
yVPcrcci41BeMLUTjbVVboKnfT9s3fn4xFEvgCEmi3+JRNyuNqLZpmt4kTXFUkqS3oIjM2GQz1vi
c7BuZvfLzI52Yj/9tJ25PwYITA76tMmW2ItQJBkIu3IyYk5Z/gVgYGjPplurSZMoA0mi+Gkx4jce
jwAZOUHeyBTYsS3XbgOYQzEWEZzpFc4VKEgXTlZFMNdweXIWhCHoprDozqJNlXrYxh0qY1timZC3
6+vXF0zvK/YjviayLnk7SWcS841yf1X2Mu4dER7VUPrmkXN+L1cqZBZTmLb8NK6iWyDo5diCBDOc
+mZGaY0ra/pUiuITr7kRou9Hfz9rDrXvhX6XfxjRzfFXeU+TMqS4TFhVLn057+9g42iAUbG1twun
BUYKcmUJezsJI1FBPX3+6fetxpb2wU3BFy46zGM9ZiaXCyf7VZbnXpk4rwPE09EmmOiTt4cuN8N/
Oh59TBbWBR0+ew3fCQsm05EebyIXLCBTY0irs+ZxEDlXIypNy4W94vqSK4teDO8UanRP6N3mvIuJ
73zHf0b1RX1FS445hsMEP39tAa0jw8mPq0Gvkihdt3vGDI2oR+EO9c9+K6NVgdmzrkgsIXqwvZdu
VX2JBoOWfEQIX8g2tUITWP4CUJf8gbG1Qi/xsK4xY0AHel7MB94DfdpnHFh/5Teb45rSr5lRg8xZ
2VNRUmoLZS14jb+V5OWbkAlt36SGiBwBkEQdDvcR3bE/Rp6D87Mh3auXMJzDiOOWH7gZ1T0Ba4S2
/4r4Y/cVctKpj9uj6Pri3HNQYJszZ1fl8+5zBgY7GpF8G+pDoVq6gyF3fbTE3FkUAeqhdkPGfs5Q
/Svx8aHibadr95YdXfwIpNBQ00RQCS8gkj4jkEjEYNSNHCCg1jutQDLmhlnPhNLl8kPVTvEf4hi/
E00ALXQh5GN0rcAiwMwE7zMDy92hiLWVuNtLDOb+ktl85CJtWWbWaj82X4Sa+YDMuPTeA0/l9M1m
/kTqZ9Ny817Io2w69ZS5RkEQ4A0Xx9bzIhX+Nebg5G/7pE8dqygx3yh9Kii/9ORxUNZuOjWqYmnn
1rnJ87G6PCohotPMBULgRuZDRl7I9WMvS4xgrYeJYhkUgwpJ+w1T03VWbEooaFUPwkelM45QFzxB
gz6e34GG0+Y5gWSgUS8VcC02gUy0TOW5xN1J6EL0/LBppO1+xhve/jGzi59P3o0HnkLt/qXJazAf
wlM22abSnw/wp0Sf8TPRQbJkc/M1NGDbn+W7I9PjiK0br10Gf8oxKO/XYAo1UL9IHxz5cQu7ruop
6Jwlx/sDrnhVHooTZ1/yez0F5756Sj0HxL2X/G7OLOmvmPyWQzZewqGChimBqOG8zN/bC7Yq/h52
RK6+D/rmJS1jgBZPd2VoQKCn+5BLLhdvFZ7aaXJI1GA7tT0PqkWWuv8Oxen26/zxwGUYJdhmgDDK
RCkPj7WOghDZnG3yHMsuhJJxAqxjywdFvmnAWGMa4OCfWp4h0bsmEjk0GaZOsG+Omd5F/BN8DJk5
y63QKW0Dcqm4279athy+ECXK39cMZ8IkxbB8O7bmZktggqFNbaYxo1TsVOYu8ilBOCRAduIb1zBZ
ID0j2cD77jLCoO68YaVByXS3g2S7OWg/t4V+oujZJPPqoVqHU6JLBv9t/gzkccEXWeqSg1zP3PBV
JJk/XHDz6HRfDk/PRFzf0jUKKGO6KF4QvyRJc8e8QxEvZo6anTVdW38o62DQEk1JiLzOiEKwOxMd
T2vnwnKiAKeythJnnt0lkctPpB8lOmJaKhoXCzODzp6wT6jjt2SOxfpaykHMZquSrd6gJfm0zWSV
mV7jK2ZVfMKbk2CCzRgoy0yOZnDXQrEjDlu/rAKLyj3eja1R6w/zDgiMO+4RJDA35Ov8iDntcQy6
MXZEFC/YAfxythmnBLSCvjusmzUMr054Hvk46p9p1C7YONgjChAc9XRqI67x9HzfQFFlSpm65k5g
NFJ+yuwf5FNdEpQglvXHl126Wp3GCexkLggcXq7a7POxa6LFsl/dfEtNMdxw7vJjMAMOjmvWabOG
q8M1DJdMGVOebMir1iW96CHu39kZ9VJVyfOyqIAZ0yot4YFJIuPu7QUSuajhu/HnRy/xkouImXzF
CxkFb3TzNsysysDdat1S+BQc/AaeH9IthYkTGCmXLaFYGeqvg7fBGrfOiMIfaPjjTkh/9jHzLlJf
F//tHTFoP9IAMPn5U6xOqYQvJvCK3cEvnZDLQNzBz3eZc9u/jzS80+fkpCZK8jWCM8T60tck2vZD
RvJSCVBVxOnqX6YXGgWDnqh9nubFxr73XPvCr/qLpnTuXXPZ2b5SFr3UJUM4w+wylKiG1M9aaV4j
HWZZKN1yqHIh85tE/i64wjohE/tyYQPa6+z+X1s1mbnqEYJDdCotqoLXcB8xdmkY08XSxsxGQ5wH
Y6fHGhhIFe/km7fFtGymBJnbkL1Fb4zDUHaURg+Wa5URqGgVVCBWXit+jQMe8vqBkFCptdPAXJLN
i0nR6CwfAEpczybqKg48eb440FOAvxNcu4ONQNOUYBQ5Ecv9g98FDATrsiSUUg9qcBt4IxgQeeSD
H3Jv7PkwaJYGnNpFWw9qAkpat6ysNfJOXBtj0IOaLGCQLCR6CvoInHcZUvHFJo/VRXUoW0GjOHzL
HoSoxfE1vwG7I5u0DsmtbEgaqoUFZ+SGIcj6VQBCexun3qgDXVT5/N+3fE/f/C55hGgpkQXnOqpe
1N6nwUFXoMODA64K8oThBxEhMsgTgBjERvcQWh/qlbpUl3c/JoViVkl0hAvx+Pko/zj1LslAiBds
4LJiZwyNa9LXO5mhvAjJLiZOXdGENtCHrfL/+OczR4eMYYutOyI3TT1usAFOIuqBUQKZsPkaNuoQ
Uh3i5lc+OrjS7KGBgMAOOi1hW+HNRNB+eKBrCEbjnwG1z1wPTb7d6eEpIulXKo5I65NZOk7Ca3jq
3Qbo+2+Za9es50ZkFwgTXmGQg8RgHNPZsroKHnQ9ZWJkEk6EnJsinVz4nwFw8oB6dtOvIM+ye2xD
06/AEfKE2U1AzY+bvZATW1vBxPtB4uvUxvjVICrDWmBUeVy7x8VBL5OLPiYcuLiC2IFZa+pJU1HH
DA4Js23NQq3wFfHAos+hM3vuBwK657/zUYZLEab+ON8mf/D8vfXWX4b1DeLLSKt/u3lIyX+K9qRQ
HiMYbuOqsfELaNlhNDYZAZLB9+tGAT7ralNTf+Qq1Ss8il6Uk2+aSED+wZGr37S1xTTSbxMZgCgt
z17GPG8zMp2BTkcG2Qt3jm3T8egc9PSwV1HDOLotNgYojMM86dIdsOuHgRX056p4g61g/t+s5w94
vs4Wn9/YNIB775ui2iNfHb0ULnLAezG1HAx2ki+sz1xgnuGT2+hnnuFIApMUjBZmrPAsL8jXcqxe
VjfkfqfN4UD7yAd4Xl0IZvjuaWLcfENfjTt/vLTsFnRG/m2+gIMhFomV8oOgAG40FU9vstwReipi
llGCfbqB3oS1WRdG6LGQBF7GO4y6hyY3Zyg9iB93Ew6JLGRzjvEOAdU4lQ+T9VnAheEpNcOQetn6
KojO+HbOy14sTGjmomVTnUyylcGVdolj8RejIyQNOvQ3djBY/CscWsc6wPlfXWGe/ImSQ75SXQJw
mA+NktfdjIcmSuzOni0wRZG1HWcDPmC/VoYJCcwz4EsAxwW4lxYmWcn1F45o1PikHg+5pWSFDJMZ
etPFVNhJeEsbjfeIbnH1PUCz+XvrlMnmxogln+fMSsqwmN6FPrroHnhPGxbKDQVLpnw7Pp5loXy0
e9PqkV5MdUy9299DR1aLXqXkerS6itBKL0nz0I+yNDpQqP8fQrm9U3LTwfsOts9ZKgXLGys59+I+
O6wIrhiYFGfQis7Nd1LpZnJRA3+pG1StNTpTwau4aUhwLL4J/q6ABOnZdsH00xMeQ8P6XXZ+Mosa
XyZAbYdpnVyxGPEFe0ocKXFZhx/7pDMSgw1jxQniJMVCfrDd2YBuaYjZpV29GGPLTROu3c3/g4EZ
8o+sNQFyZ4pFr7wq6kUWetVzsBq2DrCrgHeePZw0821+4A8Y3Ho1QTWzAE1oVL57UNxbVovZoSPF
Xzg/wf0ztP1cm9QbipWJp6TiLrtLa9Yffw8h7tcI0FtMVH73hcJhEk9qYZIDdzC9Al7MDH7dyq2f
cFmDAsxDS9Xo4R+XbeMJ1yDbsFUzWBJ7HRcvgPvmpUZdNRQ87VnwEmdtxcHgELlkmXW10wHdf4LZ
IbvXX+NgLjWbVO9xuuHQE8O79eBvc/nU3YPqYu4WyZyhD8kw/0YetP3e4CAsQOU9VLMYx1vrTJMC
rWngaTqldYmaAWLzS/b2WGRQZIKQM0Bwl1YZsPaP8u2CyS4kfLUc4xhMEKGZe9vcHhYiBpQFv5cw
KgJMfsUGaFIBGmDESG4OYZ/C6NcU7y4+Dkr7TACXoYTCOd1tfMdow7si9HVcyY0yhJ1Pq2kKclDL
8dTX8Vi1TdvaTNwuu31bMCQ4yx+lVlVLJEx+AYWboGAg9QaGUwTlEPUUTWxofUT25c65sOjNQpue
sGO3BKUTcfzDiS7g2bcHaYpdnTWMUvtTbaQaeSRAQfc6U9td/EH0NQSmZBHJieFaZCX1B84fB9ME
qRyzU3Da5fAVr/oo1WKRgUvOheXYF6K2AbW2eK6xZkMtdXl/rHm2imbIix0B7ZeeOO/A8CKq6KhG
YoLKwgudT2Y2qfWZnGXOw8AbduJ0EDT0QuSpOlmGstZ0tgIIV68YSK07HLs2akhkPHG9Qk+dsVjc
lvnyB2t3vntuPulpIEP8Wwlr+MSS2g8pbyeBfxt6e5FUWaEHmIBeZGriJjvFYVZqAISXxlXtydBC
zGiZzAqEIGI9mMH9gi2Cqu+aFu4Y6NCws/b+wI7OTV2zV83i16rBwO3F8zjno/tXODnRNSNBch7p
0X1q5CFv+p0PO82L/xN05i4iFaMMmHshQIymU2Y+wIVPtQe2hWaaFAI0ykeVX3uuFGTNLJI5PRW0
uZLW2RTCI+jJTBko71uudLnr0NzH4YImFzR8XfJpsfBbd3wFnxBSjwpWILxcsGAsPb0258o4v6rO
1oN4t02XfkPmSxJTbt4e6gAXNzXMXfRKTxQkyJ8l5L6D7I4xNPjtQYnaCmYrMDcZ4ZKi8M4osTj3
YD5sSRaudPxr+V9AukS9uL8JQ0sOENmQ9xolj13WEyKt5Qx2FDUIcdGPDQ8536C2zjkVP1sc/G+V
xOwdFF0zxfDidiNRrdhJ11FheCoy++MxGr93+gPQ34YJg2JqIe2EUcfS2xiwk4P0ZOR/Hm4Gfpto
sB1jH3h9AQtdaU9qTN3xk2a8NRoY2lt7QfqqtnAsPwypNwOeFO7ZAfaMEsFBLAuHyHq3/2gizDbo
2zQE7PKEbs8sptIFnctQcWdPHJO/w2auS+5ZLoS9Ka7KTckLLXYupWiklhizY9SvXqO8OgrIQmmx
2YP1jNDO1NugaItBSxODBlLycSAn29ChrWiJBUz328TMuCMq/0MPgq59RjoHJfJ5BqeswXYnvzug
vUSGFjqpAQ8VmGxh5j4yaSTJu9GzZtPVIm9MTsr+KmI3Dkw3mmHV4Ui+O5Ro39VPNXEy+ZT2U8hk
HM+eCWGOi2bY1Mr0to7QGhmLghDhtAeu1rP0tH2wAHyIRg1A7Uc6H6RCB7ELk4XNo3xl6lPN+QfC
9yxOjivUJBIMmN3HBb+xgDPsi0xGva2F+WLag31YH10D6YsYCE7KGCtAiToTEpPVmcyez2raAwlx
rtz7Dvf8G1wWa/RCYSozX34++pW7+aa3m+6dfbJyWN8dwGJGWF6sKh1GwId6kXhyIJIDuoSzKne5
mz58uDKiyg9GIXi45dGXeFr88Sn0/Owvp6VT71+MTVCGi/Rv12hQoaqu060bLqnpf507TEw1jf5e
L0H0tLX+gwGottLtAOmeYgy/NL95zCK0QQdb5K+WF38nraBuFgemawFqeUv0ZOl1yuVwI3/7ofb4
BTcyrepzHr2/Uar8fOwV1e6RAM+FObSRzwjYEDLSu5IkvpRl8uavPWo6yyPQz8aViowDNoGbErDx
ldq/KUmPgrT7Tcn2ynwMFSAc4/BbQV7HTzTh9XN0otlN//HAR7feZaLmeF94r7YXoMLH5pfTfqeC
Gd6/D5i8+3/0glKkOZAYB0fk1IKzx8MR2bh8CMenyF3XRWLOdhju38UeaenDk79O99M1OCr0FFdL
mgY6cqnP4RfXO/PZPB5wPIdcz4myYhjWlHP/H9LoQWWgPiU0/q8UfBFoWdg63mZJQuMUQjv5mWrd
7NwZZTHvJwWr7wKyEVEleb8T31ZqTLL/I6AJF49t2UWsNuQL0AmpOeO5fQEyAVEyA4aXtThDx1yR
V5WooZL7XB7qeUbnnok/HKk2ZCcFM8gPEoPsoYZW7Lr2Xc7AIIY1WTpJiDe1+jXN4Q0Och3XQAEb
tYKevdTpPO0pSK05Cv19tcHgpVqIPBHa0kEJVc2tz76LUbTlLcxNGDK2QB7zUkTCBU1rFuauZAvA
Jv5saZYNqSosRhw+vye3m4FeoLtGOyAVcU9vXynvAXBaHFRcNLzEFdrSElD4FUD4jzNgFAQhyZCX
1VjqhJZEWqupnGeJgatIKEhYknJxQfh2Jpu89bK2ZiCxcOZ5XX6ES5z441i2dVouXyAhtQQ9khIH
NnScydRciGHwTuuNR79CVqFzGCc1muPsdz1qbEzikOAwQl3jvRc1XGa8NeHcUGgGeXJrMgNc8hWY
Wz1KGwPVNvfDg2sj3lELmcE2DapA3clKq/Ru9+JeU/S5QJyDQ4QYZcfkqovhEDJHiNyaXdAnDyPN
hEICr71vktOCKROlJzmimXJUFgCZENl72KKSFUjUIpJDYHUS+m1LZlGqZ45ukZ71xZsuYxHL71YA
//Bxl0pOy1c/PYmSCO8X1AtrJ8RErZ22DJKkbyuoglXcD1csIl20aSGPcNlZZQ3HPGe1/0AYA73f
3Owvl7idq3dXO8DyLhYCSjdoyCvqJaq34VtgMbLPoh+CW1eMeF0tUQTijX0bxmTb/1ISSqnZVADf
d1i9o8tBV5RZlp+GQP6eADaoKXaiDqMo3X9lCC1Fkcr0whzz0WStdyidFIvgPLHERd2ftlOqjz7G
zlJbB1rdj1HfbeKrf4hiJ1xh5Xr/lLSQJCxsfGs3SkGPFuQ/6N7B8dNFCeoHo/qGDX+yNUhouS4/
axQgTLFB4Ya43gXkQSwngqN4OkBxW6+662HQfuxSCjYy7hF/1s3jVGGbYW0hR3jNFc28nE4fbwCy
uxAQGCDAjxrdER/cnlAU2vWJuwwAR/ANZIJen8Ba7Adw9NnYx+FkNp/ZgNW0vfeaU+QQwkOLBwxR
o/pGnW2fjmMElxPF5Lp45faCs2HGOLN13wGvOhHBZA+GMyERfOEiGG+JztdVfx46DOZUVE44EVRL
QipxRP8+FWC1C6SqsLYKJX8bVnPIWMA9Gj5q5Gd7AgXpkD2SY5i41F12lTjK4TqKIAXfclt1Uz10
Gc5sfShg/S5LCNGRkBcDS90QEOcZqcZiMfNosQhHA7hUUU0mt/JA9l2VpQ6hkjFaIhSwtIs7ifv5
fDrqNpoWaeihvXUAk8MnowuBYDey3ne6VoteSx0Qt+EphKGnqsx2gEX0swjDrF/jPI7XeyxxrVBT
dTuqDS9M2r42ohHl0zPHo/rS724bIvA7hd3Wj7uO8QJ7ixvE7se7VyChZ/wyvQHALsKotG6uR6BI
1NjzrisprrMLW9in1IY5FEgDhPwgsl22GBgg8X0YVG06lUsCEaVyTnHN0oG5cHrw9xh9wd655Uhg
XVvMalgIWMdOm8Yfq9hnR0HjwNijJeQm+ihxYtrnVB3ITEGsmHFy4NHpRrmicf9h5NogjQqVClyg
6oBEj2vnecCnHJofNwO9Wakr1R98Kt21+eDLzus0rFPoqKRCU+r1MDrlGG2pku9rPue/LjEFpFDt
7dCsc2yEB7R9YAMNNmitJtjVg2Z5F9LR4iEMonH8LvrRmZeV7ZMjmRh5Pf0uQgTkzq2/8GxtXayn
ls9S/f/4TRjSLanNrDg4WUP8rPEE6U1GxgmHdiXyIVxQUDk/EBfa4xEYa3n8Y8cDEgMt9sa2c9Qj
FYuaGBvExVqU7u5DRg4qnx9viXwtZzf1HtByQIJj1BcAojaAwgvS4NoQJVWYrAMQd/ibjqDEgGpQ
qq/0bi9g7XQ9O6f1WNl2DTxFgZxO/FfPpxRu7uixou0jzwo1NDDmc9RRYBYCRexfPDwIj3ei9hWp
xKy9Z/JnXJJC6t5lZcz7P1UhKCVB/JVId+kcdqAN9CEyVIIzGZSv+CXDB5nKYFfFxH70d2GyoJSW
VNU/3IBJ09rmHcLuZkcPgNgo3+l9VJCTH1ZVnpg/YyBO6VhvcBvWXYpSFDkQFbsJrExkSdktc11R
em8OdbE6G9C4N8W8gkj/S0z23uQAnqKmQbZeqHBEPmqzCI09ot/48iWc/4bi4ywuCXguHG7Dz3Ac
worptSvnOc4RB0GpZBxupUbGBo0il5Qzb/hTEVZ9Vnw2aj3Dpzn+VFIJQsB/GXUIuQP971Tr7pPA
UjFeGCBQXVqwP1czSNJIgIiNSbf8O4Hww4ZK1hzI1hpMhU8AQUGU3xkj2t9LMMkz+473XM9Ik37T
Ovh3m8P4PJ+Dig69lz+QTNtowiOHmKc0x760KZpdLWQcMvwHEkglD47kwuBDFPzvXdj6Cd5hGIfl
E/BiKb+fXt7mz7DHGKRMJ8M7g7wa/rhbAyS79wviLDZCAk419GOULKTtv3HMkAsCKJZgl+MH86ys
FCnhvXVYGeS9vcZYQ0456GWYw0P8uaram5y39P89SBjCOuq+d/eSAlAeJzso/+PwEAa8hW+Ale69
bVRgIlNCCKJhsUd/xFuGy/XmkALWT4iR0AXstf0fDpOrBxzDc8W3EtuOaimA5w4RD+8j1ueGLHmx
/3Eg/cJEpCZPJwBi3sJ505CgmPxgQD6eCNeZoVLq9bKT501iykI00LQbw0wH3re7+3jEhulKVUcv
AazUB1QWuWfvNZQBgm4ul7Er1B7qQvPXATS7oHqARwXNxp7PWpUKoY55rT485uorVVTMuD+zH/ss
FttVkMIIlKVszjKA1MgUrMNISshzcQqtGUcniIj4CFHqLHidP1rhvkP3jn83CQNesRhywwhY652i
ouRQNit7DERTfhHB9uEAOG4b2PcwlNKexFCvflr0C67ZPqWJoLOOfc6XlkA+vPMwqzsdYBxnfiB0
K5OPzftItW9ubs0deSjfLSsSpi/VWyEJ5reedL4li+u384zBpYPouxT3P5WIJRBKANz/1N/tVdP3
mCqCarBak2IJIXh20/lb4NIkESdXcpQ8CcgMKwc8w2TUYeBOPR74Q78zPh/fA172NSkT1/6OIPBl
bGzeMUwRrnP+WGLs/K0xJF2zW+oWus6+7uJYtoWYD9v1COK12y++gACZtV6QsQscTUyTx3DKhiH6
h7ZMGqB2XQxaTK6ATDGMZ9fcTcjEkBJlEQzW4S5YEslfqFy3vGKyR6/zb7TnD3A4fHa3/U3Tx8dh
YqRJR+W5AUdX0C6gmBMYFyphGmHNOCZHRPwD0ea0Q2gRlqVEQ+KZA/edzHtJPpdEIjtWGiyBe+Af
VPDtw57rJ+rh0Gs+OJ9L4jCIoQdK1VgatMmU7jF6u6EnL4CyzhEVQA6ovuZaFXTEKdG9UpDLTWL8
q6nndP8cMg3c92perIJtnj9X89ddmvWZPPTBHcpSTRlCaEAz7HgcivFf6N3wixqkH9Ug1qeNS3lc
OjzF+euAmZnBJ5MYXZdYk55lYEzc/p+LjZgYKJPX4YXSY6GcRF5bUnSTv4O1h7Kyx10EnhkR27dH
cxE1kKOP9UXwLtX7gYvicbuyrVBOJOiCzZK3GCMG4ln63SwO6J9refBdzVxb24SuRXWfAXUjEKAd
Toew4FsVOsBNZQ/sKPdBR7psJ7GBFcROmV4NOXG+ljdlIAADKp/XkL4L/dBqKbU8du61iBZ8yzxy
GI5khDtYU6K/aITr644VlDJFtYrAFCSafK+KG8uaU25aJzPn+25RNCirRt/UqxQz5nBaNc8FO4LH
cEzvriF/y6Ahta3aD7FPgFXFdVVAtLgACgEjDznStG1LvfA+Wz4TsWa9X8jm8BFUkHoGogoodn/k
UClPXXGY9I2an+m9GCirWCnZET065kfg+3sSSCkMhbwcpkzAN3i+lkqefmdbpfu/UWltUmj0r15G
mLrMImB+jT3gjlvE09L4kD2j/v0c8G5Fsa99RKFsSPgXxcVO6pwrWgMXfh9aFTbw4BIBwzzjaDtJ
KQas1qRLkbZJToCGshulo0jduzc0hz9SVFRINdCEYHoBT2AxZYoliH25+PnUCk7VY6qPkNeyUeEx
5OBCekA3nqMC+uz0KRz79RsJQbC7gepl0d6Adm6hILdxB/9t0hZCldjEnLtmtIZlRrVbesF+8nzD
BMnaaCimkKxJYdxC3e5iJ3WHpoiVNPckupDlavl40pJFXJCBmOyG4uyQ7d39OzLt02MVWeA6DGBa
UfaWg0JxzbsBhJKmZNw2tjQP5DnGbeXfgQuLhcqKH3m/C7pUjMDpPR5o/WyuJ61rBvovZpincgxk
5vCElePlvsoxhGrMJW2c55ZqIp1Efpv2qa2yLS5KZlSpoc73HYf3Gl+5hvz8+Q0WOojyDucVkLdM
FzrjxRkPQ3O2oF8ZjCmZUX1oOn0Z10Gs8D360PEGap0tGNS8BEIS45JnfDJZ7KuzD9HbmfuI7TpH
r9+KkgXogeY2g0kjxNdxEwvQwIShyhEp3AeMk4vEZJLC1ytUIJHnZQmhSR46IdZz0LJZHTIHwPl/
Ndm+zRyPQvcgKCzYoeZXYysH0PY41hwJbff6atuRIWI/F3zO6+XnV5M3rGBGl3gAwizryuS8o3aH
qVUrBIPtSaHbwGgOjUn2rcZ8nrKkimCRdfduc/N1EEGcWKnVsP5k0p9rh0OEwJRXw0RcbGJpnSOs
FkQus1wyWpNGJTY4poaWMV+LgwF4053mgzzU0hzL9sY+wpdj8USK/fEv8wU2fdYpPEeodrc2WYJk
y9+adb7N13S7euchAdM3JFd28slqLP1MWNp49aJyvYZd/GJjLUqNxduoCIzBzY1zEy5PDXKGJjCV
thw23gtjaGz9I2ixwFI7WL2RUcW3MwmdoJ3YEKg1Ew+CnNzhGozGGTtABB8Mj0aGhdQXrCCwxlIb
Ae/sDuzkx3mfap+XZ/bt7c4NtjH8jAhFmKR/kM1e18Ud8LuJm7KpL8YqNaDMQiQ8NNlgdpsU9VCA
4DhegfBaXR8U8t3zO8TupCC1OUyO02cOxdJQ0z6LHANBhbH1+RSp96tumSjSYrrcY5wUxyRwGdts
kQoV4ia/CL/1oh9/MSxo8hU0o9SjWFVQ8vphctegUY38miVARp95x0UtOdL6oMvNCHQy7EZyNd2a
lVS1Dx7OmZ6rRkqHGdRU1+J5DRpeOKywnck5XJ4T7JluJFCKJLRyPxYA8eFcMqrklcZan3sJZ1EY
hV63OQ1yTHsArpH+MwDHhzOmXKYrY0BcUhXtlAc1N0cGPVt6DvuyhZJAuIkEGVaAc3rsFUa36nby
3/923q7sSsusi09+A9WWAVDL9EzTu/WIaeijwNLWCESbHlLkghf7+qWtfiIOKCIhWZGCcbUpiLXR
mXLJc89nLlQPwPc2EqWnUFsckRdhx3Fy4P4byvDlPFVgQ7vPVj2F8i5eRYNzeDy4URxzndCgZ6v7
ypfD8cBuTe1MhNmjrcJC7ldDdF5sSJXBB5kCJHyYy1+oiJVpK6dq4cqiBXAIsGpW+7lI7PjuVHMd
lKhr2mBU14BnlRou3j2PIJeMxcrCYmR6vInAlsSiwEt+etAToiG7j15evAhwyfDFo/T+irBrfwMB
W9vOVx7/kTi+iHy57M6uoOWuq/Z+olVuZKGv7IquKCIBg3mawXy3wnW6AmD3o/psfvW6oMHZLL+q
jyoIxcHVs+58c9tzgbEv7ywhEK0J1CRqoTzkxMB35N8ntFkTvN2qQWKu7Dpr7QVr3pKEHrm5VfP2
2Q8BCt6IaKk8oCXCj+lSaTDddxV5+Ui2pPI3tNaoSEfQQ0ysfXs1Yex6IYJG5BANPPKjZ3r9WiWL
lUiMIGt31d9upti6x+pdJ0e5QLN+pAcV+hCSZir1pnl/zpsiIE9/j3q6xfqoTqKvW7lefJ4Cao3v
qyODPrm08oqSjNc4rup5VvKJkPxHYq0B39DH3OIAqwsaKtK58EefhaL1FT0sbYsyOGXGnUAMESA0
YUq0nw4n5qP+hQ9ul8OROWI5MlXwnVWh8GoerU6fnhew+R8RIB/o3EdN/jLiecpSH61qZKTqGt1I
zVbluEIv5puinNxkD7PUdzXGbfsoxb9NgMf5wMfMn6oDnn4E1iqr/h/j+vBUzf8aAXQhB62b5SMw
R6sg3QnXro9LkqNtrYEyrV46mmdJY3Iiu4xlYitcUpU8aIMbNwkLll3A/Ntcg5aUYVBmCmPfQznN
opo5IqqK87uoJ1j8L1/Nv1swsr5jn30Tzphhn44QszRse5GXtdqYSZxIacAQzAvrKIF07frvy3lQ
dkeNGpJgNRKReuXu0rcN/jGe+/JTQ6LZL5HIegmZIiSNMF0lQ1rAKhQYQUzkQh3x06KQv4DfpFXX
rXwtSlmKZlMuCuKkzlJ0BGrA1/mmL42QQ/FHC+jgniNNA0HP0eptKJjvKwdMWSvYWuxGhQmYSkPb
9Q1RypHGUy05P9bmN1guJF9anxygznnv1afSYIzEjGao4Hcrl4EbvYzZ7TOksqpU8PHNojmI7JyG
mtE7uPzewl2xrJrSwBe4zaZTUl7PRi4INJJ8l4GewT4RnEebTgSBopeSaJifE+YsAmrR34sHCXY+
JlpIO2EGrj/oF1XFWx1ME1cfD/hlEH0zw6QlAETAEAlxN1aJwl1FjQbQYx5NMZozUAj9k3bn3BFQ
SbknQrDmvZ/knmsqdouN1pDsPq/pYQkALRTgpXIdnrNVGG708kStkyVf81g2Dw03FPjZzOGiBMA6
1zgiohGDeTNmBDkV306EjcIF6zTRiAbkmmQTZbrN4YUiLNqPjtAisNqrokKWkHVwAfeGiFrjPOcQ
mJHb6FnSjBG3S17LCHjmY6wb8ysHyb5+D8gHKEbfkyfpEbuE2Gu1btPkA2Hif/v+dmcJaPMBxTsI
jJvhuedwmqI5bcXUCXU5Oeq0gyYhTVy+puZotrTeZkadqpRqS4xD7S+5kvoM4HQMCHVX6U/x7fuo
P89jbn1kGJgjt94R11AZR+I7IU/eCIxLZeN69WL9TZ1aKZQYJFV/epPlCZ8gtPVi2PfsNNeRTz3k
IUVBrFzjKgSex1Wypw/IHXC3Tf2IXJ69ZV5FLNJUJJreDERERwqoCDEbxIUbYArSkuT/z8K/16Zy
KM162oq0cRYr8Ts8wvyDH9QReWMsWX1zCXkUSpZ50dQFIQSTs2NhmrcIkt8mi+MI6QYnE1eYav+V
2WMS3+9ZeQoGl8hi8gAyrycKY+vEPswzkADqMWXa/40A1xhxbDbAH4WeJBiB+0q3lNy0e3tuFHHi
/kaI3IEXmRK9eabS/L/hmAEu3hiR/zFzHd3PhiKtLBwh46IqEQoJel6SPIZiXUUGbbL6CdNFz1hI
9FSxLpsAM/+E0gqbZ4h3/N1LLq60bE8g4ajYaAY3bjm6BU6kjj7q3nvvjOdl+loqY7Dngdp2SJAA
9g1J4CjCf/0W2WURQYEn3e0H39ghQvMCrnvpEnyOnEzsmZ3kJ+eUuCqIGfs8DkWFqM1uqxt1i2FT
UqjmxrsHaX6o5HAhIwazjtvZ1VcqZSAw8qUT2dU8K28h29fg9pltcfH5uV9XOavB1xNrLKJINpEU
q6GYtcRlufQoH86rCGQ3N8l5WjmHXxr9tfeYlepGJWSSBPl8rei8sSkf6rfG41WNqibNGD34NAqH
wkwYEjq2+W5o+uAIuDrcAlOAXBF50H8+vWwIsDevf9oY3k5WWrVxqxv6wlI83/SSLITY81WoYiAK
uforbJ44u2s1A+F4mZ4uP38KZIvFSyYwSMZI7IZ76qAWEgxZ0ijOjY6s+WnyPEb37tlXOz8P1xS6
1tU2HsMgRa0KFvyP0Y5qMAQ/GHhmnzwKr8xcuBrk9rTCyfGuUYVzaU8svfeEAe13Txnf6ppvigrh
ijnxVBXTPr9rfOHLu+5Xm0i/DkHBm0R6aAjQyDAA5b7yGF1BG2tVnTHGQoA5NN9jhKVJXHujivLP
4o3+1DgecwcuepsjNjvZ7iRD9fI/BptScX/iYzByFYcJkCwGfZZ/7dFKq4fknyRUGjSKV1pkl3PO
k5MNufp69ZdUY/mhbhjgGpPuSUBqqbl1TJmChoSwMu6rW1NZGmfCPDuTdLy9ovd+x3S1Dj3uUiKD
nB71kGG8QKmYpMAs1fqZu3BnHnOcs2LYi0yq599nmEq0r9NJxpZrRE8uvcqeaBS3ehhGVqR5NXdx
ASwq7tq/Fsn1wgbupgzupfqt+QZdpLM8cn3Y6xbIvvNkH8ujOYzobp+mrgs3Vb2ugnue4IochxuH
lYtgUuisfIoXmC9vDhKYCQ9+0OwRRY21WnNcu3o0K61zF74HUL7TyiyObC/or4Ibva5hznTa3Xpb
Q/NnQL3bJyQfUtn3GEVYvLwiHCZhlkyy7f+0+WffycFsxqqHuieqUKSxnZD+RYB2aTfiG3E53nMW
A8KsGbh/8qMcVE2AbtgzdSF+K5tOwPKmamVigGHyv6T4XLrq91KAz+0E2pigSIr3dLcn+44UC5tb
FLA64EjJ3Q75WNh83UzmFHK/y71HVtYp/e5poOaWy62QJRtFYGPzJRIEbjPOQLXtWQsN8CeFEFSt
lIeTRyfkQfgwHyBxD/HJu0R2pkcTn+nyCxG5MlNr7uK5TzoNrYWXTGL0NbqWoWTp6Esbu0j/8SF+
560fWC1e7rTHbA4YJLGdzm4opDIPoOG6CX8XDG+v2qORT4pEX9HSIhtmBhqGqiYmNd8m9seAwsDO
5wgTVbZjtRmzdjNYrXrX31XWS1KYN4AT/e2j25Yne9y6IJJgYE9Xn3x211EGFvMs6NsDItfsaJbA
/6Cfz62rLnf+EfK4tfqvHKTqs7F+LOeA037/11cM6KTmgs+F0+XPqxMVJMMjMZZrEwruamoGHith
bdNNI/GrI0s0/dXQYGzPn5elsabUobdB1BxieyqcGbeA9dcVa1JF0pCh/ozyaaIZxse0dLtFQQPM
XVh7W6+KpnXX2pbzC7c7gJDUC7rLxEkNLoiaN5BOmYnb2bLFVn+Kgx8QesvG5zWT1J3/j5lxtnyR
XMsqmJoUnA4Rr4MCWEI58JvJPF9qNZKosydGad81PJxw+zoWfgWERNSaLm5p+ic6U7V4c8ldZJDM
+tUUZje8PzLThbE6mAAjJjESmYwZ0xJ+Aesu0jJT+YzebuMJ8sW4E6R2RC+v5KjYxLbMorRLX5gm
Q9DBVOJ+5zEw8xIIaybEiXzbUyaaUAaofQsP8a4uldcDxwHEf1KCjvrVYHAfdyKMAT7nUYPjCRI1
xBJQZ0Wb8pazY+f8Hj7ctrLyq07u6sz/l3rLSTawBAsiDSSuCz5hQA9k8uvck9g8Dw84CfLcVGAE
E7BWeuurBo4uExFBXSyrdSJyKoJ3uYXpDFny/SS0kp5SnElsRDf6k4hrcvtAiIN9qWfAvmMoC6tq
Fk+xPuvjSremh+6BnUHlZznUFSsfbE315kSQGMMOxTtSrUt8LDJ0z0KAJZSPd7ns6uFNboBTNYxP
UO+sKi1thL6orRoplut2+rISTpXvRzFz/Jp1DtEgI0lZFyBJic2/9MYzeOokHpaKHo3kzCJFx3Sd
vwQHsENmuOoBQOLC/00ilzvTy8pIZm2u/v3w34IvfxpXTubtJuV4yPNjCA8BK5OWYU8jrGitgtI4
96EVdnnonc4Oy0c9izOdDIAQ5/kp3UqLclp9eQsJbbZrjwwAlveWG4VNQv7miNvuUGeYO0/uewM8
Z/+c8WBhavQ/eaFGLU6YN4UiH4ltoWK9VK1kYCYtksw+axo8b0k25M8hGtx42OK9c2/42q3+XFaT
sS9+P04z76y/KwqEXaWNiXBGAYoG3CMFEc8z0h3/W5yPRgGYgE8z+CL9tqVcguDSg/ujl7aoaV1k
HheFZp+Sm5KfUOA+ZTo6F2lYoS4FHwCNfRCf+owx3Vxg3TYGY4rS7bXwVViw1S5l7QW7Rmyvxgkt
2/cthY0yfG2KKNvhxxVcRyYIZ8qDGobRljYEnqZiCaJp2unXFhbOl/kfDSDtWWIdzX5ghDcYIvw1
1e+Y6GrC4FaFEGt+BxCPycMtZyVvscjqhbTb8fgv5JiHwuKx/7zhm3fawzKlzyxytFQ8grAxLEjE
1GNz6Xz5bZw/3ldlkNQNt1uoQ5rx2SgsjsamTdAqwwSiSvrwjXExzL9FQ0a0+7HoRPSsGyt2xPLg
LygeRl/M4adb6lFFlTqivKjqCI+0dSBO06PCPMtsJ+2SbQoRZ2WT2AfBHGA5ssVE3Yu0b0CNw4ZI
mKahCR/sbau27+tIY5hBeowDCJZUaJ7x6UqeQNcqdJJXHlWZQ5E9eXmXLOU1wlTKmD8Ab9mWocwj
1DMKj42n7sqFJn75/7IbglEgsESLcKTnSzX0koHzF6tVe7mEXCbjKdnr9AUe/mkKvLheglUThShj
v3h7PMDRdsnbQ0eidyy/1nt3TtkmSntB5f12r0LPNwGdIIXVBkTw1XHxlyaq3Lkc6JDBqE/rAXdW
PVTxHS63Tb51TRGqCc10Ak3fxQu5jO63hkhgRjoLDJgz/jSNvgobdLm1YV4OmXAcZ63Tc07sqHj+
8VZGkZzRIXMPEIINP/8pQnIuvZWPgTnE/VnTEfsa8uzgcw61VkX6TdAf54FTufz958w3NCLwpx0f
YJ62xtywBiY4TiXFhlhwH10737cvssClsCVJYVqEMQuA7N/z+8TjXYidARfkVrTWM3qSvnrQcyUi
62vmYfIH0+lzFeGsaTXUOT+wVNwf1tGY+qqxViljh6HplrI5CNT/lQpMRYctHF37rtr4cHUwrNxe
g/gWeWspr0jDtKjzOXOwMIMK4JRbbX3uQvsg8qD8z6JrNyjG0Aidyfbck65rd0KyL9CsF3yB6T3H
JZKHvZ93nyOK2zdL+HT/QhonubQ2FYMgrT9lBAcCn2tj9vyUhKA5Yl9hQAI0+hiJwiAyU4HC6R38
e1g9XKZL/gsi40XF4hoG1kYAcvRyDgLy0ioMhNFDs3SzvK7sgckod34suqrmXWNBZXQG2HOFPHso
o8SQYvTAOT2H6Dd8nAjq4tGgb/ELFR9CkMRddemUqepYwLcz+4394v8AMChdODrS/VIdsDufFbt0
J9zstMBCq5Xiwaoe18vqP0jsgm4cGcn+NZaZe8LYvaW7rJ6WNydeT+kBEL1nNOMScvoa0OoPDdD3
8Lfp9spU5LM34Ug5+cwOCvMfmlMvAH+BgFArpWrSALAJ+8vA5X2uBTH5xpmWTwL5knphlFEvCVpA
AAY+NB2Fq92SMFCQKsZ8vIh51B0XV0uzuAUcrXRT/mEv363TZfwlOCyT5tzzORkDT/MYcC+KKvxR
hKyXH1YftUUd29e6iEV/7Oc+EC6UvJjEP2TFuG6qByNKxV8Gtei0yDZzDc4FIfImhEKYPO/5+wbk
csVk8xy5JhKVLfxsKQTFobBNbYYF0kgIPMaqTvEqGKCz1V/ku3VMCkoNJUx8BuDQ9II1s0I3z+u0
3WllhsjrhH4M05+PIh2XK1GTR0zWJ3VenC0RL+NFDoy4kWhFWM14KfMtP0ZezIjAAwfFpmpu5wP2
1IAPccPla0FchcbCKgAV8R6BlN7cGS7BaFAAIUph6GP78opUbb2JrpT0CLyXh0XR5ZddZ8fSu5wZ
WNkBilyw+UImw/ivF7UGzqPqHTT97cY0S8XYKwEN5LpED+YXLaZMoJg3pJOROETovEccD/1VnmlV
oM8YKMU5kDJAPkES+EhlygCklzKlzYkUAdb4/pzLUq8IMZWE1vr7Pzri8E2r6TBQeBZvHuE1wSX2
XexPLiAbt4Fic/lZg/2hlJd9mIpMZ+W+2MpfRfs01jIY/KnhqMPrAOcvaCTp3qe3JC2zbOhlvY/x
lpM6I7qKY0hv6hoBlxuCnG7uIu5xlxgOk9V8W1iny16SFpJYUoJSEjI7HNFys2cSuTxiC53hgBEb
tJ60kwhikFJBLwIuoLN/4sLeHOGrcKJvFUy2TLIDc3yFppZ+d2oGngCx7s7UaMljlJsgY6FZ61eK
qvLunByraedQg0wEx3X63IlEFGCSFvYrDYveeI1cG2KceXB/TtHBVIXKRlC3EcYJ3vCgria+ohwO
dni9MwNMwJRMZTl8X963dqfq+jeJyC+WWieLOAdRZQwnaK0tcwePrZZcSe9piVC14h60BfUck1wi
taPn2UOZZ3omzEgodrMcHvtE9xcxJRSUmRD+Cqcht0ncEVRvqg4yGHoyqdCVUPE8GervCfEIlQr9
54Ms3W1TJf1MZqrwoi2Z4RMhSBACJKaA4iLEo0pnYpavViXnIcZljy2ooH0B/IsfyHuh/cCWM4RI
25uDyXZmRXvDleRDJd0js8xksa2mLx6+0kVhfPQQNz5qph6xScKbuaZWzPonizNyoOYX3xoA+4Cq
EzmozprPSr2s5Jni5a+2Tc35g2bgAWM0cXIztHjBhRr4SjMZ8Jbezc4ZIgXcxjpHR+hVQLGDBzfn
XauegDQiIVzwnqUuuTByINDlw9tmYJc32C0UiOFRrjtzbVIF4vrCYVqXB9qrNQGFgUWeFKSp1n1z
sK6EOwfTUmr7SMzkdMlN4q7MeEzSn+kHetq5ilxChtXsyPX9H3BYNzQhafffkms23qfMt3En7/Hl
Ws8YxUZw/eSTXi3WAg721u2GyPwTR2xFpjwetYnoYYJ3zxNQiiJucX2p9glx/r25u+yHyuW45V6u
QSLCtJWxHl9tCB+nc1MJ29KcCJqKKcWBkQo5nW1suTPQWSdHErbQsuBPQLvmvjsv1CpZcVN/NDmq
9bcxQnftmVwaKBNlHEYo9yzLA9k8CYfUW7hlR0vtClLEJB/P2X31wXIGMyWqyMi7HpaSDT4xBSJQ
JO+bslyV4K1mCOWv/cvEb9RCinQkxAgyAY8jcWcYoIRAVJlvl50subZ+4nBZtknnJpRI+Dobx+9c
DPivkAKPx03PA/AmUyWDH37qXNTd2lresFHuMZqpkEkAcC7EOfntfRRxWw8p2fk/fxe4aVypCZjZ
S3qgviCApkYLtmYE8xcJjrcltQKzGbmJG9R/+wCtVznCe7u8UhQWx3dTSLeu0LJhU7SRbk+4X8Go
UxxOaQ2DUWLZFU+6kfRI/1/mnPDurGfF4BX5HWeexEJI4iLaBIRp2M+nB7ZHpAbn1sPbgwSxpTjS
1lhbmTLR0G0aRz+R1OvHYXFeU03CbWKVCXjUpmH4OA31FONSlyzNJlAVvxE33KpMUTtigJK++70w
xzrxSR9YP7wJD8PsL7HZfsqSoOjYZt6D5lMhVUprZvqS3OxZlwq76ZfN8nhp4M7CW4DLRM5F7kAE
xfOK9Et2CGVaRqBfH4DUTcsH4VBoaHgxnA1kMp5LOA3nn3D6vdbxzTwMt26jcYCvRTV23H/vbBtd
EugpLxyj/EC2v3vZrZTO2PJJ1eZgydhuhDKwa6Jo/ZBxtBhgUfCkYlaj/fnXruaeyEdz5FIBZ96n
6IL05jokGfejTWeO0DNbARHrIJs7PGyZSHNpjGRuCowL3eIv91nIkjWMzRCm5GnEnwRvOyVWJC9F
cTUMwS6x6DAc6BZxHarku25tCZfJtJyahOkvEQ62rsMplMF6IPIAEbV8Ej9epcbSbR4Dspe2AHPh
Jhfc52VTVBwhjhW0Hoc7T6mdKE3DRppCOKT6HJOMIrrYI9rJR8GMDnYilsOV7dibf+QFszFqj0/+
x0E6hq43Le7mOqDHXoUpHSw6DL5++YXVCQfw7QeB/AqDcrCPLB64UU3l0SmCLlow3VZeyD+hX2uj
Qw7b75igUaSZ0m1YjytK7gUCY+iwQbzyg5KqAMQ9kiscbkFM90KKcgzb8OioN7cYLR8NugpuTPwd
1895rBc8+/OGhQ97s5lBlPJiTPNfn80rMsUV6smE1Grsuo22TIChzCc15Pr5hsH/dvFPEr5h4q4K
cN915MrgRLsJEGi3PFVgFTI5KO/6f2YhdUW/xCrrH/JgRRUf5Qhz5omOCBHh6Zztvs0Y8hnBemSN
aUIcAKm/7+UQ3p0mzQVwOj5ipg2Ln9/M6qcbZnQgMiwYH/INOHhRAZVl7d9DVOUtuHi5pOjr7OuD
c5Ikq5L1BzzSnePvtdtElQDmQODoX26+ycbC3zBI2GHO9zOBKIb0oslWQ7cVAk4164fJGyc5tbQG
rv/QcxP5ROoewiMWjcXbqo/6GMGvMMY3zSCRBuPhd3WuQpT0aZ2D5zyCSVp7p69Q+kN/FN8ynaMA
bqjexfejl7oEOBhJwfvUg3h3+HV+92eZhBwyrmFtCAurvbiBYEi0ZmZhSlIF9PFlhD8DJzFza6BN
zzD8/uEk+7ql0eTlkQTvgf/QyLU+Gj4WOHi6ACqfhNlkQbED3MXkxagYKS+ybF38T9dZu3DJgNso
ByqSXD8n5KthWDfgSgGcW//7qy90/P/VASS8steGeOwPbvrlSVAMX/ntyj//Ur72yBKZBVB1
`protect end_protected
