

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qbCebIw2n8+gN2UzOmh7axnoM4dwT2xHCHsKSFB0KAVTaTY3VeBTwlUpMviyYkfKO23wp8O7SpGs
0Wn95oRYAQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MOTbFTv/+AMs8CgHaCOhzDGjJY2CXbGvrGa3rJLL400WolIwHStE0ZS9HCf5QwC/qlTKHtSKXPFo
IKgluTeQifTssmpfL3kRH0S67h8DFhFcVbDg7MudxUvt52DgkYpYAzVfSG/nUYQr0UoPZOGdWNek
d5BNE54QoixjvjzvCn0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GWCTcTUIemqhsdR62OeZRXGpfrf7+14v/PYnlQE2+elD/5AQSNezw8Yh5LK7/U0UILMPApnh3/AH
E8gsLq5Dk9JFecIp+TrRarBrPzdkLyp/yDQZefDHIVKK2//cPrCux9IXp+jQExTJ/wMgB3Pk/8bX
EXcTuij9bNakvhh0qqcvPXbXX9LL1qrTKljruNhZ8fj+nzA6ZReUIHP58Y7Ee1d3Xsop4p9lwil6
6qwN+Lhx0npqK6UrnqNlAIb5F4pmCfRi3mvh8/WO2vx/mksFcUOTOjcUSOA9S4Cc2fWFZaEJu2Jk
nSdbTDU9JPBBG1HOZLBI4PeIS07u4kvjL8YxuA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWqfi4eW93XaurdUTFdBvYmgRlNt3IP2HZZVV3EH4zpzhLtjfG9ITAAZ2wgVBZ/ubHVDQNx+f74V
7yqRHt9FI2nIXks1MGER0/CZXcSrokzmAY5FFnm9jVBaptM3nivib//wb+pTYDyqkgJnA/Lik/xE
5N+mBusMskQJf94X2yznI3BP0RzkvftwacL0/QByYbp8e6B4oEzsoFkwinZKNJ2vNWKLPcxUvmlb
PGne9+10W8+J83DqAyg/K8zGYWdHwirFkQalIXh13D6lOtBVr0AzGpUUavift5/tIqjagi8Vba05
wcVi1W96tvqzhLckg0QwF4ZrgLFtGXEYBLEWwA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T2Je2NpQz222u+FkFMUb+rWAcPEE4CQIHwQeLw0xXMrIAVVpaq5m32NeZx1nQkTHVHeERS6BRWqE
5KXKZ5QH/IVcY6HLPbXO3Dm2EHobkpU16emyCApLCsUgcmA/MRWQ1gDfMjS3AeaVHULoQYQW5w5d
K0sQnMkknyB54GHQXbQ9LDcdo6L8t0/QgEyTJQzA+Bh1kz6FgmgpxVnJ2LlXH2CxQ9jph4sAcht8
4D4AliecDgulrafA2JbdAEK/+S1BpiG4ACtXDtpGUomy9jKwXZ35RlimisNF6bqfSQIV4R/H0ItO
J5XFboxTqNvqI4emJgnLzw49Fg7ZKbuwP+cntw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eAGLDWmORjuQiifMQjmPS2N5D50nOZvLtva+eMzhWZqeQDnHdoI+D/Z7CnebSoJv86oC3voi3uQO
SxQ9InTJFQxtvUyucyRaLG3IUGvvgRJVL9/LE3scUCA2tTEFitvwjYXYvUghUxVeN0l5sMqzky5n
zjDXmH8VKNGD/5c9uPE=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HEgtpre6H4t2Ov3YueDpHwa/86EaHsc4/+NjKCU7D9Yxbmaq3EsfTvD4TQrIFaVgkWk0x47Z+GXZ
XP5UWE6u3RBO1x/Mh6hoOs07p3vW8f4+CpkxsVphw/PlJLMA6ViCtY1RT/gVyW3EMzdsWyMhYd0a
eBNyTGx/qVPHDSwhb68iLOncdRos4xvixfgQDHKuQsNL+3IolnroIGIVLQcbMlcya/UeqXPqMG2Q
D34oUJHsZe9pFr0sH47g3KLSIk5+85C9v/KjDCDxxt+J5rehkZYhGiFA7BCW9XzXHBd3bdOzeYwe
44cUn3Y1z5xJtLKPPWZMYlyJ9qCWupZE5Vsg3g==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pKyysRDfDRq2uWj2DY9SyBumhMt32UbCuydjdoIBXHnCxoa9K8W0tPBijFY7TxWwxjCKsAj+kEvj
VtrLvHtrCvuITfo+5kyizBYnGecsUq76gq1jiH7ibthaaoTsSZdz/yX2qho4AswTYeBrNIFRKKMe
ytaGu4E3+UdZJ5AmlC2hS9L3lKp0rYpW7/3ga79U0NGN3PYu4ctIQY/piPLQqm3mLXgYEwlLSYSH
bF6Qetk8JiduocsQ5wCC6ymA1HmnZVZWWMFWqekwyt6poHD5G1+Kc09rJ1xRCleye9m4OKUo6xJs
EyY5+aaPBaQftq1EZopQmHLf2tg/+2D1daktcg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
0kwUHTB2FgSqrVdqcfRInU5qfdGwJsBIGkz8ldTK+KTBBraYQ/GLGBwrrM4sfxehGpguuDv62X6J
lPMTE8nMi6G9ce/v78YSYpeI7q/ZeUmUe8eAPmiP1OmvXq407cWk4oBHLriD8O9hefFuXKZritGv
cu/Uo8qnLtKvWjb6FEecS2BD5aRnHE5tYxenNnGfRgSJ5UWwzT9IL7NaiAm7ub5Y/ddtW8z8HPZ3
rYoQ6uunxJ2vn1Ssq+J8/Kr2eX0e5rYXvV8pd/vj9LYUEcgGSefGsnUNyANwNdqGG58LTW/DXok1
Glnp2jXB2+rvdwoOiUfSjwWfT9+YBjNK1XibuyD57hpZ3fqNNkNdwOkvTpeCY9ScZsmWioS/XpIe
ioKfcwgVC8UvrSnAT6jZtf23tXUQ3vMF9aIennUihuhrrFttBFwCq5QFgD++rGkmRe177MwbGyYL
1uGPWJeQuUwvB2Dsk3fA+Xg5yuMy72geWQnhoMkVqY9aDRPLvbY4lblGlkWUv5lMt+6g7sP7yTaI
nZqbnlvaYHcOf1Ehfca8kxrLM/dgZ+D/MW3o4lGJ4lc77hN5gTZWAOCAXtwm3N9C59IJGX+PfF0O
odR/0jDXtYlct8BapuLnl864SgfWpUymBAVEJrjuyCxzHG6uZEpTQPNbIIHdtTvb4YJmtDfmVH2f
ZCc9lNBkT0tymWy2RuyPMFddC9q9hGNgrNh/HwymEEZuFj4cFGrtkorLtwn8js7sz5L45MYAyNXl
MW0bNN0ON+DkfGa1ZHybACo5J7XKCS9WPaMeD4ai4XUKFLLVISYX3MjWIGJhb57pQwl5S7zfpnyd
mkhm6nuXykXo09EGzEawLXQHRfIyp3MjF0pJ3JEsbs5xQkDIXX3xbjI29+vUPrklURRbsNUFGA4Y
AHOx05UMPQ+vtsV5ClBx2WJkKyQn+qtqWr/TFAyuQEFtmhn0S06X9aK4AKP1C5chmCDf5aeZT4Z8
nnrYFUAbkkQj7iaU5LRv5Frq31kQiaBcl/PkLXX7WxIFWhM/ebuqEvmn6kBUyJ9RjS0TK2p2r+uc
QNlEvwM1hVQbFxxdMZCaEmS06enENzbOxsySl9PFdh0ZebVPsxrolz7Xh9tmmaUjgj7g8CYlQ+JR
SYowhEKwSwsE/AMKHHQVnKy/KJF3CwSASR2Gf/edEuQz0lg58DI6k+ZyCd1OZ0+UO4vgRgv2/ZWG
k5cLI0W2En3FVpS0FnX0myg+Ybus87A+shENzehAWJCo9LbQt05D7guR/2LzCzPB96MaBZM8C12q
gmT+dyjLD7cn87wCEwp4V6rQOGp/3IfUtxCxdwhJMaD6HGFivbRwE13EegPDqerSR4fD8r5QF/bE
t+v1LxOqIHzFa4SA7j+ByoV3vZWxtPk6eGLdYK/NURLHV9VRvx67lawXaZXfmMOcFL4NbbI27M2k
IXxtt8DRj3rUrxFuemlJILC1240k4vLmAej68Gm1sbji1FFRYHJYWqYBCQhR68UGbLH9F0vedHcO
KgKxhnBgl6lV0kiaDiRi3+A02ydtYVgW2dED/OrEjyZI4WcQ/8nV4WN3J01cCnksRWptYvP3YiYf
H0dX8KNXJHB9NirJsONxNjiO3iCOP1T/bP9B3GjVdWdmXKfs3JpFq/bSZfTHB8vz55I0fj/ki73+
96AvMMVL6nXVbWfDuklY+TOjGw/fIN2092Kitu5iiN9S8XR+wXZqAf0sJupMDlJlzNLcMxnnh8f6
QjvTbEGse1Wu4iE0Zn5YphD98rO8D3gXx/WhUBGSBFAyVZNiK3Kso2BlNO9VYQezpIRPxNeGABcR
08HmNDSaNtDB3uNwfIvZwmmXVd7j0gyQB+Kn6PWnj7Feszc3f2BiHNdRf6IfxMf6laceu0R9BEaA
FBpZA3V0NNI0YzfufQiLVhlcqetxTX30blNCO4MTeKmpYXSkZg6tX2cUwPvAcrDFB/uAkA9j6k7g
29xZztdBTJKz6pI52g2jhkU8UBmcmqmynP7VLE0SEwMmLVehDW4GIHJB0HdY2sSnfidOphPxvD1o
wTvSdtYOyUBhx1N+X1qFOq1SSeVgUatVAPOJuOplS9DKOK/ig5g+U7YoscDfaCpQSOzKHEJ2gypE
3/lEX90MR1AVQZUEnzuG1ex5FeCBkT250Iq7bjaaaUK9/1rp0gMvUNEwRmAFE7+8NLgbygblCtvC
MJKINfRlwEQPAAHiJWj2dnr2dhb6nxAqhk5qjdAF684yyagvP7dASp4iCVbtlAC4b+eplOEaMuMR
1jmwmzOhrE8oplcVjPM+B0TaoZrjGItRqQXKbP/nNnUUHOa4PFRVtToltB6H6MJkAECuCOvN6a8Z
f2CQosEABRwh3Tq47/NBw5DUT/zEniVdTNZwVJK2KqxbTDg0/Rsp5Ft77yYGm8NL6AJbRyeXf9LZ
BD2/X7qlDAXIXS7IaMHwlDN/Dfw4mWKBjSJaXk1O1pner/dmwOm2YJrskI4pTDBMrcGzqryclgvc
ljHD6wTMX/hJU19HSfydEI6MYzQ4C59OiKBgzC1bDaFzAXnQAxEL8VKRyHtt2k0T5HaH6y7uSfsm
UYXgJZv7v08OfDc6SgzYipoqK0dOC3u6INJahTFVZ3+nseVBPaIE6z3G6HeJQwL8p8xmpfrwYV3D
7qAtPjE6pTn5W72ZLUhL1e0itsMNmIg3blQ7jA/4PvusOnkjaeh5YMwHEjVQvh6rd1jvZgoLD0Y9
QfoREUxyCpKCpyPJhyfmUwZVRPakFz8ehU62ko3RltKURmdDprDx7KsU3S+O9sYCXNe1GrRUpGH/
EgSD0WSviN33K6z6tSnjXSjRxMQH0loQobCUlEp+jWIjRRhXnwzK3QhFGzsee1WHYu7aF2+KDxZ6
M1kC5T3F2MSTfVUwsD8K8UsK13l7G/LaRxyp4+8j7lTq9gfqjyfKfEuR5xvGXKCWGrs9GZDbNZL9
aNA9dtnNSz/74TEF3bdiNa4GL/BjWUsE1HhZ4tE163iUUedkS7ZI8Ei/C1Jgn33WtQ8VbX52thJo
ZxOYVQZ9/heLgtgloyeUs4lI2uWQdIavKe0nuCqBcP4p/A3dcNJC7sxpzBlgXnTD5ds7pXCFG/Ri
P1a4KmGS7zRuuit/MU1gCJRpXIfcQVADJV0XaW0CoLBxCBkimxWb/C3efbC9FgHsJAR5k24WKb6L
0zFN/mVAZ1koG1ONtnDjPiUwEn89/OptOvR4p23+90EHYVsCDdPtKHzSAt1N4HU70/EvVNXJeGxa
oxgYGRuY2kgbE3YUBI+kn9v0I1cHAh11YcYBgU3oIcPXISdTBZ7K2l5VIKs6cKPLdgIlCm16v0d1
ZFXKB6xq1CEZL2t+myXZiqX7tCNmTigQ8DCNaiTvpAVLFbt8NeuTinoq4ExYHAjJnlNpyyQwnU3d
+kzN8kLCtqnHsr3SgJ7VXFQPfzRM4L1He2mhcFpgnoSeloA+rpcmw66mWQdlcUKPpKiVdrRbgiAd
sC10w/NAiMNKURS7Dz3d6WqqSF8U5aOk5Ns9HoGWWBwmxjuljCdY01AsPMHQBRwHB7sbPS4lVr/F
W87OzhIneiDzRIl/12dH+iDj1ChdBEAjvOgxRmvESpbo2An7rIP2PkMBn8r1LDcDkPQesgDruJkw
3wbNdeARduHFtZXWD3Y/4PRz8EAUoTpeyPjeC4iz+Q7a2RzMEh2Dm+DyjQdJhlvj56sJASTmN4uE
QcGYssezeKtObQjBMDziyC5Q9I5dPd5KYVRzr+iiDlW6owPB59vIIG5cS7e8/5cwCiY7cqFu00Pg
L/6j1z/wh6CVDcSXCwNREXB5RQ6/G2e4WQCQAXgodWVQZxlOWUm0ksDbrKhu4C4CX3VG7WMCGNUz
cjg5/V2zm5cdy5TtcV1f4qnshl4phPc00rKNH39kMNshC7QtJhUthrqcoAZ+sdCyg4pkSboKmYTq
tB2/AZkkNA+iwKbsPgbdZOha5dxBrrli+jgxa5H65W7Ha5cuETSLnfPRUtJ7RFcaiMg6awLQo8gt
6sZAKQQp2Ra9xDOR/rzVX85F+BqSi2sQUdec+P9nO0yBSiWeGSf9p2FVu33WomuNUt86cTtYO+8J
iaIg1uoCNOxsqHruNtUtyMHPkDGHpcOEdJJZURyOVnzHbK8f/Ppk/1+i2YV08N94Qzh4dbvJfkCT
aTQxuRA104tU2pbrDuRfFZVutY6Khz4OBmuJ+hscgw7tY6xnuKABguLsucjsRAr1kmPSccehnmyh
m0n03AE8ThfZH8zbqh0/y/Z4vU+QoxQJwZawJWIMfFLHx6m3tsSfG8+GmOQBGtSbtZpT3pDpJR0N
nIhO6Hc0Ep/L4dI88XH/cVDavh1+fzHtIQOXB90Wl0cN6fvxeRoh3eqJ8owBm1jiS5vfj7VKhY6b
VVmBBuUGyF3x9Fdrz1cubGa2huNIBbJ/Ip7N0zDcOo06qji7xltuVuUjDb9eEJ5iJ6ayA4OJGV8n
3S96VCYHudIeljsL7fhWkcuXo7dACJWaysI9AwN9iHh+4b7DMeIaWeDg2/xO+Uu6EYjP094sFlTx
CCW0VnMjgkoPyWFBIUtJf/g1W6h+kwaa/j9ENDC5y9qPGkc6LFVRWIstY7SoEUXHfOHFIQD6mYPV
vRJ5AFE7EQ1EgoPKZoeWpXTnCc+SyfTLrsLXCivqwknvO2uz+xxgwmlj1rNleuokCGmNpucxmNUO
8rfcOY1e+s/hcnMVrmF4cQX9zydje9xx40cYHmsdF74jp52gJCPC0C3SiEwDI18ZLuEMkJfQfR3K
JXAIDYHSOeH4w6SMMVkNOVWOy67s/g3/sCOD7Z8vfSYK0UYT+K1kroHLskTmPL3+7giygmV9RlUl
iU6AOKR7UtnckzEiloCsXgwZKVkOzPxNZcW/L8JHmrX8efkY79ebKxyTT1NohEMx2JqtS1sEN7My
mqWz0fLPTydOXffqXXCKPnLUJfGS7Q/zm755XQ79hQUv0CJ8XzJIHCQEr3xGVlxOBYa+upTKwwSr
WZTy7MNs7LZk/m5t8e1PeD9aXMViSeBy1E9/a1UxvTsskDgmjnzZC1J32FVS2mIyRA7bwf/+t/fQ
+yUxom0iWN0pqECjGVZu2lIGgSqhcjbWJ+oiLxALt4sMyPL532piskLJqCCDYBQHDFjfmeghqBie
WzCTall0Qh7b0Mq12xDtXc0zpTTR9vcLeWRhGQaMSzqyfbQnc76ysVVqfID6ExSPpkbxgsSNH6Ql
t/HyK+N6oDGAFdhAKvCxxrzRH5gd2uDWHCyU3CLuwZz2PR5ircEaMrtUBLPGviKa8PjxjC8+sg2C
bBw/ozMTNCXXuCYjOpu3gsGaEWTZXN/tBsu9HCMMhkQlTrxq3vhoOteAWRCdlfEMfNj7W8EMlCom
/aJyulvVJ8st3Y/gLb/8q+n7macKF5jU7jZoDwvFNversQTS/u7S6r5h5NeavnR5Tc7b8/dZI3cc
O4QR3MtJhgaK3L9N2soTMp3PMT9qn9JucP0VCRtiMJEC0Y4dJFBXC15TVc9vL7KV7jl//mNJXGsP
xYHT5G8kchzhL/6A05GGDcd22LBTcgJevqYr7nzoAvPo2Osz5hlpfOWgJ4Pbvdb8Y+BO+fQpprrQ
QDWPl4LprMsdVdQ/YikjNxanWM8zze12zTvXbqhrDiXPShJjK3ClQgdoojrPzJLiRrIQpthPLhX6
UziGNoiGTc2ahWEnZAM72pYjIWxHhH/5r3rLsyUAmf3AQEmN43V1mQ+HYwB0HxBV3wFluId3iuS/
/X7TBC13XoHBmlP3Vqtls9La4N5RjLncNUhK5EO8sp7mAeu87qyoqg2i7t5MYUd9gp2MlDNyyFq8
KiUz9LOvbIYt1Koe81+xJOFXuzAeMAEbIhD0IAUHlgL/zw2bX78MTaMCKzN+vdAYvky8k44EOt7A
ZHSIV0v7CJdFrg8Jm2p1k3xqHA0JWCA+hHQQJf+ZSWOUEZNS1+/LsGp00aa7/RfVx4yX6+6GtDQm
ueUPR7yLp5eexOgOR9VXaEV294+mlbDN31sgxfaxSJtVkGzqXeXkeVZMEfO+x8sq+JaztUxvQ2ln
DCQlNi+FWU8RgKBgrJRxNaIvWHg1nsrKkcAgxWHp7U/9CcYSwtUsRTB82Omtym+jJBTc1CQE0tqD
klMnnPaDZ0PiBz4FsUUpRRPIQ7WFwBTJ4jxuRlXkC9X+xWyIXc5FiCzw68vzCg+b6sy1TxG1CWiv
E8UjH6Jref+UVUsT14KyqPM1xz3QjMcFS/JZJaugkPhqhDIVA7j3xW0yeaxFxKc+NlGGjwB4IyN/
ZU7BOmgKqLu0IZbHHqOJwcFumGps1U6eSeSPBV8LYhqLuOu+gabllVvYaOZGTBZ6rcvIZgvhU0Ic
Qv/7CIfYk2upqn784lv3hkn0NpIhfnp2c5yM/ZodeHYWgThkCPMxmaZ8kEtXl1lX6qmcd0WFZbJn
sQmQiCwBV4XHtqaVoULIJTY7vGnodLpXFdPR4mH3iFPnbOoOyRrnwm/3bEw/98cnMbt6ekHsv2bQ
Dxn0VC8UcdWAk/ohnX5GRkfDRF4dqKWXvmrnIpbDtuNBi7DeMFzZA1lNiKk3FVK8N4KAkzeiwp4G
P4xPvBzjZeoFC8l5bUmz2FX70jpOql4tvgNGjvrM9BWeEyCu5sAAOAIAe/h5ZtD0DFSn5jwEPG+S
SDsc9d3MHuk9wrFra1n5aC7aCfa4HoFOenK3IvrHvrxIfiowMpbjwqeA492wL/diLV72/TFrMwqW
vZvrOaTLAmAhw8ebMbn8NHjkczQiJjSRBWoPkWdNcDGIcfBRzhKUO6VuwznHF50OgZRu+shh8c69
jYifEUXpMWtfPA6knNmtFB4xxWPm1wdRXeYHF+0b2VYZCrLOehFY1BT9A83YxjKnFbPQ5vkKaMEc
Bx5ndRC2iQ9std53vEKqnd97QFZh1mZ/WrIwwPuxUgr7g4HPCTKScOLL0Jdp11AtjYn6R10lx741
eU2rnP/jb2J4jzyhJDUMb7GkoK2QfSZ5S8Ih/27NwCYbSOhu8a7TRSmVJdtCyj1DN0QVUFEPq3Yc
dKfnVUtDkM7oC1m5zs7TvzANi8Ah2cP8Uari+IGLvRPBlXNdGbbvkpR5G6b5hAPt0jF2WPZ+ASe8
f6L9U/9xUD/B6HTYXbmtRK/ruvFKB9Pats/U9SXSHZEvHEilc/E1nR3SaSUzlePw4iyh/1RAGHbh
OgvqdaRFEAPOadDYUbwk6hx/MSwrLrgqVLxyWJmhKaK1/jlQMqiEY3/IPI4Le/iu9ZAJCqpLohFB
NiAWEiCunNdYT5a14TCTybOjtAbd8ASPGrztbStNsxI7j8hRQXc4N22v1K0F1v1bNYbtfQweZp+v
VNfOgf7n6R2FklqI8THg4cXEThJxHjlZE3vdDSO6aaGZ21uticL6HQvi6Mx+V1qcfZYzsHsU4XJW
Hh6hRb+8x6NgPOAQfAuZtpFXQDyXgSXtEQ9YZrIamADjGGDKZyxFxSGQYjBXttnfWxgOUkOsHkC8
us1cIGpcmVIdw2tB/xeYAUDTHKzzp9WQAkbs376zNkQVGGN6zr15ky+oIpevppdqa/M0ZYXStRNv
7KDX3XTNd8JwZnXHLQ5+uBcra8AzxCXzvwnh4Fq1isLSrJAiQDvZ6XcBZZQzQmN6oHRcgjTYHAmW
y/nwB9fkHMnbDgwsn9Nd+FbbAkdvYwMy0HxWq60d4q3jUtzxvDJSZRzA83XbbZUX+BXLbJwoppC+
n8aTqrbIi9yx4SnjTdWYsmsSbvjdOu7KL5knKKfoEWtHmF8LfiGAaBUdeEFV1hq2w9Xz+75QSTML
SRugWQPT2I8mo4ge4XQOaNP/NS8H6qu3zvQfsTWQYXbWiydbESOekNlD3i16jDFILnCEcEzVFgzp
JhNYzWYsOHu6+ghEvHCjgTC8YOQM5EABjSuIwcc0AJeIu/1upmxRyJSgDbds3d3lIHEbyZIOzIVh
0iFXC1TVTaQkhbXGm0Uzd+9zfqdwloh/NeB5k1FIY8gx4YGvY4clQUANe1ZFXi2lKDaUQPS/fKwl
61kVh55QdCueulzmRm8eKolTQ6nWKYy/XUKfxU7chJdNpG4lEm4AVH4DcQ0b6KxF/qINKTaQQ0e2
GnXy0MbeaHsB8B9HO4wGVDHD/lKm03ofNF69uFj8ZCc8N1ByZg96SUhrX0fZ19e8TEJ1PEbws5HS
Hh/NOjTDyCBUephlsH6OlUvja7H4aXWNDNbCX0oJ65I8iaCVMYzIMrasa5ineam2pNgvvUQZB22x
6cuHd0jjV8ZXi9Gw38FbDEQw8OIHUVMa3uvL/a/1Ne4i3M4IPxvoGkBrXvX5oBnj0LNzDpSJw5hc
av+bAYNBq6IEG2ccZVv0JtnBs1opBnDP9ik7R1wKURtIqAKIBPjFDu631dxhvtMgjkDs4iB7RM2R
mFmzcLmQnGZnMRgUE5AB2em2B0+aWfYiPaR7PQHG0eNn9irMFGeoLvhVqZysb58xtxV4KhjVXXuF
gsWTrsLAKsuRPrErsfJBml+dhUYAQWeyO/soVx8UQFNj0fy63Aa2RXvtUL4+yD1vmkVX3HDTt1RL
VBgwTIRTjMho0NZyYvxjRE3oTWiJKI4LuHXKA0QDdc7H0rVLJ535aZpyZp03hrQbPvIyHqD0JFpg
iKdlKgwhfDaaS9kBrWixSuCIwJQlPZ7QIDj5Lo8zJ0iwcvG1s/BrZ4RB0gqf9VisGG7JRx1JRdT/
vyPClmTQYbKbchMGKcDAnLc42g/FO8QBtqRBsuQ2ExPVAkQEo5PS4zm1Cqdx1oX61cbFAGiXuoqq
4tCgFeVs4cUudI3gjJ9hI0rsLByOy9xTL7lioKqqmSJizedaHDNnPfX6+afzEAnThiCph/0+d/sp
HKFiZu0wRBHmj3H9qhdSihUbCyetQzAJDmdCIY9CMRwnrDVRJ3o+sfBpqD1esiOKDbCCrDkNFpfI
RDaY5Z/oatRRaZgJBp7gg5fLRYf48VCZgkV9Zi5m7xC+cVFwIN1IuNJdryd5mHo2ZzmFvkiZ7Ao+
EaThJL6h4NA9C/NK7PrSRl4+5ud4eawBSSoFRCCsxuimEf4jiD3/kmESfZY88GCmOI5tXL0zdkvm
UhYN7QfLuzDyX7+NV0OQDdzP6IuTtNgGgvuBEDg9e+KTOLnO0r/sOPlJ4/7p+bYV+eFoiz04TlYN
o2jvsR4hL7d5NutuwN474PCyK20cKq2mzcduCUDCGp/C9VovNyw+OIuS3afB4gGO7PW4QcE3SaV2
C2VbVKeqI014s9uxk6QGcmTU5iRYnmj+U6zFOgMKL031uRHKL4HyadDSDGczv0k/4bYYM7Lx4CQc
xH4BfGFUeoNYSLFF3KuSIfZg65rXVVHmOgkDx3thCeYN4V0jOVk1/cIrWllTdQdvv5ZFrzJNYMXP
ULx+tJT/fG+Oa36FriGDJIW0C7qQuBCCokdwTcE1ZbOt8wJMAXYFrt+16Xc8ceoywZ4t7UghbMkR
ectjYsJKBzuXspB5ZSSNSNQ2jIxK2sIkMIJEPjSR+bHwlKfWjHC/2ag1Cg2fZzz2SrI50Ag5lcJ2
4Bi3XrsghHJ51VFljQwbaAnpBQXzt08J6jzBjRPfohGmv9pQekxGIvDCW2IeQf4gsqEZWRdarYXu
VSMRJ/Rjj5MlVunWviU+VGCFFYosD0D+1Fd/ScnWjP+4pXQAFE/9nNAUqrf+NuDKJDY2tMQB2smJ
UPgqfaphiXSKJODr/v2Ip/Lpm7oiCVZtqeR3b+Cy5+ndO/BvJBzjjIil7KBbw5hI8B8O0yv1nQ6p
5lo80e8WUhCC6D665uxacNzuRkt/zCEuKoKkxWYU5iwt2krtxBawhiojA2IoN42Xu6HzyWkqjUAF
tvmtbd9F1tBLdkFv1NUkU4g7No9p1gmkqt07999x/eSmAtsEAf9J2glhj01oLCBL/+h5tILy8Tt7
lNwTF4+fWBG2z8/fzMWakpAIK/NH07zweJxSKz8sH+wOQMziukzbhzLbdEU3kRjXtTHgmTS3RXhp
44xqGxeD6xatYNoeVo1J+KYayefansDXO+loppXfzOF2ueGgCZXuY/EE9trs2Sfy0cQAKx94zwlo
7Y4CpdmW2MO6AtolLthFBVOJLwBW5fMrmdSDFODjHN5Trg4ByWQlAHFW2jEnSVRRaysX62QO2YPA
1SFZPWPOnViFXgl1mqThADzaPHyfGu1/wtj+fnq3kF1/mfbHVDYinuH4llX5OAtSSUXBcSc/hqke
pL9BNMHRkeKPdcaKuD/OYR3aV7NT7FXgD/XJftC/wnbabM1yZ7rZmrQwMawtYzHDoM6SXCKLUEq7
CguzdiZ9DpC8vSo2h1jCg1wIeRLMMxXISdbER+/Aik0G9tijIun9xEGKBjL7YmMvuc3xNC912O59
OeMHYOQInlyH7Gnkjegs8RxlywZLrMhx6dFaorLW+QvsClq7GYGUtq1w/WIzxeoNtSp+pnZgk4AQ
p19gacbT5D+4qKKF6uWnnCRE48nBiahdPdOAToDk7Z71RkMYHNyTqX2Ey2PPUmUHZwJtfpg3OXg4
CkNZ2DNOsVVFSRJfd6AtspOVK+Yss7l6Wvnc4B0a1UOTIj8O6cciqvMBvWDLRfciHYxCkgcqh2Z6
q8VbS58KwFyNim5nlbxn1cr4rWTZNRuyl7JzM8BGPzaMrTzxqdZO+szib7SG7aKZLTVs7hR6pYfC
BYZcAn7CTCF3/rtzNVSu9SAM6F2/WDdX4lwfRQ/02LN7zS77KhG0PClWZSdwW6nk7o09CDKA7a8v
VfOsBexgFhMdI6MYzw1TvqQ76hPdJyX+fRVUYKbQ2ouggTy1jCpRJFsEgp2StmXCzhoDok5GVj7s
DQ2cVFJ1Nosq9mPwaDAQ8rZ7iHnPg8p2Ip2TrFokbKQvxq+nEzIa9vK38wRW3Cpc4lRXYIPGeoOF
E6WiSSh0xn4zzzSU8LuwSKSUSyr7zr9KWKNSFvffMTgmdARyWw1kXR4CEsJtUv7syFRe1YFXAmBT
fsUP2re5FPCiH6uDpdMYpEt12VO80zeiekdtb4oRpAJ+d8cpuWMJgJHSbe9KylykeLLDEbqDw2wD
6IcoruaXVc0aKW/hvxBIdegvl/+rCuAGo6xhl3g7PaVH2OnuxERxeVcAIeeDQW6+wt3LpEx3rGyf
FdL1VT9MloyQ2/vljeMJQq2BxzyJnKmxAeQjJPlR7c7ZrzzQj+JO1h13pgyFaJ7g94uOYLizPE9+
fFCVKkSdTOHFBJyirgV3KOAASrHuAlJEXkZM9UwM8NJuG1l+pCHjpSiDieWXSn+T+jY+RgBuZReJ
AaSIXZyDN9Qj82uyz6yRls7Nutii+11AOJXTRlacsUis398v4ikk5VLta5fkrzCG3qniD6UdYvJm
2a9w2H1ut3QxUAyMCiN5ogTRSwcoiD2vZNm7dscCbTg/bjD0XXNNMgGjLYAodYCO4W3waqf9ZZGC
1M6QQo9jPGsAN43eetwVN4rw+ZZ4RkNgD4v/N/pR6/pvX2rR9HqqeI1GF3sn/OHQj1qTSY8muK/x
1KIztKZ+TECaEgp9E7ZqiDVfBfs3lx34DahXhGJxJoQv+Hzvpa9TGCJQhw8FvlmCes4XmjFGsuZm
otsTpAg5cto+Sh2jKofQ8bpv+ZhhV7/GNcvOAXmdc91A5LtYdJFyZCReZYSZSmXYr/aNnldlYqLH
4csZy7aW8yvvxXmTSKGUXDreom9pe87mi31i/5UpwK5pCzWtIUpZjucXOPBwLJaVf9qFYD7dd/YI
VWvW/JQVQaSNCCjSQUr2b3vJtq3gn45rVOZAttfSJLMMM476HeJ0kfrnrGNYj8sXE8EKN1mXvSi/
ajwIXqvG9G6XKuBtH0XG6FCCZO7FS6+BmOTP7B83FyVGS1WenjbydaAWTB5SykhFRJG0HrIE9krn
PmaeL4jAOZcaI56dMB1bRZmtolIfkVBlNX1rizkuubgMRyV+2o2IuAOs69kCH0XrZdilzyUunXRN
vRN8vDpkIX8W8MKSljd2v386HXxPGFxS9gOeS22zAyQV7Fcot6OuIQ2fpdoYR0nX+iodmS9KMmn0
lFu1gBEY4S5cNZUlB7NTk6G9zuKYj2Y/097dOYlla7Lq08sP/J1sl9IKLMKW0Hn+SAkF1MjUzl7I
nOVjNkIYhZK4Y3tMiAhP7vvYFGLkRjl9BVKJzPKcJIkgqHJPoKePkoJr7eD8paxeKsiukV/Sbi3N
XXAKhP4hNU1rgv6mWebRgORQ24AHIhnoe1hH4HQUYk+PtgyjpEuq7dL5TVNsa5AbPEPVdI929eFp
pTIEmctLf7sgz3GdCU/KkpD1jWFxlP8/vQxL5tjmlk08zBnUPx0nF6DOz6QF8IcDMvNa15L5uOzy
8wJapLENKoTymvWY+dYbMNPsuYAJwnRByKQlkDL259Xnu+z2GOZE61RKY2TV4ppTej6ZuOlAEKoN
YZqPotH8L8+lr5fo46UYrk/K3cevDR3j2uZJg51KWFCl/IqCrW5xz5DRc5RPwHNqIDDVfkrmTk8L
alJy6zEFyZO2EBPPZqbnPJ65uowhz7dU3uhJNU3N6Yhea010iLtso4tnIrcrmTf5O5k2mHmjsMah
pus9525P4s9/KSOkJAewSHqt888duX50WUlIXBV5R/dPPAeXF/1VaNuVQ17xVgY+KAWF8SeuoOZU
OFU9rRtiR/JetfLXCI66WvTpMBX7QeSmzi/ZCYJGu7bUclhJiMIWWt33r1gV9eGoKyZZdaozNspI
chX+RbwUW76bZnueSgJsv4YEqjvX9kuo6Fae0u1qGaX8WKZGpP0oxlPIikyZYPywdQr4gEQUtvue
qgCQ+3DJW2/3qBn2fb8gUWaM1KY4YLLvNw1oj5+8xjVGbgUIh8QMd07Ba1HSXOBnlrKrhyz60Fmo
oV8tgh6wIpdKgH4rSPrGwJ8rVzA4lhgvlF+/dJAn52P8w+vPOrUkQe1qLJFGghNhP4BDVC5ChqvY
zwVnd2jXMfLfi92qkD59Pb7AFfyv5xMzYk0hr/gqDQ3QgcTsxCgiv0TyB0335gi8+6wES3xCKixj
mHagchPfaFocr+rwFJhwnmGVLsK5/QrSo29MXqBeMeB0WTkTMxZ0fbEclSMSWD0TOUaChNDlCYt4
ecezwqXExcC06Emt27WA3mBnjiOp8mzN6K8U/KBsuDn6jA0J9d55q8RZUR/Ckd9hArJ1DfoJ6K03
4gO5mVzHvOd6icaeDV0Gj32jmQZ6PJElZo3OE4OxV1cDV0BnDsjrY7iBpukXBNw1RDqzKb211Q5I
YlypEUbYl1dqALz1njmjKr7E002Ct6k5GGqr4vtIIzt4xbpE+rd4NNlY74RAAiMf9m3mKkmGijPQ
sZtITdJmBCoOAfToyyc4KJ7nX0IejalU6TnyJ2KzSUq0LXVRWjGv57vT0aLZl6o/B9l71ZBBY7PZ
V9W9PbPKVjZgqTUWEHSrkha5fVMLKt9gLTIw9w1cAQYCqh0kux9xVIUT1IFmpbh6cKC1qHTzULAn
2U/jN5SaAm9bTddbwpwFWFHlQ8ohoL2KfPwe528Q10Dg0JixYiSm+3zOcxaAs+g7mCP8nDUm8cEL
g/P5JUBlgM5jl9Cy/bDPXpnP++xkVTJF6I1VJzft9gcxDpwu2KDXDlad4G/22HWhXFIra01YUrJf
5ZAFRXlH0BTMd052LVH4P3L68gG9Obku1qX/zrbubvBoqUAjgJtN3EnVjHT2/rSVOtGgMJ7uUppH
Kbre0LAwcKJMkDlCOs6wEzukfRPBvIdZtBsLT2CMqU2ioqV3zKxUJEWm45Gv1WCX3KRKKSrralya
s10AZP8wb/0jd53BPLD2wa52IHNMC1W8Ykc/U6Sl/Hytqw7pQT2Z10nLm/FWFqRUy4xbJZdYDM0U
I6PmXIvrEN0jGCiuAvnoywUu9FfDOdPN1fZFYKphIlAO3t9vbcMARZ6tiL8x1jtGta64bOHgp6NW
YaQI6UCRPhKt5RzDc/cUxxyGc8vZMYeZ/OjBgbOO0nDmJH310OOkyJc7ms8ZEedUR6KrPQmcXONJ
kwGrLARQ9XISOtYTVUerCG2IIAgril6BygOTkx2MAVlBBrTnipq9jND21u9calffJjs68iEoNtjE
bawkIZmmGNl7HxxrSk3pi7c4NlH+8bxhvmXN3r93GRsHPyTT8l+JC9GtD6YdgMKdefrZK+f7tXk0
rmVDIL27jn1RdzufOZwXjqfNYCVMu7w0myLQw+f8M2NsSsEsWlw1ok47gnlxhxohGA8iJxWsI8rV
zlI9xJLLpzFwdnfpIQHspN+rU6WEigOYcxn6flhLGKOzh8TITC8Gg8eZTco8LNt/8aCYr9bXoi12
BYrgNS3WrrVZ591rYf9LbCWiAkZwimErmr9itSIWnO8+5WvJgKnSBpftgG6cxVE3eDdiJiUA+9cz
k5MtjBMYXmRAHiJKMBBiew/Pb/Gj96ev/6bx+3HQSWQhW9bUrzCvRZF59xZ8mG4h2tQ6OshVkCwo
G/qAaiNAzfYlWQmSCKfNEnZXa7rClJo9N4lSfi0CJfkaB2JxLR1ZU9/Ya/qOkRluWiSp2CZR52gb
5yEUS6hMaPLZm6VWzBkE0VeJsqNu1pT0ryVRFmnbxPL2Um6ss9DC0hT2v8JMcw1BDLkbRP2+oAjo
GDekG1MSw14YajIt174XIlGivr7bmn2Ly4gjf2NPeiqpAYQ6G++8V0hSTwQJsi1Swsjr21TcfhRJ
tCHZIR6i3lhwEsxOcrFpa3bB4JjV6YceBIITsHUL/P6WmlZU6OWggEfeWDSWtDPFAxwZHNeLzHQr
TFB7MF/XPIgUqVdS57aFa1RxdZ/ZW7tr/KJKHV+BBv0Yys1ryWKOqCI6WpAr8Idd1Nki+pJxOqkm
FjP5HhpFgeUXn8zpa+DTmZjk61b5IctLSKlYN+mxezkHOE3i22qjs7uWlGYXVgQ9mtImf8bW4Sg/
oZ49j4g/AEb8KFAuOyxGxHZw46IXbrx2qwlhL49gZR225rLTJJ6ZQCLzken9EZ1+Bw8NXe3e6g5g
SQBn/4jYdDVsuOGY1Nm/JoXma7C1qsnttQ+p/C6hroDNZ1wJ/j4hcgQGKHc5P+g2UoF7yk/zqal+
J5BUMTmsdM9sFlkpBzFonL6mcOIhvxUee1G9ActU/IfYoLvDFjcEcSWAydnhS16E0nsD5mwlv6cJ
0jadaz/zFGXYSfn+OxC3V2gdMIny5LNSHUW4Ti8SiIVBVPLjNjmRtxBZctvsJ7FzRKJC2zXhQPpn
zXctlGstSxy0DrOMUwRiAIBdewrUjxQAeWfu1UxNJQqZrPVUd6D6SlU/MhRDFmyCJrvs75OKWiGk
z1TWbQNmwAsg93I/3Qc4xlemuu/K6cNhERLcLNYmGEP0nwbHXetC6Mhcn2wkKfKSg63Hxp1Y8sXD
8m4/jf0+FK0iH0w39eJjdN+Joi27F1sU+6Ug45BxH2eLBdU2CPtlHwzNpuSHtyV3bpQSmS9Tmpbg
PPRceZXFOR8zj1b8CTm4aKVMvoUzXgFGhS45OXSMNvlfCVjh80cmu2m9Ph65fmApDRSXM8p0uABz
/fPDLBY7F3J+dOm9C7B+E8rBCr1rRYB1laHKk0ZzvLC/ILUrCPF3XOnSyY5eRnI0/qMGxEHDSU8K
TyARfuOwQKe9ZcKD6IJVgpkEiMeQxCcjFRzcgRU22nXUXwmheBoxsxJnezNqVQoXyqQldtscdY7i
msQkb1KHzrqH8zsoit+u5m/Y6XAGSrcerd7IK6Cx3T17F60OskAVkVf6Ta0cTml96/B5gOSnZxOr
86ZVJ2rhZFZv67uR3l6GOciZXjuQA8pjzMnVdh89wYhuUC3vpjp9XgU+Z1g20g0MyI46ApSfiONX
gJrpdzORGbVgZ+LIN7EzMfRWPi64nvIDDWidznu1sjXFAyCPCsH0Ad42h02sdX2NCO4qZvSLYMap
j58yD+uY3/VVxAesobyq/HTtP7NsxoOpaXXtgVssbRkBha4BKuC3YDxBQej6UkvJ9im+N7qc+nVp
BJve2eOrOZNqNMUhCfR03uJ/Ma3/sSnEV1zw3ymTmcaA2VyCBXQiCJHIMjr1CR5N+5LWXLGB/ldA
/lMIGwCTDyUWM+fC8+9WN3bnANNkdwtPO8rQGh/aMxAbZv8GpQG9wtSpq/LuFhg6BH4u01IMHZvM
g0gN2mCkMItHFQbRTya0aImD+4bVuqxGEN8yQm0L1e8dOdidCL3RZyiwRDIw/nROng0MT+EVzyiz
L7vPSGDojiKr+I6RwRnyhLR44n0/Xb4yFFY8GmMkuOgwROinAD5f6KbZluAtJ5uGltlaGMHDuS5S
cIu3od289bptOo820YdiL8L6oKvIKoF1blJXHkJWoB9PsDHt1jiAgStAQMVJFf1HcU/JcVSVAZ90
ouhHv9hCG+vHrrF3dJfXqHSx+fvWB7TlE6ohgntxw5t6S87xSHM8KUZQl7nIiCuMARIzyKLNIaCY
Eo/4p3dA0XLXVJ1MCyPZGwXDh8G+Bw6ygTmWzhj/VV7issJFMXJRCpW2Zj5lWa3pCNItH6lQOmnU
wPIQfFuuE6gK9PHrESlD56RJrvHX6EUPUtlX3X/8SObxkMuEH3VOpLIeqZw014K4RhTAtodwkVpT
2Q9WnjlQDbl+4QcDlWicisBrRM51CUgz/nsTFKjXXLgohpv6t/LCHUQNkq3ajsYCfJHS1nJ+YU3w
7i/sh37ojb+G2FkhWV+3v0zvRnDN4mABV0gAz6oklpot89aDpVQFJYu7gJh501xuM01VxkTp+F/c
4jUA65exqIO50diFhTVqvPMftPSajpkFZBZM4WgV6EolS0KjiP5r4gYiZkYSlVbu3P4kUl/lUdxx
wIKGgn/fPMXc2znONqG88IWtZE8kmhTvPYvDAffCdo0O0HwQOuVuaUDHvWlbhgOawYXXxmgGzylx
wSHhqwT3HYyFkQpLSH2EibXED3BAOG13jbh8Gp3Cv2lQyu3WGiMr0XEKd5yv7T9ws5fqB6Cg0MSo
tGGTotZs97nNaPUgrjy43bG8qArVj1+4J2eQn2tGAEAcdUET+e5MN2LfTPlZd5FIdeync6zNvPVk
XsKJF2OF3APDdK8KwNyTTF1TaS+DKpxkLcci0iTPOk88/B2JeqqpbM2tAVCj0/3X/q+xpYTfeYRh
SdNWROcIZ76Iy3WxrCUowd08IiKcImmucaieXDIOcCKLZTKLykIZMJ0VO+7bW6TKt+4EUlrD/ydU
CWqatTf6hzbTibuZZmODJT156vXgHmBGfdGEl+u71lxk8/uZ00rNl5ZG9Ra0bndjUo8IZPjoVDbG
j6JrSb0dFoDzZ79lCYF9IInGTfh2HRMjdWoZWaS/5MJm/m5UL8n2wJrzaGdhmLaAbk/5hNV9ZbdM
/IjY8F7RK6ix94j80MWVYAwlpHcGfJdWhuqTGBYn5d+vF1RofO3CAfyXffzYzy/T/nPdp5oKtBW+
8NHwyokpFO2DbhhOGtorPNG5EZKTc6Zq1uR8Nm3E4LtRKlpX3lLNAD16Dvb1fQO7Cz3Hg0X6wxzM
XhK/DriP0hJ8b82+/wQX5rzQ/yUUIifGrqWhw9zHpmVx/+D4Qs7Y68ixV51avjx684imwqbufhPo
P+Fjdm9nBE4fvyveXPMhreu8Qy8ER3RMunezMBf0gdbRb9X90JRcMxlDsKLei9dWPzZBON8IzI/q
hrtUpbb6kENcs8gk3AAfRiUx6u/ylPKepfRYw2k9iWYzaV984ggvl6VZJYjQxmm4lHdHc1R+tBlN
zd5qYnhEqn+PaAWUi+Uyj/3fLRiVTBH5sZlkorRroKH5hgLPC5jt9vLsEwfSJoC6Ossb5ZwXom4t
JZ9mOF46MxsHBMdcJMhvqNAG1y6jXbm3Lin5bmsGTbXeHt/CwVQQKoQmJZm5v1DoRMRzDDgtmD49
riAJ00kbbHtIS+cKZhbhGIzaSZXTN6GCtNsbfVump1aAWmnmhwRm0g42Fn4eansY8n2XEV4G1Uzk
+EIcAhfedjNBYpENOmR/PzONBWmzqtAslm/dwNqno27iHpX6tI+NDnti0vQJNFbvA9gAiVqE3qlf
hcnxBl4PufP5gSCZ1/s6iAH2a/YtW2sS9UipNmApg5neeuHrJfXLK2D9cAmvCrFnoI+HKO2ehPBl
S1cx5jgJHlg2Y1rqjkgT96hfM3EsL7tLBBJJ8fzeriNZVgXKxrg1JT2ijIAxViTzYEWIjbzewEnZ
kXTuR4XpXtA8nxZAbUBFbrIt1ZFmO8RF2LaGfr71ZZFUWjoZ3gVHYUaEJQPFTwLnRzItI1cC1lYu
j5vMnXd7dtKolOtNAA38Y2B8GRa0D5949TBhN4VzoKnD/28g19m5afStTOxTskEm4i+v8PymQhUN
wOYj2yTS4Ke6X9zWEIENH1NYkETC9i8J3e5axy5qmjG2+Z37njt/Vho7vjghHkyAzArE7v50sAJ9
/89APF5P9FcvMo5UkgW4hciBypPJ9JlH5Cywp6KSwyJ+GKcLhCKFMxa60oms81n/FlpO0aox9/h8
u5yUNYxM5vc41lCVcxZS20Jnk3x2Z39UT1XkVoOeubzf1Vp/ean8sfa3hGLRzhz+i6Yo77pnS1TI
xlr4XAjl65xTOP2BDvjvZsqR0MqwVTKw6rdEp6W+g58KMEBfGBE7UEhD05Jml/4NYCYTYiNHajQp
xuuepw35ytLAAcc2Iho806weqiYUIge6H18+KFz8XTXqehs1nGgmvDmO9MmTkYg4ZAAO+ogutmGe
KagLYkrPCrF/eBzwhI4n8YvQgbwlHYdHihLZOZi9MBO+63cSdiwrCtrzpMZnqKHyfu1s7oBpNca1
L/u2RRS7VnJrq1LuIVNEjK4GE03nzyUP+WLuvmaf9nxiYcn2iXXpfcBnfZWw/NVk9IR4A06flOfP
ZTxpMbcZ3w1hWzRQn0Zyj1YuDCtBblxjK8qbGTbuAxHEjT6qdvgvUQVt275IV9gWOd9DgZBuhwmo
rkmaLRShV/0EM9ojvFqfMUMU55QabZE+UXOy7j8KdHZuluEWuD7kQzvRp2ZmckPV0gVmIKgPiQMx
ULhtrGSMylYLXHcFI0zMB21eaH0WPMoqAWugBicYDUpNxkMoQ/sAYwmu7X7DRN9dqBbFDb7Pxy6J
wPEynhKD2mtw1SvKYPGLtdTyAziNH6Lo1tv++9MzQG4w/Qduy19TiGF/HshHMvdw1uIYJeJtup1n
Zd9GNKUrXDpKdFQwRIDIoBrCCGHJegP8YalmBVY0qpooFwWDD7eqUS3bqz2buseKUAqG+19i0AgJ
vQIJ84Q8kKZWlbvUqXdoneL39cNmhCHt4laQ9x5YQjTvYZcWD/gohiR2BeAzILFq+LR9t0UuLXyN
Wmny5ONVlJBUlVq843ViuIigxig+4GnyIQ1EisiZW7Zjl7nSLxU0CKPcl4LQy0rJWKc7nuWCkw5z
HK7dz1wc4rwFRqvcboPYavVPBnUA+vLwwAZ9lsT2crAH8oLspOO+WNFdyHZKROZEq0ynVbRZvtYn
8Xr6Fb/UDfrLlC4u/AQ2PYmraDD8um4UJMe2m4lJ/qiAfskQQHenBJZg47++Y2u7ZpEljHIlN8Pp
UqTNUCYb4m0Vn7ZqAnvgR4C9K3qHC50VtqyavPjpFSgIClCOQFwcQOzpuVxsctwW825mpEVA5lyw
U87qY2kE8qjtw4Oyr6C42hmURy41mkcCJFor8LBvc7PYLyWzxeIyxt/WSDn9mA/iUXtkdpRxpiet
oJvwIZkKjOtKy1sBKGz1uze0i2Kkp39OChg17fmrrkBVCmFGZQLlH3CEzFBFxkmzQlmxJ8AhpDB1
aMKkIcrMYHDsLSIre48QIDWyarEeclVFEari0kxdb4gD8K1uM7iMNbKXCcCOvP1vViPR6FYHowK1
8LlLOJeqvxp9peU3hPcuM2iumwKZ+7b2Aa3UbKvxe08Gm8d2+TC0iRR24GT50BxdNCE1h+NxwVnB
V5W9a4vfZNBauCLSxVK+M7S3BzkfbSQJuRVagbMBpO+XryYN8Mm7azk4w99grUwIUFobAEQYu131
bzn6kGLduq5oUD5lThlLdJdPkc9PHInSOdO41/h33B1kqkr2BBl+3C+72cVMPKNNJIwODVMrQEgz
3uV4ujwqMKhGQ9CNXeCAubcVmL4jAPfSd2tr35J6q4fR53gqNOuq/IFeJZMXlCilV2s9FoL66SWf
RXvGD2oflL4anKRuQE1BeAga5ahplDG5I29//meGEyiGLV8GZybgjDVpOJJ6BsQ+T3/zlgJaEMeM
dXbMZnZQNjTeu4ia/y6o7+UBwvMAb9V0FWnroahZPsIaa6jVJh61FMwf4QuoU2UjRADLqnwC1xNI
LiQLoeGyJuX+4BiBDNhkv1GDl7a4lP/h4PjbFZg7ZQMI5lYl8imUZXMmlAdP1+KOAAjvbs7DjAWF
tN9PMuJbTLhZSYYOGH25SWvBCDEVBTp8xx5VJPlbfYLQvnC36B1tTS8IU8cS4vmaOJa2uzpOv+ma
ULpATwYOWnq6cH/X9S5ypPX9r0q4ZHhewdjRINtR/W1vAUpvFpmZ9fFsbKKDEsuxrRFu9Dwo9vPm
zY14+AjdMAVGv2Fky8qvhsZyStsvFf1Da2HclkMyRlecL/aehZX35YPiCn4Cv4jXhmch1BvTMVMc
iswZkNi6zi6U+dJFfLh27JXT+EBBbJVtbZ2C+BwlcfUnDLlvpU0pZOfSwIOQGlOvADnI+t/dhcOu
0I/sBGOJ33tPMmKQbxLt3gDVJ26d1TfHumTu54fIzUVZKxLA7CZ4JoOZgqKWlh80TWnxS9v0o2Fx
X966NKHwsNG01uaoR8kfwIwEAQGSzGhBvcrqwQGwfPz5hAzr8ypjujQFThRtA5LcYQk9Ymj9DPrU
yzvZGivt9M8gc0D9JY3Fyg3XetTK902PaYzaGrDIyaDIUyaLYDF2mGZrHqJesU+C5EaVWvXn5okK
Uf4Y80QQ8W5knSVCmCuKLzAxuKT3pQbKn2/hv3i80szZqt4Wrnzv06sEuSsblrl9lFWFxZ78Zliz
FWIHpiQzvU/wYBI/rKLuS6R3s0IE4FrGYQJ9N8rbfhlKXO3W51Qp8ARqyqZfxeYVAlxQMi6RHFNQ
BXYka7T2jNWWAv6W9EUf6w2XdX4hBZCp0E5sfmr5s/9cKxuRGP9OVD/eDtX4PmF+Vh0+gpsiOcYg
sN+RuPgcF9drUMduHdVbgVL2DdAdIk9vW/j6sgEAwq/238srjezC6owIrEFRSeGfd0yVa39JEukh
iS7dOqOGoJRFZ6A2Ac1/8Mbf7EbojUDlG1GOryemGuAsJojlLPLYKRuH7qIUW0pTcX/nEpIxLBGL
0d0+OjVgg2nA7OWOt2C1HFH++oP9/VZnIUSLuNQ30+5rsD3n7dnWZTiffP53ZuMF9Ko5isYujvAj
Lyk/awVvvj58FqUMifZmRkWSV5mZq4nEAzG1IgxnY1msN1EOUSlVgwWP5VH8W6i0EbPwcQBQxuDF
gfDo6uF4FMaUhP3mKobCxrfKaKrk8J1s7AGpp3wDXmREJmVeSq96WlWx8TvEUE1tuinBSgBmxjDt
FtujoUa+dmFTAwdNO1rWHQUbfn20/CbWFfAh7E0W1H4m+STJfD25Cm2vSoiTGtyN5D8QtHTysTLO
YJU5Q/HYoIxIOSelFeyoI9MrTVYmf/bLAkVAG4qGaLpcx5+0p75uW92e174ybNiHUEds/hCD5KtG
bdIWk57DdQtRQnkCkTA3e0P0LVLB0qEzjYauv6vdlEYksB+3zUWU0xa2ZxZQbVgVk/uupSg5owf8
7vGBhwuzfa0jsb/D0sH2aCbKronLjqp9MNvkDWWBrM8+IPUVIeDBPr697Me37rqp5xVCQjSpp18w
kwyp9eKYExuCpAHbR89okvYAQ25r8U5asdy/V+ok14j26kdwVG4l0fWHCeAxT1WR0QujgGWjUGpi
runHk8NK3wsgre7UrPoRMxTLyI4jWIYazLh+qGzRY3pHM1FmcefZafD70N3TsED+KIxpAGr8MD3d
/BUf1loECXydfURsjKyQfcS2wgUOVzN+rq246u+T2rz/UKD5cWXppOuxDTNNBdAwDHq6CZDBGfFL
T88oFq4GQqqm7oSNbHyVHHuPgzxocBhLGitHoWw6MRopeaamPxk/j4CxtkrHa/4zplPHLnWlcFD2
SEa1Ks/eouN0h4K5CLQIHzsFPS/HdRtZquimf64TEDPbaEVC41Bk9lKphYYRq+UOxO86Q5QnX4lV
xqMnnm8pWDN2nFTFZuvXevF2Ykc029jj3ZQ+JXGQMezmgl6GO6Tizb1D5oupAVGXxeAmIOwBlBvb
Kjlh2L5AMEOxqRcWrckZsPndGT/Cn6aL+/iA1XxfXPfX8qgl+ty9Z9E6kVFw2rIEHG0L6/UzN/IQ
VzRtEybQ4f9uVBIt0e9M1QeLZ4ryDp0iPUdKb0iU7OrMzhy6jnjouIFxGQPaP8Wx54Zzh+qLFhQs
SLy0vjHX1X5gdXPgBDV47GinAimpi/Ikz4QtfOngZ42v3azhtOfKbxN0p73Z6ukA4O+BWEGBbNOW
xyInGalyRXDh67ITq1KhRxsuS6hMqd3/blAkpuweWnNsmkk0EcdhYoIZNB6ZVHEb4Pc91thBiKUz
sADjz7LaaUuyE7r+TA/teeHChd6PciehZEFrt2feqUzx/XQiRmwbcqzspKes8u+xCqRosorvHh3k
hZ3MUcshqDDLy1vkGshoVccBb+YEA9eCeDasrwEEMNpm5WHnFJgl41FGadPdWj1D+Ljp1aJogHEe
IVDwKxAdZ3lSjvB0kgoCcTHqzNO8bNSCcF89ljqLPP9S0f2t8CPv9RpqazmSppgx+6/N0hS9sMKM
XEyXV10ulNizzCcjEkZ72C2psWVwObylipqisJiSL+e0G9GDHlEOLw2xd69SIotJA45loAr/n1cH
dw1HxqTJ2xoxl39HZ0B9+reK9PL6O6gmp4qIcHeidfekYxLLkc6uO6Vc+esdSYNDy7+Imor+xWW9
Qo03V4Xpy/vmqWvD1KLPHia27mLvvLRgkP+EKWodadMO0YRE482xln1xLzZK5cUkDFDhaGthfl/8
zPJzhRDcX3O3frYluxN7oxkb83891sSuv89kS+owARexFZKIshMwiTZUh3iQiWyhr8JFkNuxeKX9
wBA4nulXJd2e0gz3MF+Ho+c4HID3wNXFtStjq4cBkbkjXGCSPVNYQPkMtSoY14iXuY3wHAoZ12LR
Vcq8TakjoEvZPGE1hVzHS+N8K+abpjUB1k4rxVgnFuxgp9uDHDTzGqCc42t820D4w7NeXMV8qjFz
Vs59zq8RzpfwgVvE8WMedpsEVIHAsFbA2n/ni3E7v4IbUrtNhS388XS517sPn+NJKdBvhEorzuUe
Nn0MchgTwITTRtbQusgm26xfpN2w//dYDVl/YAxHa4h2+F895Ge9RNcxBNmJOIXoatmbZ4uyvKZf
ryz9nBqZ04nrHvFGuce+XZiqwS39MeNmbArxS97XR4KQUmzBjx8po/WTjEPTnOfmG0Z8cz/f+qpg
dS3+pb4/Xtwkp5xSoyrmKWhcCTNV4E7C/qRnvG/+KVaxEDWdKccD5tk0AtqMP4CBhst9P2l6kIV+
gD03t1uub2tGZwcEnNd9KRfqZM8QPTRDMIArNON68QPg1t09hIhRpkZM/NdHKMkNZO27bY/8pz2Z
ebiVR/ndBz+KRC5eYzPJEcAC8WXMvEFh24EBqcuCxATAkLLG2MsG86QJnvn20E6ze4paBTiJznut
exBCdvHkKL1ZDXeBpL5ordOalY77L2zawv5C+iAxo3VNVd3s3cKzgS5G8V1l1ix4Da/PljttcIQO
vOarcHRa0GtdHM9vUdHsubvcDXKUhkpxI84kPSFIlmZ91+CVfUHSinmz92+YVcfpMPOfHv6Szm75
c6S+yKzQaHKeSBWg/DO1ut0UcAKwr3cereUF2jNJsKFPFi212VqRUKyAzh5Dvk+H1MnNIjxXLNgc
GgFtVkXnfzwO+i41sj+Ay+44oOzliyXm/iWJvbIXL5yD2cgOrqEH/+7HDh7kHEkhZIsyJRdexrox
afWYVFOLYLkvAPdb5NJgxLHdU2vHCLjI+Rn8sRUCm2fAWDHJnZpD8upyYkiOTSQR5d8iFm0Da9n9
IuYjqJFRg0dbbBb3ZJ6oz3WJPqm6tqfzxruhDAJOOZu9jKxgJjb+jcUO1xdBSimUEcYtSHUQ2nch
3S81EE0JJLMRA9s5uWnGfdPrvfvQhSn3qpYoE601/2D9dBBbrOlZSjo9ye9YiGFYHhnJwqQFD97y
P2nw5hANPZ8KsaByZiYO/cydNchdSd6CXf0gVF0rfX32Tus3ysv5WB85AvB1D1XRGrFv59TxD3Z5
pnSbjocaMtMHOwA6OKmwQd0YvkodB6VdFIufTh8bjVzanzSbPvgrfpCunjr5TSBsaaQi9O9qYmiL
X/8zOO4x0GOAkaLob0q3hyzPZrCVgoQV2OZ4Fc87UnaGVfQuYwTMeJpbfRqF+t0LFCFtoLC1Ozwx
nhyicsi7XSDou1U/KLzWJIihI0qRfp1mfUDpJIvS17NXs70GOOm/qVkqZZKvPx0jOHuaRQiOWQr+
ntMD5E9X5+X1NHk9FrmlBvPfTg6cQjEjVVPx04546XqGC6zq2h8+7kC/nJCpYVMReQcNz8LPBnij
0UomfIKlt39hIahW0iNcx9fxOeJ46bv8LYITJOk0BPJYieRDY3i5e5d8GHQouGCP3Vq/4TfqEwE7
TROu9F0UBz+DJ8p1eQzIK1+GnRQUM1El6kCQFWT68vlro9M2YR63njGWxSSqHXmqVKOyEgE088SN
qvYNyQnxtG1ZML/N0GW8hlDZrxFLkXpBuef3ooOPpLcqDMnOt1KnQkNokLUKxECLoRVXSRIBbBvE
ug92RRirxu2b+DniO6g6qtmes29mwBx9qM92oKmw5CYQ8sor1hjkxQvHTOit7DEZuTt2C2sqCPzZ
kAvBH156c2ZboV6x5Ve0DuV+/VZbnb0qDtHbi8vB7Nsy9HYC0Ac8f7VPzOZ33xAGF7yhwGDWuplO
R4QJlV0GEwUmTq1soi4jg/6vrWuUOB61VVJaq0y/hg24z9d9XrobNs0oQ5nFlv8Y8G0IGTXp7hvy
FNIqY2BuGGGuXlrd3CyYoIT0+hjB0xZDKyomKmjYLyAXIUia5dVDKNzxrS2BoCpByoMTnvrXf+7P
NH04cKEnXNqAGIbqzVymymJmYuwxi7iU1GOBkRVXRe+Ma227fbnik07W41rHh1yn3wvDql71vR+V
LWfborUX2Et3g1GtNud39Tjn7PNXsNEVK52fPLnjIv3548ZvTGeHkbv5L41yuUJF1DPvzFSsIUtj
cZfERQq5J/xcQlwS9SJ0+D3NlC6rm1EBY00oI69Vpfn7UdaKuU/shkeOIVzXLMuKGb50JN54bpXe
IvQXW6PSZSvbr2cUFU0pO9yBly9lWxPJ31QN7TXrGFj6iJi26ylYL46FRMpdI8sdIsxviYPQZu8c
6eD6/k1+XfSAHpULrbB3NXO+oIvG/NwBw3D5Q20Dsl/9wvuHaQidJxIDCBPmhI6YT06shDUOeTKA
AWqtOS9HobdiQ9YYXrKLKX+qCU89ch2+sBmcyG+XQn7vokSFgFXP2XUDhcVG46Dz8gglO+tkPsKa
qy59VjA5ZaAN2IWns0BQeqBJsfDUUvJ1x9CsOy53AuKIm1JZAD2w7Mz+NKCs9oLRex6iigrq4DWS
ZSzHRQMlEhGRkf9BEVEJ7wy/ZzYAvg3kyFaAAAke0EPo4kcD+OgwJB84avRQliHoDz37CKNgqoKS
2Kz43IqFjDLwDjsx62Aq55Bgpm3YkOiyCi4RH3vbFNuHGtZ7243OTMrVx4bbUPKl29UP/2iW3j6t
mF+TYPAsA3zMIX4MBa40qapEwWQ0139KTAmNEukcD63NiiRGWtBtYtyxSqHQpI5f9Dm9Q3ZEdf/g
hl0r+NzLRW0aqthQM4tLz24/OsP4IBnnBHOKzanI6+NR71zVlFgTZWP18BN5KnJ0wZHD6Wh8wduW
y6F7H9FkQAcHFIkv2M+EqsDK1i4jWZIyypV0yW4CUJ1w4pxuH9zjQzARV8N6cZqA/YlvW4OSZ128
L2OTh5ueRQIkYxMl9ONNLe4A+vHbbEeY2QDiOe93ojmXPe9CEjpyJHuUJ2VZG9zjsyXXCj9oFpmK
EmkByI8zSTIp/iByaVYnBYPVPNiSb9wJ0nGZpPX11UQ3OgfgCQtQg0JJ44p8m8cGjDnwS83/7Hfo
aQbN04KwF7+MwALN8I6CtPlYBBc9uLOGSEiiyr7z7/KFQUIol91+0co4C9iGByyRO7ji/4Pb2VTw
6ct/Pwz7WuAVJGEbnDkPuYfRQVH5t4UhYJhJ6614KIdgDEzN+RRpvioa+PIMvCGIDXi135rTHaa6
9iYixwTdnxqMnQqmVwkucaNf6EZyvT5T3erbTxVRQAyCOzLtbsfP9K7AkGOlw65UGkQ7b98p07Au
BVKhk5iBYLYNC4kTdN1oNIPyg28hB3gsQleDEn02VedDZnZHHI8bV+pSkW635/J2vjOi1S5yGtCT
K8tWevbnroMhWkuGNhLQaBfNCuN2iNPxXu6FoAN2qCCNZzarzsoAr0HR3Tif4GkJWS2DY3zieAJT
g1j1AkmOp9qm1xJNQpSjHOhy0mlKeOnZrcwRHlF+0VidFczBlL5nP55ms1KPKKEbQf3yXdw/qxuM
8fn8R1/0go1fixUvWs6HeqFflVoPyJHcIQ/E8uB/3MCatf5zhH4NZZ0ToCr2SVp0ikH1YFge/Tol
+bIYp3FskA==
`protect end_protected

