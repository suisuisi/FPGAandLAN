`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lOovj60F/36/SmS6HGL2YoZqU+R6HMaRWxyFEmNfnbUwXUI63tMlaQSgHxSzSPBQJDg9qS6YEHxY
xHTVdrG0Dw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VRGCd3WQIM/QlAXLFeqeLkJonwLPKfgzsiA+iTNkSyhmnaoeFXllv2y5XznGwnukYc6aq2TmSHpo
sCmaBLCnTkuk6FBvkcKngPCPDvI65AbR8Sp+iSUsBodg7Za/P8WblbA4Sp17AkkdU0US2JwaxCkO
l6aCv6PUhnFHVdonSPE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a5W17eDlPJRf3DEqIhWY4sCFWmuQ8vFQ2TYiMnZdvyW5ti8fsz0fz4Cx+wFf0qqBfp3t4NJLXnTN
/mVV9NqBoCK3X1uMAZTSzpZKJEEURoBzMNOauReFuZlFN8pK3pqCx9noU6ugNyjAqB+Sjo2KQRQV
F8mlKKHAO64izY58gl2ZoeqENV0h9Ak+la5W+rM7V3HWbZjnS40i8OiuPRsFZsLKAw5f7sxbNEKE
mkC+mr16HgsBjCGS3hGodhUlNLAMFC6bbo3rPWk+Sp62LE6Fnkij7hoBJ3cYoebFFuVrmdvRaad0
AWxJusk1cH/brTz+rW/Wx0NAvdrgmGLOswiQzg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/Kf5sf9tZ4xHVzMm9AtacMEqNH/0YNjKEh0GQUyxICblVa3UkBoDtSK8EV9pzxphPSten2yV+Lb
gsOS6km2fKlQ/s/sG2tAjnhJXvU9CNBe7jRykZzpFmqdInRzkEgLQV8wbdL9sKvYEo6Mz/58q4iq
7Fha7KJV0GS0gj/Aekk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qld2FMhlHX+jtBJiVJ8G1TlzDdkfnrRXO/gx0+KIAl2YaV7t/8CzEqAC8ah+OGu+hgXORGYExRAs
NMcIfeX86MCrW/EW883fIdupJAsW1iyUlXBtezbeE9+UzTmM/r/7rAOUIVau08GDoeumvt7Y9X3X
uR6CTceHr5/G83hLgUXKCT0Oi6lSp8027/k2WO628f8Veu3twv6MksloNo2XaIIGKdxYOCr8gCd8
AH84A2lWPMMiUrAse31apCd6vPk72GYY0JjsD+gDCtaHOP68iHCZJ5EwtcfnphfQ45rgK2X3yPlr
iuAlGtmeyBhX7LO5t+pGk+1x6WYxkwcxANCOYA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dXCMxoBFa4HuiNpnO4iJDiL8354Nga0YEylkDCw9SfhrYiiaWYdYIPDUboAq0inT/vEM+bt3/tBt
ept8+U+DPFCJAkX05h2u++Dtao/lE9PB2S/9phDTIqrqc1wFkmRiVir+h1trMVLi4GgU3svUAzo/
O7O7PiW+VNB1oGyQLyDtdnpkAWKs22i0E2HWTjU2jioNImqXCjv9iudNOrSDIE3k0EsgWDO9+Nkv
fq7GAK08JIu3nx17lWLAtHg3JrAtYyyLbcUTeAEcSikaBcQXc6ExpSpaH5f8gshMtb6H+4/LEYwO
GDQNl6AaOOKGwORorQZ8BVGNqtle0GIYQkeXHw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 119648)
`protect data_block
SRnPres9zl3dEAaeg53tBFzT4ZF3qdHLCFPfIsrqvSBNbOrPZ8CyTJjqJE+1Oxu7lw+P22xtetL+
FBmgFG2VM+fSODc4IetzFzq8GpfPaYyP5yI8V0COsPUJVG9PuVf+O8mBz/Uee0dvn7J7UMUgET7s
SpIt7eMZwh7nuudFLHwU8MuS3V0XioPsn30YqZzL9DO2Gp0v7DRg+rM1CJXE9TdCJOpoUEUIr13i
XM9UrbntIxjXQIIlx1KBSNAXRaHpU111LE8P3SJmbyjPEpC3yAbfeevaeSHnS8sRq2TBFzmxPbcr
bcp12YGDKj3Ad8shC4vOieNbm0j/dIdjEPO3lQ1m6UTxTfYMF3Z1PHQ68C5u+GsWN/i4ETdOa1lj
M1QLpjDsKubHlyWs7gs7GLIXJSxLEG9hBH5kKWOfD0b10CGvDMGtdDqlqkMADyeyiCOCDL912faj
NNDj1z6uZfQYo5kbeoRq128netYqeVKi42pzQwPV9V48Y1tqwOopR2RVRWjjdzk4WoEGABPHsCwa
t6Gs9zhhpeX2YdvGC9h0GGU/LOTkKn7EidhhbZVuZP4byJBtK71c+WiuopcuKx5Jxk4qIPri9/iN
YIx1m46SCW+jEtJJibsYSXoRheu2KMAbyxMvMba/yhJoCGhm+MB/vLOexOeUfj8g5sZob59lA75X
tmY1rFzGo2kTlSqv2WHBz/Ue9CkKwnV0Dd1H8qBLEzZ1TzVifw5isJ5Hbj/yeC/pk84ELgNzSiV0
GE6RK1y2AZdK++WNg7PmLCq19DSoWw7I8g7PmWrBzqdhgJExPDZOot9cOyyn3zlk1qFqEIL47x/V
++s1a2ZDkndRCupu818eTBXxbWxkr+rcqZ7RIn2z/jOt1SH+jNWa8d4hH58VWyTHWFoxmyDnMLC6
2tNLV4ZgSszuCe8nPH6yXCGB87mbkOWVcgONXTBVaSS5GHUY+fZod7SLjRimmTz1+7J5bqth04xT
VMdqb0HvtBvxzGiF+lD2F98p6eCWoXwmT6IUiEl4tHzzLPTMkj5i/N6YrVZsOIOb19CbQM+M1dRt
PmyKKWGxXXRWYIkzUHSS3D1FvqkWiwdnfRiRPsFhFaSDlWpANYebuv6tHwhwMvC1OWUJfQmnQk1m
RoU+2YQk2Igh0E8lqIyq/pqYhA6K1QgJzl6UVDFILkwjI8pZw9Y23bf9SzFpT5dbbrP1Vjhi+4Ju
BT1Wa1DLYjkx91MVkJknP+1vM3YYE2/NMwa1CLnOqCSmURd93ADowYAQ4zspZuc0+X7X81thB+uH
ue5LS4HJxOJVYueqXk/qgLhznicNiWue8tvHrzukU0RFuEnpK+99D7eXwdLyPUVFI1wCMP2hTsnW
6EAqQve4JqsdJgsCYbPkt7Iur28amRZn0hwrizOdfZgppxvimFhnvBxIUS6JThwJslnqRDF5XGG9
sfiRIabkMNXiiJ2h5Vo4Uhz9d2kfCKzrgDzwoJtYZqVZ80Meyz212kNwt8TfDYDzNS9il1YHVEg1
ixcaBcEd4L60TIi923/dPGqPnE/1RZ/1YYSTCb+EIt5R0w7ZtJdE6mipREScaBzxsiUjZ7j4H5VU
ZT1dkZyM5H9TSRy5HhBzxS2CYZDlYPwc8gkA/uoNUlB0fvpzbqI8TStuDpVQD8xU7EYuhAGUV6p8
j4jo3o3X5pxFoGVOfVpDOH2mDHVVyUTIxJMjcZfQvBfc8ylCZYlQUf2JpDF9rpktRjeaCwwziCwg
F2tyTBCDTKdKD+9Xu4Wd1Fg5r/2KVkq5ejrNgPU0AZ0bxgCURok5qaYx+t0e0dn9F9Ftlf0gI7Kl
Ytn6gEM7SQOfAAApD4NagWNFj6jCDoJRUJKpujDCVxLEqQ/ZNnzYyNG7UzKQuQbIn/9BNNjCoos1
lpcz2gqNYAqd0mxbyzTeFmSu1Ud1gY6vouejCYOwC2dpeUm7JKMU4gYElGj7AfPUCUaselxTjkKQ
uC1U0qcAfikiwlkR3loSpmO0GqnmSeM9A0CvlIE0eenxNNbAc04OJ+T9PyAsONmiECIObOd2RJuH
fxDGfIvHiIoBPQKdzXfStE1YdPY4y6Kr67WASQ2r0voDLZgH2kpcP+tuCkGQFlqz6tYXqjgxkOEv
R1tnwUMQ0meFXo0WD/tDEyels4BRtoNsqMIMJJsTiqz4hGwhtl7qBv8UPTRz6MTr6Dm1ZmzSzcXe
xswyA1/qXnKoO0TZaIf+fv37czPGAtEYVj+DmGX0Nz7Ab4XVYAgwwMOY7XeYF7HaopJk+1fWEhSq
iyfcKLliSgbGyXoojqTHIn27vK4qDzS17sTqda8u0w6ahBglvANB+Ep5yx+mjI4t7RA5se/blqqX
Lb/F4grKfvbe4e0R0uBHSLXNO1S4rn5wvV+1Cq0cEswjqXuwWzkqcv+TAB7YQp4M+O3bvgIVpBha
y8IYkfjkZ7bWdZ/VYctOHv8TbQNU9xaREJuqtF39zZeh0ylBaynuC4kkWldLSYrdzqt36dzaajMN
X0G8KuvjT0KmX8anAKa7p1gNaWuhqSY9L1jGXefMHIXJ3PdU5bS7Lp7w98N/4ADh9UaYGCSPLJxW
LEJ3zrHVtWilwEf4ivO5r7gQH0yJlYCK416drAk3O0zOOlUmpckTDqJsre1wkAQlhADiTv4HdpmY
U5Zcsi8w5a+TlIFnJv/ApqqO6l2SXxtSynAf3Yti1HNRFoQkEzRIntudj20iZJ/fv39LgmWl+iur
P71xr53TqT9QR0v2/5Xt7tLhWv2OlAOc/PZxXY25q66uAxKTLe9njD3+6vrUDE9Rpqj8rDobQI0H
iwFyvp8ii/hfF/qRIOeSLp6fILbYDsVJe75vkyGics69GkOBfv1JA+Zrwr8rz7KwHG2dgdkA0wPT
Sf7lGjdTaaYtu0zjgYnSypj68R83DKUPpUsYNWE0eUf3J/PLqrIH6U+oziUyVmdZxNh2plv6DNB9
/XeW9iGqq6pkWGDaDK6fERaIG8yzIoO0lCFciZfkDy61T/lq0KL8xwsGqXtaP/UpCCMAV4MX9UIX
uAdsd2PJRShV+F4Fw6K6H977fMtyDBtwttzVKml1Sco4itzBjKWJZKSpd+0NbHPUKTufVxA5r2d+
4+a3OqFZ3xuF681lC48Xf9JajWxPkc98t0An2hoRDgvYEpWvtKw3unOfRjs9d4PKUqmeZYiOXgWC
EIuIF/YmDY5FjcyU+04RN58gyRJO+EjKfsXh0MKJhIr6GpjY70BpZ/B7BWAHTCgJGod0Gk/nlcap
UiwnBIjYZcpelWn9RUwKfGtD1BA6QGmCohwVg8myGoKUOSrTxnU+fTNOJmEvdoE7YzvGkSqH4kDf
/IZ0sVj5dUMjZ5ZQ46NzrOwET0b0PpO+5W4Y1E9Uj9CeHmqNkxrQhrP5F1D9xh7QMnnh8Sk5aDG3
tKW3ydyNzHYTo2ghGDldE9cBFw8artwi7fkgGaYlNNhc4WbdZxnbyXfYmsXt7Z9N/ymVryU0H1tS
ClL3J43xUQoewMuRfM738W/6m5Z2zmSDP2QOwVsVoU3sbqM4H3kZTpcMSeuEXvVgolHeG7bxa8uN
hMBe2QFCj54BaQO9NIcLsSDUy012pnfOwC4jMBQV+MYAEYyC/wEZzJq4j6UVshrxlbg93neQTY5T
c/401NFNCQEOhamXa+yp9MvKAsKuszeTM9Us+D2xY8jAnLDFh9iM8jye5Gyn5Ygxe2THFcMLabsj
p6yD6/NGClsReIV0giFuWhUUTxskUT586SlrKtsV5hkDRGejHf5Rl0Nl9qzM1Q4wDMmc8y1/Q1xY
RMzqXMpp20X7i5Vdwa+zIhgDTeH+Gx6Dn0LrGOo0Cwi/+66D9Dz8JSfPXKdRuB0pndBVBVJKyStM
YF67m0q+Jn69dutu10TREi06x6H1ty2PD7c0lX+5dyNf4+6KT5mEzbrZyKH7San/IdM73PXcd439
jJYwESbaxlkSaok+iilcA+MmL+Sbx/sgYPysUQcKkjU+NAy5AFjhaw/ScEUOkWRgVYhXs90dy0ex
5Ix99ld48L46rec1dx/HabcGy8NBnrI35tEFDTcOxHtK8hBVPQSQZDWzGnc3pBHNsjzzaIs73xmM
p4SwUFLD/zVK1E/ASTtHV4UxT/2HP3ad6tF4szMEteG+dVDOn3adn/2anbp4YpHmKE3D+bT744tf
T7PjjDtmAXDCtIXLkK6SrR4cYekUAx10Kgb00STbZKk+K30L0E2jDnLe85S9LWY0VlEcAXXP8g4f
kDFuZDkZGculkysCBP+UpssFiORWkvjCNwb4k0U/5ahyDB7l275Ek1HKCrixeH0vVYgHETlMVayx
toLUoRG0flJHsdjBMWF6d5BaFIUBt5wqmM2RlTjs5OenxJaToSVWCBqi8SX6alpnBZHLW7nIm7GK
+8hwsUCU4fTQExCwZlPxFDRFlt1xJVkChL7cr4dbCZ+wQ3ED42/ZT/Qw0P1XrRvkr9J9uzZfFKiO
hQWJzPVGWfFTPHgsOcY19yhf3h2hPrwXXEVkHAlKIotCitv/rPGjjy3fJP80QGx4r3vhe0lDLB+1
4TbwJx0+MlETGydWNYyAbqpEJI3xm4+t25NkFYJm6vp1fl+7RzrZkxS9/IJ4o0oU6VrQ9Ki+VOk/
21QHVGKfB82/w+8dyT9bGQIxlA2XbfAFQuJYhtG6VV+BBIad+N5VI1VSgAxfgyyyGZCqyZvpjiT6
cfW3oHcRVT6PQSb53ov+jRuf8opnOkwqOZy8XTy/N+zWkRcbKju1tA1+38aRglnnm+nJr8OuDUTO
9IbxWkY22wDHcsYe/MG+FYQWCoxzquhw3mznyL2jElKd0rasXGYUIwD6jnRuCO1yjOQ31c4QW8kL
Vhx8EEr4xSSwwqcIFn3N6JG66lvvx4j7MQcwJP9oPP1yQe35piTyHKXMsGO9dAGAfAqXp26ka53W
upsxbouy52c5gRrQur9+68AsSP4+vaYefD8a79TiKX9b06gy35/eps+XOo0NrbMGseUVH4iPKjD7
FJrcL/k6wf2F984xYUqAHbTmAwhAM2Qd9j11zDxfLR4OEao2slQastYL88pkTAU8sxSBERj0jegS
3mO/3e7qTrWeEJ7fXaXDsb+fjuLIor0HUvYG9m2BMLJzjX0VyBLef0OmD0GFcYFgfRxCEdDkbO7G
ZHLOWq/ok0onm2oj51NPQwW42q4UHWFZC4lV4HA0xnLkzmVbdgxQdNT8IrVCm8ABO5Qa7fMePr2h
UuMNennNPkzJtkzPUX9xNYZCoUHGOVPeTqJm6py45c75xvk13Py5rs7TQWo8O+8rpbvg3yc0ynbQ
xvWT+crIVBmJ9aeq0BfQsdW/7uljneeLCBG6a151EdH4R1Upis6zcmfYFGuf4vQ3tNoiLCsnJjrm
tP9/BNBHM/G5rlx0V4jfN/6+lTFy7Muy5pNdOdQGfUI5UogXFOXxLnBsy6dIBD2pH5LHNt1dr7uH
1ls4r1SORmsFE2GHZ/AQ8JPpIm6rHwbkuI5FGZ+c1TRnrjk+O6Y+PSQa0P4qZs5VO98afgQ/9dNm
wfk4swBXNbIhkOlmL6Zk/fx3erPl2gpxjvpK8pyCJrFFFSKGMr8fe7Ab/LZkYDvWYP/1CaEQDXOU
6OQJHwRn3rzaSEg+oG4uQUm25xwwtORk4JCJzy06B43VeQjrcCaBIB+8o5KbV9cOeh+9129YlHmN
FHYdcCjz3VOADkvk/KkFQoAcHoa9GY4uV78JfQ73w/V9avHFOp8+TusV8gSMiefNdfyoFp+HHxk1
58PrLjP19jt+WaBPtdNA8y6eE2zOjrtOu28S5NZntuc52cPij7m5/hpxrz5BKLt43sRDItYTSbM5
arBQ1E9q6p/BsCIf2ZREnHNLEq0gjy/Gz1mqOazB6gGG4KtIffhCcSjXfHo7cNOZ9Qxei8Aqqk+s
M0iaoFIKg01SsfJJA952xlVkB9Gw9DfioRoU5c0cTs7zbFOJK+Qe+bLW7/r/k7FKjAte8BEXxDm5
k887isFPB7fOQrbmg8DXaGxVrmJqWy4fGNZEhaf2/fkYQIa5NLFIR6A/B1APYpx+Edo2ubx8Sx8J
LHUvQIFvgG0HdNHqMuGeSopGVeE8DWECHqWKELy95Zytpx550YfPauMJxLxAYUsAgGTehqiFKe7u
EdSBWeIXMNJGPMAKCrltDxhDGudUjD2qqUhh8utFyag6hWmQXXVX5rGR5hIwNOT4o7+S5H6dYwqm
yklu8Ywm7ekqF/uTkTrzjvrJCVuK8i88N1HkYyhrtDEF6Bi/rZ2HcdNl5zsfk2TWhP4GqWrdEBBX
2c9EZQ9ekCvmCmbzlbzrapkqXHjHW8AiesvZrTeyzSf9qjeGESVhZGHv8z+mTjamGW+0kQBwWeDS
aqf1paUiJZe/xPuVGJ1NL2tY5niAXiPopeG07LSBqzqePLnBF3GkyRCIzR7DBNeCvPnPcA+0Fxr/
jCkP3/y9CeEefqfqm5OmnWdYO/WyeDpV/fFLkG29ByaSGJdf53ULjdegq1QSUHG1Be77EH9Y+cAY
lK0VDHAtuh/ty6u+4DWo0cI6qiMg6+RDU99lpY+BZTDwyQeuks630hQFiZPefx/OoB3pFQ428GuP
DhvNuyC2yIgJdgZWZXQibKSJQB2UadZvKUdl5WAYkPjaWApzMy7fSPMykKnywjumFl0+34066GRI
tZf+pjiPtOsJJAB29K+k4xvlSsHD5ag9i9pZ5HMAFNdOV+KE4MoW+RXUUzE8oAwr1pkyjM4dt/AV
teZHmgfiQ5Tr4KSWi83JRu5WV7FVrSUOLaK8urL0NbPN7G54erf1pCkg6jKGa0pV9bLV93Q5Uupj
K88dHhLGwSkyINiadVEVfJO3LPevy/AEJnwIY1mt9B7QDX37Dq3bInTFi0nAbPVGdY25mi5PDgKd
wyOBaXCKHW/xJmUl3iE9dkhqHEHVPDH7kCR7Oxz89o65IoMbofdhrwaMClprktxGj8Gpab+KjfvR
w6bLlABp+Jcv1bZKyb/wJN/SxzAAAbMmCg/5hOOtKotpi0YrkMBjFasGxeIG1V2VrWVdngm/Z9p1
fqf5U8rTNipfoV4gCuSPQlYlfVPOdSKSHEjNAKhVau8bLOoBXN5SwTEve9v2Q/esdGaDpH6qGYlh
g1sYlyy5TWs9ha5TNEcUyb4JCU+PfC6R+2VSgceMcl85nhpFFnY7BMffFW7qh1g9/M8QuYPOZt5T
/rvo9hQsPRHPTvxznuFpp3FGXVguekaEWnebZEvdjHVV5cbYW7fsKMbQYwOFIOB3zkFxZZH/KMpk
ejPh+9Qo07rsOUdSkyysA7eWZpg64d5n/3oUyepBbr1gfg+Lva4YaN+plkIrwSUppIgNIbSXkoky
NBkXIUMrx/yRNslebTZTOvcDdhAziFFJG0X71WrlG/bxlUxNQQwhkxTt9FJNcHPiGmqzSC0va40C
1oumQuJUl6OxvTrwCfnPaNoGq1jS1emu21ZSo29ki5w6CQJR1BxXnWsreFl3/pcKggScPXkp6PMK
pag/Nv2Nb7HFpRl4hgKq0GinSHIlfmOVv3YRrvqmUg7T93IZBodijx370Y5RzUhASl+/FT4NwKyl
ydAyUKK3nbT2Xx/a0fAn0mQBgAeAb/T8fmbHWU8EgNcy/UyHUZMuFBWnA4xKSJmBfYWZmWhOLVG/
KHp/S+bfqZEKElkk0UTDUAc5d4iXQhVyDAZWs3Ay3IX9o4c9vI5OwZWwcAHepY/qePFzkpdTFve8
vv2D+OWzPVmq8Eurd70dZoHWvUrHv0gfWh+4e/KdFhFtGt6uMSQnML8Qr4doRN4GvLREM/eYBg6i
n1Q/kBGPK4W3knFnLV9k586lQ5lxP4kGTBSR9xrFqvSItMWzEBGemcA7iVnfBSNuhHzqNPHyEC+O
0jnFoeptJWVunQXouplizwCFXJUAncOx+/xlNSdZKBUZhaxyHHKOrsaYYi6RlDnB5K8rqW/xvRku
WRU53awleu4cc+qmi/dT3eBjjS/PNucC+rrBnWeiFjyLhexTXt0u7xBmtTtewlO6HnfGxdqcq4IS
0xwymkM3abLfOI79WD1GK0OZR6wFHRpUcT7iAPOsaI0FGjivrBe13AlAuNmKD18qfOfeW0Q28usZ
fIesiVPRkEA+uyYDE2iBvMkHPcURIRpFFUZVR2pdlFSj588smSxK950A0/3oX1OeDV3lOsi4IX+i
a5leQlsiAxPcNZlU/HHFCUBw4NgpVQ3aIZlbbbCx6fJEaswaxi+XGhQ/k/NMDG6LjUIDltdCqr5j
3+okujI3ZPV9oyxXqZlHL8tZiFqxzQAvJDydWU3n9tBBLPHqJ05XESLCl4duEGiCM26WKzVWyYiV
PyOwxOJiHgxoRh23d2UiYcunZiVL8gcZ4HTpbQmW7kr+SkoBCLhLwY3ynnx4o44qTCj4dPD8QvkF
CiVDzJ20KrjZpnoHT8r2jMxzUMcYb0fnz3pX1w58OysTquCmUHUhnxeBUyTxX0f7nlD4c1rTEViy
+OfTRQTLk0mL6JhhHBxVflngffZZUPWQjKcEcIFt9FPhEs+YNeL3QPYVIOVDofo0gubY7Injqqvc
Aj+FQvBjRklujdrXxGvCJIeywM2uSTglFkuCThOqEsDFT2a9EIs95MMufSLO4ykf/t6DsRBYb3ZI
yhuUsGqj+36BubBbgxWDN/OOdzaFQicKe7VXc5PQLMeEvw7HdcyS6AMs3tZhuY6a28Rx4Gtd3sHq
N7YpQ7LtKUOpcersOFaulkjBb7ic7MsFsGLp4T9mgt/tGTQunQuGY/aZqG9rIFpPM2M/WBCuGmM6
hFMmH2kdX1SY/VPOb2U56cPZ/mHyoI7B3E2WRJQ/ptm+pWUuQkEJq3kdSS50Fn2XR1T5hV2VheH9
wr3s039WX8Mzb68dnoyHGfUzJmTvr4sJCkGAdavDp3UOLm0AeXtcPIuQpMwJFq+Xzy/ajWiKuUbG
i+tA8Ul4K34MEI/P3vxQk28VwUqlLIaMx0hrqkOKvEMuzS0+OhU4+yIhsw1Zj3cMG+RaXH4zS0CC
Ac5aOr5VlnmJC3ShJeGSvHZucvfMHzkw3S2ibVS4rQzFSrYvUJuPS1trStUCJZPSK2yMqjAcetod
b8F0R+uzuZGvZeSR7sjiWDMhspulQnTX7WRlUFHC6I6OkAw+dSgn1oUTV3E6nCPtSj/NbeE6pvTe
pHIRGCZIJRNHaCvi8CRqHrhPWPagFdOgBmqB+gVfGlEoArdegfsOG8wnNII4u9MvfnTFePNXdPio
EXD/0rEwCnF2LjPNJF7b/GvPQOFUfqplm7GFSD0rzMSCB2Tz2+0yQ7oRRsoVoQPvUL7TAQSiTjxA
20MZPFSNFiG8+0XsSBl4jxtGg4I0WC9u0LyR9CkmZnrdCBUJeYv3nQLsOBI0vsHSSoIqn+u/bvIN
PGSblzisOPihVc5uUwQAcle/r57hI+Rpu2B2j1ur6if/pcQguz2wh/knJVeX/YbuIdilFFcywhNP
G0RwYf6fcj9kdA4COb9o9gm1m16ouLBGWtAxpngDNxCMMspOojKfpQGSHTdqnHfdShxt+M3h/1Su
ZkYMkDnVlFMS4xH248nQ+sAMr4Q+Gsfwcl/4ARWUPoc09OG3/gZ+s2PYSnLl2xgd9Chrk8qLwY4g
T8CCMUemVWRYJhRU7+4phUmNi42MSVGBiQoMfHus0o+0VC2+azdmCIWWcnc5MbNLpFch/gNrhkc3
55weaq9G9x2qh30QWqlGahxOuxIdBic8ZC9sENqKi3redRMq0xVNldv+1rAXAynEhjKpOT8P314P
71my+c5Zw3C3vRak+cxwVqPhVpiU2ps2GataxbIDQDJfrEk8WoDTVWws+CiuPO1SiWkpFA76/gus
eSfSBnysbpvc17+5ajC7/N3++7QypV48wYB/FTm8NZYvhtvVScARy7qo7KTRji7BeeNu88NqWw40
5MIQ3u88zr+8pflN2rY4WCqizHVNT9kZwSi8ZLLlmt4xn9knUFHslnD80f0AD4tWIWuUoagVdL2+
EPZTUpD3iSeYC64IcO+kv5QAk13kPRSlxlQJe520Mc0Khj2eHoQ2ETz7tdszm2dHOY6qRCNiwCfb
ZGVwJEaTSIFuBMeCOlcCX4g9Y+zvfMDkTBoTxEtmv4MOysaqm0n9AEqHGkl3oyJvbAYdvHuH/3QK
s5niUdmCBaHwReXE4elBrX9EEpmLxipm1kaota9KDNllVZi63hiphM8cezdd0TR2sSekdt37iAZI
HXRxmu7VFX9YjD4AFIFl5uUsOoS3HI5EoNmg4QKMHLf2lVIcElDxUW311XL46Qxb33F8WLmbKDFR
2BfMiS5rKmtXGUe3y8DT/uH8EdItdHwx7+c0YJWP9Cew4GoOb/yKWo6P8Cd45cJXYfstHcNTIsKj
mJaph3RAIKaRBzF8cxNYbPYREwaxp/p9xmypGhbLMCFHrCqzA7hnjW3qq5liXlRReENUPGS1iMBy
mC3gHdFzGLvicbsUkl0OGB52O4yn/dbhc2Kch4xT1lHa5Ffcwvy5NUwKdX4DcGlyXEJhF3244KwB
gjJSxpntcruUaTUfLndjioaOHFnE/JqgrO4TYuDPE8UhGdUcELSSgZ06boHdpoCMkIQvUdHmaFxG
PEMwHJ4cQ3cUjzCS6qCaNeJDs6WIdm7Y9/KBoxM4/GXAHwrN7JXEvMt5RWfmuuyJXs1HwHOvpVBM
2LZCohC6fAC63hNzgrIshcd5EtsAdZzGDkL8TZxLRUdHhjeJvUZZPT2ERSjGGi/ihlBW6//065tE
mDJJjosP2qPo/+9Ht/IlUtmNEqvIGbX/0pSxQYOPJpRD1+TxJFB0sg9taA1yl7K75QQ9qy6ygUNc
Nbxrmy7Vf6BCaGG3KxTfVjSy38vjBT6bUoVikAMpQrYH6ZDAfDDNCSIiEH3fms+aEkkJA0E6cPQb
cdb6M4oMOJftklCf02O2kt4+ZK/xvjlU3Eld2CqWr2OmvS97aj3JfZk+1YdffA10hhKCPiYiU7S7
iaeoiwUCeQXj/qX6OwVYdyD+RQH/OVGt51G20Q8UPYrmqB16mBUMi3iKzSf+NKwf96lN1PTRKNSx
UEaHDL31UkEPYUSS875X9Ga589gYE3eNGh5wSovjT1GgQxM3jVkcjANT9SUbymEmuOrzaHwJoMqm
YWjtAUCphGdBiQ84vihW/VbwI4ZppFs0kTw+OdR4sn4drK3f0rTqkPr2i05+ZzMMeV9emTLPT264
EVjPKKXsgUxRMDYBk/+aoFCTuFayXJQKzAchxgRHt6HT3iLLSUal74I2Z+j2SPAwXRdQZYlj9D5K
FRZTGSpk2jSi0Tyfdn5lls8/k5D6uUxxK2X12oqCXXAkcUWYT+5Foheyzu02rcYt03pZfs/wc0IB
NvVijqauiQKdQHPfZ99YWCzPaTpmuyZT9Dxe4KETQ+deAS++CI0SObdKvAQjdv1i9po2xzvo9axY
uYKjo1mziMQZo8IZaWtvwWgJvczFrhm4QmeLJOBx25BX2E13nYdGC1hEjzy4TuVHPPpqqAdgTN3v
PoX+9qAQgM5mqO/PTcxsvO4s5Chp5doqPehFr6FdeC1msHBYP92f3kS6k0RVNS+F1gkegQHzJnzj
pYqH8jB2iM4A5zsj7xNGQdNxXhaxpeiM25m1f0gVZ0zThE1sG5UFymloKSdU+ibmcdM+BUq5BGGH
Bp6Q9hEzOLWA3Gfi1DyKmqjHm1/vO6RpftKmIvcZsHrT9jVtwjpy54Hk9Bp3swpI4udhFOk2BdFH
MVHUZxwwPRTL4LxcY2qe0kP9nZQ3xkZEHgaT9ls5T+2TBD5vr/9q7fiSBpe7IYume+lPFKxhhq1U
uwFaurRr1vlPjr6Sn6IFbdZLQcJAf6ElG7wQZfexiK/MyLhYZyC6XxEVv3LICrPehw+8gANtMubM
1+525fzHfK3zs0Ue3/qdeSTHdMmTxVQFZ9rdZmPtJxrmSGqjE72Ok2cbxputvyI9pJ8kb/4GnVmC
Dc9Up6ocLdnjAZZHMHRPsorLC7pIvh83dclgYE7O77gd50PyylQoslGLAuQGYHX5yo+0o3jQPnUr
Jn4i8l+cvzdkntldJZzZTWsfu93ZRJ4JquDZiWa9JfiMfVKgLfEsGBvfQuE+iQuKlpsno14klRxQ
Uk8LewaOEuf6eVP1eddmUq6v7JN24Z9/2zp2wY4kXInfV9W74cRfUAGnOmeqy86JA0NPxjoUJoAx
xFrrKyuD1H5WEr5RVXZeyPbPi8/KjY+7wSSMqQ/s7x3ixFOZME3giW3fcglvc/FciD3p8lgSrheh
f7HAYNfCATLCkTiFrY4rRY2JA/2wx6Lc8peeA+Wsl3/Tv7y86UQEVYNdo5pBmGKvEzMB4DQbmDG2
nIssBwKdqzkGImWAF7z4yZfottQM53Flt9Ib15QyxeKboCV0rAk46BULORBPNlWoF+yvT5FjXT//
yk/xPntSGc64SQUtAqATwC2orBDf9Mw54HIsXhbeCKOLKTJSimwCxFHMfszg2lCp76Ykbq145Rpw
zSf7kSQQg7cD+3UlOqMz6zX2Ev/ewPOUS6eDIfq3yeb2IaDWqZeMokkwZ9j/TaXLpFREfnqClIDG
GRRTIYJe86nWOC2OvxqeZIAFfmVNiJ+j5Hn2PI4gBYnsJeXTRbrQPaR1mSzCF+IjjmUtib8QLbw2
X2E3GqUVcx7fELvcfCwO5xzqsFhqwdAfDBhibg0lUJ+/ZJUrdUY3yQeG7t9j87YqetbkPjtEdhnE
bWEE45EgIEPHpfZkx2tQLFFxD98ImNuAs38V7fj4HMrDeGUmW8GcrZVXCvrtp7N4D0rm0BVtWjff
JYQ0ZP8xbLjBnmqI7L3Ex4/YVNOQqD5gkKS4HTXCpc42mdOIF7G9kVpMY7yHNafNY/OIWMRmlV0C
OKB+13WwQ/H0kBDwnmjWyLBCjYL3sMlLbP2AH0Jfa9PfYnREQvRN/sEppYZj22jE+qfZP4U0kkLz
R0IVcoF0UotSC7S9Clw1WYUq9MNstRzRVCHxv27eZYRvNY/OtJv/eRRMA37WZEsREpxWMLExQp1e
S5RUmPOxjbbofDA9r+m3TeHdlrU7g42bTf9NJ1uwYj9ATyvFriWnlJu6xpOTCTuJAyeGMXHYYhwt
/17BlmNGDixfMYf8wCdokcnHYgnZw7RB1zAB3+zxgr+kMg4QmM39ttGRgB/5std7k2UJRVJM9ASR
JhcpE3A/E/qRxDpqjASlT1VTlkSnUeZz+K2MPeBgJ2K+icJpUz86i/p1dsSeQt59cZ9gXM1RFcZa
fpPrpqK6E6ULO/Y0KpfWBDLy5q9pi/9NiuID5A/UQTS5o0A9DcViNalfEcSG2PGHmrRmm8OMy7xa
M4qvuhG+h6f6igBy18EoIsekvnE3l4rfXsEC/YiyoNVYmqvcIU5OlmJi47zZYJCNrhL7ESPSCTwa
QuV0bbzeMebhBkw5FwrQwIajzfeBU4JJ8vwJF+7lCLYAzkwvqwTG9qTx8RXoJ/zFnjrS/lCaXDDY
SUooF+9ttN2osc1NhyzKF8o7XUXO3OPdnoQRwr5pmHo4e7Cc8kaNktObNods/khQ+iSzszJi+40w
z4c9yXQU/eEcwXOlIzCKuWTgCNxQpx9TIeD23EyDW4VWBjWDIkkwPsVLsste4qHGYCdK68GjWG6x
ON3e9xC09WEHBZTcrOSvy/1YlFsS0nTr5LbJlXRpMAUOxR8iw7ySYDI47GApmv4etTHsxZBhZrFI
ibu2j6kGg3F1oqvUSBwK87e4B0mBc8tFMOZAklEIcexm8J6VmJETeH0lcknb3l1xTI8rWagEV4K7
UNDMca3fV6RjaVe00+lxO1wgplXFHtuHB2caB/DoPBmuATE8uwwgwLd/5UHDxRpGPlKBNqcZMs+s
2PuHoMUN8Vc8z1viXH8VQAzBoHMcub+LXfSEi+dmctYBRttJfTzlM98hTI4FrTJXFoHgh8+BNSGg
RG6Tt7RxNDT+l51UDoD/eqPyXrwq07cjBEP7IFvaxxclMF2cPAqk+lMElMTgF6aSu5X6UzDakPCE
D5iUk03UFr/DLEqoBbceAGGr21IRtkoXH0w7WASGCkk1lmd6KIzpCNGg1Z6FbETX79WhMFyeACHt
8RmSgFnnUNWx/f+sDBmrtwQwN9CBKBxM3m6iAFkmmnwrN9I8CCTT1GI0U4KjqWPv4txhWXf4IpQR
bmVeasOQ9XDaoC1xDm0y2E/voHzqcnaJ2AoFLEk4VLykxQpyu8SGRd/j6dhTuvLJDXwdFT0zZJYF
SDCSWaE4/1dI3pBrVTQn5No6dyNOLniWidzGmcnijGar4A4Zleg4XQrsXfntHQ6P9I5+dmbzY12w
1cfMVssQIN4ocyHj1LXFjfrc4uILLFTGT/QE1ROTivGeHc2qgkuALM081173zThZt7iwGvY+YEVP
2lifMh/AYBYcEnxvVV4Ta95GTeouzUIPUCsIMMUpMRHrDVKVs/icj2Sj3YQN+mVk9Lm0NJ7w81Ck
dyJiPT19cd1iLv32hUPl+YScxthFQMVLULTyivx61RAiKQEHdS+zodeft7AZPLdicM+LQy70pN8y
LH65J0v61e5zEnxzRc4TimV/yeuHSfJ6zZcA78Sqj/j4YP1uf/1C0xv/dkQD3pexxKuvZaSYqKvA
x+8NL7wq7WpFXJ13vqxm/xZP30/sPiyQjrvUiQ1zzbWy63e5sP9wN/xHVFeSxBntju9BLvhwE+gH
r+g4CiEpdAPOBUfiFZ6cY4OT4/oDbacKdE5wUoz/yBowP0ODO9qZKjb1rFK/zb4EX1QNYWK30ved
UXaqV/sQng3SoX/p85/Lr0tzhZImyambI4GoU/NZL+Yei2XNSklfjTbj1KYoqv5+8KSb5cx0KU+q
YH27OvMVxw4N9ogvxSyS3rTBSPRRdmekhU81xPmyKFD4FRbHRCOnDmLSSqx0DFTHyd73xNgViNrB
PsjQWiG2D1tuLBA8i8soEaO/7WeXUsKfliPAdxVNkBPC+2sIbZC1foQfL8K56G/0mumKx/AXE3lh
M42ewi3D8EIK87sWNJkwXlUI3zXjjCZ3/WH464KMi0xsIglF5YvswsHZ/bz0eHOrSSeUmD6FwiFO
KWNHVUjoOnKh4w+Tm7Y6SjzXf/RRC64f91W/HXf2RBjxBY7yjRDlfqNsm7sCSS3NaznxiQ09qR9k
8Il9+XdSEgL7nyRFLoKkOVWS+g4trFejMale/bquJDaiJ+JSEdAxe/Kq2wgsmQXpfMK/NPhfttB7
qa4zzNfaLxZ5RAUE0aILXujcNXh+6lvpZHpvGmRJd4VjqoLVcv0LHaxJxukP2MjIX6AlwYaClSBj
kyrf2TwIoRkVkx1gefdfQXel/YzjoDScx+gTcKanimr/jrSX1WSIHzjGMlSlngymKSvGcSMAHa/I
0wOZjwcRL4Ks36Ufuo2K9To1viJkQEhKKLS73DiFiEGEtMtS3d7f1sUR0evyp5Jc5PZrIfevn5eZ
ojDAN8LZTduxOVub4OLLw4vtOrJ1h/uI80eDVrdfK/BNbc4ec3Q4omNoX4fi/LWRwHx+f2OtNmZM
02Oyo1ke7ph6Sw+DZLAvDVWW6KYcSEj0BIkDl/ZEZqjC+P4g9TlJXw1/aDOoukoCyxAaXJt8FNPQ
wg3AzCZ3adYnN4N3Wezgp2BK5CFkOW1YKGt86Azj0bYlfhH9qmzzqyWNGv68sHW7PNeVMJwIA2q8
J5Lohfz3I5DSJm/lobtN1u2OPoEKwJbOSiABjZr0tK8Dg0lMH9EMDXfd8vZ4wRUTzK4ynAJA1N4q
5s1UdDxJ7HlmvUe2AigH55qbru4w5nWH81dnj++jYyf2kNI0j72tPAMUP5MVe10F7rRHBVNO4u9+
8PxIngrq5luYoiVhohBoqO8yFX6BEUyHYlI1G08/9/GmBotK/hQm2F5M8XdlIFfAVpAP1z7miX6b
+jijV/RpOJa+WOasOTvH9k6iEmk6pMk/cDL1qMuj8uEKRgTR3cZ0sZTWWX+CndSZaE47DloIe2Et
e2MkvWEfJogSIP4gzjaxpN+WGy5RcDtiH1LcvAsmQTfN4wgPKQOxu2vwdcloV5oX2FQSN2lHOYS3
GIfnVibQ3qQXkOItsLPsG07G0qQXT3SpK2IDqiut1xDUz2ua0NRnzV4dL51jZMSnyPKbljc5oJ5S
4y2CFe2JBj/cS4wniyLAFAJSWoWqBtwrtYQZvG4HrzfmmokojIuhFkCT8ooetUVeR0NiNtX/4weQ
80LJWV2Wq0ufAeovRkQkREsG7/dHjyPJvA8rMB7oF66RmCKsI0Ku1Zmtco1cTZe8rCGc5ke0iUEa
FBmuJWybksBFdrkv3aaUKM751gt+lrL9E/dAErwdzqIKPsyaz+DDg+v/brtKWgASggdb4d245W9A
eMY69fKMSMNn2R/1h4fE43qGauKJ3E6vOqd67jcCCRon8ztnsco/0qxtDDzgGFB3HQfH44UJ9yuB
WbNYj+nnA6124b1Frpt1zMqkcLeJg5W/O0sz/otR7HZ7+JIAhneCrNE/1csEvsPiXeqt7qE1PY1Q
ioGSaCl7pcpufza7CG/Xywqm/mtZiHG73M8O55gkyretB85KmvZ6tSCdK5GVTX6zcj5y3RL+uvS6
jbIrswYgR7zhmruurOppK8G2pyfPk+bXZaawAXulV97vi0Ws8DS9fqYop5I4OJfGlq3itoQNefuy
bqTqw5qxX/UBHzEiqxkzb2WK+xyTwodLw2HI8/iCM8Bl3VbJ8N5Zu3KGf97/TScuErnbYjnciypZ
YfvxTqoh/RajSPOwhP4Sgl98SN7YM/mX+MOs5k2nGVPiBjr7zVtFI1WgPyJ2GngZOvZKAq3+wncx
oC3E+6hmL7gvgADnEqLsYwGgVj1VaJdvqpR7Rqy65SkhNbmrMEhtjGe1ky1IRWXCH48lfADg7LYK
WtgQ22majL4fptwnDtLTlzpeT51eHhk2vGN5X/35i2pnE7wVTBD5yygBz3kMQ027Qs8nG47mYa0Z
NhN4wpApxeVNDO1tZtbzAynPT/OTgF+jeG/YfYTlZ4eA7qEgg/Ep2ILx+IDput7PZShvWGX8xceH
dfQpnm22VSmu/Jo7vCHYZs5uxcgXEogWSZHAnRDY78rERO5l9nylOZIbAz4CNLCFYVndRCf5XLcy
OB1ehJqEt7EHExdJfLDlKd4nr3gq7IDkULJWBWkt91cLQwgdqXzq68/CSyu8DfW4THAdGj9DWoky
NN9WOCae65hR0yn9yfzjSFRxQUt6ZX5C4dcJMBYqfXXHNjGUAFjcSe9QZ+e55th5nNR6sH40MxBH
TFMnaM3RISuXlbtIVeWKXBogO6lepO06X7RDUKSE3HdoHKjswIFu9oP68ccmBq7gG1nNUHY+rBJg
+wlsu6m6zNxe2Ny4SAGG3sarDYqckgyUsAk5gvU/FqGqjaBTSPjzIWZdGhwnaXR99r9YE4lUpAmJ
KEBR4alUOmuLKpPoZGFq6p/7Z6YuARHtw45RO2pMJL8IqV3l7+6k4RL+UcA/B7e5rPcC0HIpnWM4
iWALKT8clN3R72kqUjCFk0w36e63cAOqutBXJk2KbQff9ZK1LLsbJz/cFyHvl0ezNW9xF16b9G7F
o4Yu0J0yxApFbjThacIWxRUPlIgPZj2yoaDfjNkrEBRRbMykj8f6SeLisnuqlS0jiNmDexdCyodj
d1uHZ8dueUZZMcnwCXtp/3Q/XvuK3uSBq5TDlLgwI5vlLUXIJEjC9QjVyWKW2VDtgy2dhenPm3Q1
hxzFtff3hkzmCQUJia7NJuOgezqfsAX28HymZTkwYl7CZT7qmj93zGGMUAasJNs9M177Mq2PCcMd
ixuhswN9FUJ192O9h1Pfajqz/gWmEQqA19FZSr7eiYu9gPyihZAnePnV04IFaZjVwUvPtloHmoRy
HX5FGRZ4M3A+h9/JXKivz/WQT2dXb3CpgcUmt0EWkz/7L0lTXCQYJJroeByJhXFNMSPZ9a6tWD1g
bZaUbkXULbh0dC82tRrpgq2ZNaH11yKAX7BXTBm2rCBN1AcvBaWRSNKv62HA/7bghErC3hJo5VBA
CFO1VeH/LIZiSdm4MRA6DU7xVVRh+cJvocMo0Ac+/eKDZk29hYAp3QJlDyCJzPi4WnTklh3+wsRI
phyaPMbaSvSqRkcIGuGcfmLs7dHmU1ZGZIcaOvyrsSWaCEPJM/n0/mmjlwz0dg1488AxMlLqo6Cu
KbtyHQbdEO5A3X6CIfTJRnMyyLsy/rCmwldFGkV+XDzEV7tfypGXu64znVbHyVwCfCOJwgLePIlq
LQF/Pr902fyFA5bPfIodTTb0dHekWSIz9mZoqvUs5H+7754v7bEVswH7LrIwQnvMadIUajIJuZQn
VKYatp/kEon1FnnK86LuZCKuAYwvrMfFLetTWycFdRNtTgYZpsJvSQ4Ir6fhUNJa7qa+wAGJFTVc
uSAieTtfgA/HIhh9OjyKrkkv2XYkXJfej1TOT8dEMDjwy3QmJLX12F3njI6J/QhQsXoqbEYNgFbG
b4vrBP9PR92Wgge8Erm+v1T8zP0e8PE+QtAf1APtg3mfZFAOHCerWxhj9AtZ3H9jGyd6uPKNzpNt
LPMO8L4o12Rk2DZTsePYUu3VZEijFQNHpO7drAsD6du/eSEhPsh4/3Bzjq84h7KIrAdNxdddA0h6
TjpHjAuSMR1xy35sIBTjCicwmsbNcw2NF2Y7GiUfJ4ox1eO7Yj7Zc/eMo3we+wGgk5PcMZ5L9SiY
eycaJYTTtDilnMxwRKgpCxveoh1E8sYWA57jGrHQcNCds7aQZ6BaldhEz1fB+G3FPcVHjGtL2KqP
Xhpu4/fmme10UWIItHTa71ufnEndDQ3nZRwUpqO0uTt06O63XrYTL7z6MfcyPK9pRSjK62Vu91Lf
pyx4fl1L0eozhcVaW4QIpYUXLDAtgolAPgnRFOOBM2Yu3AX/A0TijUUijI2Lcs71Nppcg2EcC+qW
Nv3Of/hmvfuB6fpCloAWzD1+iQKgCofI9YAiyNJvODxLcSu8sdqEsrrgHg+c2xd4KvCiNuOTDr9G
9kLi0CdP3phugIauupSiwC7WsVmOBlbtaDkMOIxb0VW2f5FjKebUTQA09KD/SZA5ymwaF/wsY3RC
9aG2fgThNK0G7D/nHqlvJAtsGKkfHyU5Fqyy1ORhRSIDlmZupgs1e7m2damTczYsoYVAUjINTrwX
Saz13WnLx3qw8AnFLgbJwYA0zWkczLRP2rekEbjHCmCxly4NS+moZq/qeYjvhcU/3grjrmYLo6SQ
Dia0+zxbc2HgOLvlVfZpG/MqzTy4ga9VUcSzmshwINrX+YNXf/rvaPXTC2NtLBPPaRFOW4k7EPX1
NSjsZesHXyeCl24tDSHP5fH84Yb/e+YpNW0bu1ej4doU67dBYs8neOWkDvDtuahurDmwc+RxnGGF
WAdsac9HlHp5BS3sw0EYjoDwzFCZxHIJDbAPrZcPCScMXybnCYW/0kytgbtAcR/HzEmVMKqFYfOC
0uVl2IL/oRoUMUgt3SEfSSqEFA+RHiWzEVEPQja5RGNidygPrhb/eVNTiW9/nsIzaTqmkIHp/iC2
F7suvll5dyuStrnR8F8hHMpMy4fYM/i+FhQxQaCHlyn2Q8r/IhkWSE8ILwVOiS2GAk35fUR3V4zj
v2rNF3DFtJeJYRz7I7HuemxX9PTNFlFeDYURRaNXn59jTL5ZYL0plEOb8ouXyZ6y0LcUJisLTYVs
tJjCvfkuO0xPcsCw0CKG+2ip/42ddVkBTXHcvLV/xJ/SxC9ypeAnVFhZJnw6cuZAMYJk1X3S3lU2
uuu/zxic+z2/BnsPGaeefF2e02OB0ed33FbkaBdexccuB5lTy/tpSIIs12A6vwbHsf4ZbEYWryfC
1/DEXbci4BSovTEPLlbvtISOytZqH/3bG/9ZPgxxi96CaqHjGWZ1Y25Iephicb66ECA/TeWaNahU
x5PWCjnm3/sTiiOBPjguJXybY5/PfoZ4Ze67ncHA1EX4oNjMoSl6nr05PGJQqC7HOuXmHHoKj/up
/l2BoRz7chTOx8miV6sG/AhVltwWY97i1+AP2+CLbRAWJ+7CKi4lytvsZ7tfiw8NmLRRZOxt9hr8
wqC7Ij2+YR7LiFNhnckCzAYQ47muIrj8rBn/dk8XXMpJtKxqwcIQ7C6qS2wTzpcp0rXM1uu5BU0I
tnW3SUBNxGbcp9GW+OzDEYGe4Osv/XQqdr/hxx6rOjMNRRqsxHRqKOrURNSgWDW3DU2GL9TWf+7U
OErBUqmkdNRE2zVENGkt4KY0b6+KmHYwd/Icz8RYHIPvi92hg6IybcNshnQO6g2ZVn0pFP8aepRS
k1uq0ukdRSxonOZgT6xMLhBm6eyYqfXlODpfk8JoiAEtvirLevMjuWYLoWosxYIuszz4mcX3uEPZ
gdbjZ07T/iqEwbYtfHb4Z+sn5hT6bGBibpBnppEcb0BX4P66fIyYWa96M8pGi8B3odPh4eBzIyT1
eIDECzionVmfiAyAiz/InKhZVOF+6LRTCLUxLZ1AGg/lUTFYryW2JxNKMKwT2tHVIFkqvxs1zGQj
dle0XBiNf3toeZAwOxbtOse/rZXNHHx/5GrwYIJ22tkRhYMcgYWu+no+mImSxipbUvY8LBcErWF5
dbdN7hkWZD8rO6aTyObJxznmPqqpHfNrVdLT4Jt3Mx9hqjesc20Zq6c/6tFc9+6z6nnodnnx6k2h
Pvr67xYD0rizb6N9IIhRT7747Ci7cPjpiYZxwjD6iU/t/nEfiPeaR+/oqdZ75i2TMFBW1CeBbSxC
7mNedmuNXHrBPUkPr3YqxZmzBu4AjJKQQrsPPYduwixtTUGHe7DuaaefjNFL1Pw7cp2bs7pQ65Fy
IHTdEmMca+og7KlhjnxFDBgww8Tm+oTPzjos0uZVBImYkGE9AHjHAS/kuOiXS5+iq7Hvsk3fKwVC
3blIU2vy27uBPxdagFf/9XRXsrnB/vG2VaXjWbM+tjQ4mbSKUDWzGAf4aqkm88IaWh1j9qjbLLnz
spZQUczfyyNO45TGSeY8k4sn+G2L15iRF/Aj091fi90YdkdCW/ebGhkawYBX9SZbgTtBHYskPsdT
BA2skqx1cD+QomZRXeDBcyzdl2qS5Pc196mvoUTrGl+VqUw0YY1nfN57b4tSTKe3M5TmdOzokc/P
tNEHQtFZN1sDyGPD4AyWTA+guyaLgHc0+faOmIm+lI7npTQPIncYdQE0QoFhGnsKlQ77oA0ABJLe
IEzsOB42R9uFlswbjUJd5Cil7YhhxAFHRlnDSzOiLjtS2q8JMQEVSBaB1dQobb4m/TpCI27hinWR
qamieKoIP2rOJmC71v7kqR8lmhto3gXJMDVMi31XhsQ5xTmDHnEK9EwyCA45tnYGTQOQFCPqDfQO
kR32XlFLY+/alRoyx7XJnA2RvVYekcrYEZrAzdxonDlq76PfHSzLfnSX2VJZ/PgX51s+rXc4bm/5
Oq5ZstwfoF5iX5tBScTSv0GnIPQ76mxw6WArf26JICzcwcqkmQyBsCecw012XAd+poFzZCzwt+/m
F3hzDgnlA2FEA2ok7Lm2pd8L1D8GHXGPeCQ/UrZGvN8GO9YLfin1lJkqnx9gwVXYUcFJjMo94WuN
NcSVZhX+kC17Gg9Mp80HrOfS5PcDoTdhWJF4Ia0WGxmsAP2/NZsaI9vVrt5C3JS+knAvatvpzIRV
UuGQfbhSRfVLkuPSAa8xwfkjDgb5pxGX7/bhnJ3rJyr0TavZKOJbpRR/4mHatTD7yhMcQtIGKjQ3
hLFAu2OBcvnXmP78GEO4lzk8KhJwCyejtTyWYsYx0zEI7QFHWFIUy3XXJ1XeTleeorksgDmGE2xB
PxXImcLflgJlEsuVWEg4trKZOr3eLAoIgWqQnFbOq6qAVL9XGC5+oGwp2zakVfJrpyCknY3QmjZt
IXyFYC7+XlyKRGcVCHEsRi8PTFnzrH2fuP05sZk7dTSjObiNAgPNV33/JESz9ILvftrF7qnmRg5D
cyKzhOmp5Ovz3QIFSRMehiYCiotrJtgFMW2juzYj1Cy5akhBjiWnc0i4WpFXeRt/kMkDStjZsfar
I6DQ9g3HErBvO+IbJUlieWKLvUntsgS7DmCbJHdKMoGRp/8g4o7gS/gwwhHUgJFl2X0GL79g/JCD
a06Ej+W83UsD36NhfxDTos1VUueRa1SO5yBBuaYeKTbT7rD9+sHHffTrobyGlhb85JDgzRq+/mJG
c4rfEJM/JBOcFhGe3DD23V78+RsLDX4Vf/rG2k3XLdgttmOoVJwaBh+eWqSGrh6jyj/nciY+HPQT
DSQqsk2KxmvL2BSW3etz6eWnGOteUg561qawm8R6Rt5idJnA/QKwF4sRNSCloPY8zFgyEH3A3fER
tk5SlVughb5H/FWptpR/WRIWQ7nzjIVuCmlH2XxckPoQyvg70jivwi1l+6M8CVxIozkBYfvrppSe
93GzbSwAyftZRZAisT4lhWiY3eNsxjFZxqrc7qDUFGIIvivSNDy3XN++JbrXLYx3XcUdj2BsUqRo
fLQh5d4BQQ84JvlfyKrCHEBmXJzUwj959GyiKmjK+zH2MHRmNpq+Ze86WclnOKVxQXe26SBdOZJ2
Ih92pB1mLfRmYsU7ijIzJ6J1MorqufBmhxt8VcvHYF+Jxbw7drW/fJ92ByVrMMGyxt7Mc0a+w79z
l+j+ZjtZ1BadvIj2KWsYbA3Pz61Gq9QIWPA7kBNypdMC8laZ2f1SlbDXknM44W5l7VQ1vRxhUfzl
DGnPF5uL5KbA2/SNFpObA6VMvkfNZW/zz5jUVAnYovcTvg/wi9gBamw3qhOEFGmX9FJj9nrt70ob
dPov1R4nEN5giNUJBDJaeEL76QNG8J5Dw75yhTK1zY4nCow5XDn9QPb15qgarsvowQOH9W75ScLX
S/Csd7DHZeLYq9jA0qXFiFajDwPBOhl8N3snYj9cQaIcAAiTsPsSR5yv3tQ6ZFhfLCMbbhdCfkMA
46JvVDLWnb03O0iG2Q9R4uPpqhF/9sN4FdH/+5AuBZA1dc3wmGRXXGreeomg4+e6B1mQYmLyXV8G
D8H+5yYBbWPfFBLC4gAsrFLGjUGhwzMl6gwdjM+0oOx7K3MAKSWb4inKSFBGMjOwUA6RTeSIBXYK
O8M6URKzVmUaM+Fp7i1o4phzos060WSK2S78j1QjRvRg6VTXaL8M0spnLFxcJzWq0UYo40e4yC3Q
D7sLHaQhlSVLbs8vSr3tFNOosL9VyQOaCcoar4CbIeMdJB3HxihkZq1iT3AaqK5W0M6PCKf2vRTw
qrwzxgJrEoRb0+hMb+WlG9xJhRvim5SAI+dQEgjsvsPAmHl9pwJu1QIROiCSp7lNMhUJEvR1XuWM
qPJzcmQLeuu46rdbE+T2vZNzrKSYFXlb35DrDKgIBAG21QlPMFXrV4cBa1PcrzrvUVapMxp6rq5v
tP6eksnoZ8YRV8odrhOW6JuqfApBBDkIj+Q1Er5quGFOrS7zE2gNYgWd/a6/tjffgd+RLlDMm9yw
qM3hyeag8g0IivzFMW3KHYrQD2jcCA3BVpjo9u251yzxnUq0qJ49Whnmhzq5xhA5GDYeMWSnGy5X
anT7JGgJUuD1MCr4JsgsnCZLVo/m9zWMG3kMnqc4Lk9ZCqIFBwClTsufMKUjB8huOZI/a7e9sCVx
J3DgFHV+hLSdI4q+6K3WciQb5pL65EdQtpRNjZSc44xwK3n5yqqxeX57z4Oh363K7Kpq3rUCV31C
p80irrXzDz2qgdwjcP6tOHkD2VY7lmhBfTLLgFEO7nTOR3Jgj8hod3Q066JurYJNDVBwy9SAFTN0
hdgzCKK9ijUJX1jVstWUamIb1YI3MPVaHWBcUP6UiBQ8HpW4hyrB7UJNqEVgHuphaUUR+zrpWRM4
OH2OF033P4dgG0maM4+5jbxCWVkWC4PvWYA0IBiHAe7wM1Dt4P+G35JG3e/HtF9E5H/dQzW5dI4Q
z2WSQ6opSeeR8ptQcrHO6pPo/Ui/L+wAL0XMKYJfyDEmQ4m6d2+mdCpIy8B73+MZtkM5SmfzP0ZC
cyrIiaqIkj0KTUgjtQPVuIdfm4jZavuOnW0hzoSdGNZa4yEOIjYszqNjiewWwWYty36HIzNyBKIN
X8HzbiZUs3J5t3EK2LE+C7cP/DOi7hetEGhrXGk8f4dFYUVi+z9M8hpdd4WADG3jxTVrzEVSiXLY
Be67xw4A9jn6ZOI1v3hGL22MoDuBujQed6/Yv1uyNUVIcSjQPRtRcLPW6XgFs34U3B/Tx/S6nC8o
oDr5vBz4Dfnn3AQUrLqBrz0zQELYexfovioHylUF4ZzYH6mHGd/z3AiPbPU5yu1XFOZvzKEgcfoa
U8xriOYix2VZMXOLGh8bTkOQtbZvXs7U3JkzU1YHH/m0mI9FjrL/b0fO8qfV+2t5AjQoCaifNlpo
x3+s2GrqAVQzJh76amqDzrEc7OeclKhNfOL9mgV3DCR7IVH7tJAxJNCLRjRh7VDZiHpMz0XTClWv
nCpI4rRilvbpvO94rmQbLjmOMuCywFNxeQ9jcEs/9EV+w9i5W/afEeXh81sng/TC+rcpds5Yx6CT
mYYLehreOOzrlgeVdzTqmjLQA8duXPgf+d/W6pOlpNbPtEcTJEOfW1nJo6BCG3H2WkQv0mid2Kua
xog4Fups0IVxtEm8+ieY1z3Pt2whpDUmhLRsgGH7DZ9PrDFTRk+6UnDIOHDQ59rQHew6nlRUcZRA
Gfc3vuvQR5EljN0CyQ39iTnkpRIyUNWWKsWXmz1ISWvoTGtz8cAeBUnR7PoRbcrucr+x6sgvlYZx
vmuODelU27Ow2K7EwyutDP/aVQIXJwXlvwa7JeLu5tFrbgzvTYsyfZUBbci8Np1qEjiNyl4EAqAt
LJR8fWackLS2x/2akwoi7eS/qbgBXmS+2sJ7cKgUJJ1bSxMJMDZxwOvyj6FD1rk7f/guRn7hSP+e
a3J3vz86NeE1PtoekzCW9zS+fIE3skRQ/kWVY8A58XhGgKJK8nl05cXg1veiVP5ddyJjOoT8Boq8
xW9viSrNNNdY41Ken8nywK1Swa8ETxOvvd1wy+GHtFRdDi7755Aet8r4ssr61ldUX4oBhWHKszqT
qR1AAi3IuAEAdgpAUIQ7IJUYzDUV49oelWtnyruurFpXe8yFzTbd3jImJKEbD9kwQg4GtdPgE3aq
D2ZNEYYHmLu+RcylZetp9XoHSXBn4vbH1Cei4E2m5Gc3SauVr+JNc8Ou7MSE+nNSf+ehGWCRF5ku
2RXNbdV4YCvk0ZJb63ehaIBBbRaaROjg1unMAVDI6JATGRpYLogWS/hbZtevLckg5YYJtdPQFNlS
RP3gxfnMwnezANKCATqhZ9NP4PWZsr64GOZDVkLjHI9LTVLoUdEyXngkpV+31BzANYujDfLUV8Eq
wWWZ3IxaXJme6t8ox9/xXHUIPK52zaBnuV1BtdyTjunAWc3PmVbpavPJOHT7ukfp/4NVGf/d6frx
hui15LtDzQKbcEemOLJKsG7yJ3YwS33BpoLla1E133ynZxuU9eXUb2tCO+c8buurqkOFBeuf6/aj
40WCw05Fh+p+nbMoF2oCpVpAH62k9VnWMocg5TdJEZaZR97Gs9EYUOtN5JJN3Ja/sqqJw62LK/Mj
KcW4bhs+Bc0x3r+QjvQEz5u7fLpmfmSnYPXGBxOAN4T/ONjmpt6HuBm59kKFegSVCGEaRzk/HcVs
sr1heo+7l77KA42TdSBA0hvk7RvggGWDMND8D2tUgRKCcInUjdqr3u7gIQsbBPDauGVvyLDZrq6Z
lFCytSoT+uUNvZk9SvAbEb8LTwKqpYPtZBfQgMFtJDESSRVxZlRSWr+ktSFwP2fIPW+ATdYLSgdB
u6yRDbCxOj6yRGaShOybBhE58SrQLMaMQIdnFqcpA3EEFYqT62r9KaTTpc38u8Qse8mXxX+9f/yH
ksr8KOwk9+aTFyeO1xq+3JI887Nmv7mvLon9b5K7ljzuKUU8M957Re5z8Fjfp355VcTE+FZOKqDj
c1wVps8xcPbpIyRR35Yq8CIO8LCtxq8/52mzbakKHVUFN1ZaY9qQm4rR225HuFsnI/Axd0dn7Lqz
EHKNV0JAmBCduR4Eg8JDbmE5UfgJLqf/2Z9MnUG9nh9LfiKdJspi/I2VR29K/U/CzVa7E7cR2tnr
x73STWYWOgnoK6wl1Rz7xmCc3Qv4a0QNXidYAO0nnd0Lz+HP3KmhWz821lZa7ptyvpKw0IuAdIC3
c23P5JLoLYJjKhL4nYMtRtr4q/bXoVIusOOzVUl5z1JZxp08zvsiX+emMPHUZ0G8dibI8LT/7zGJ
xXWVRYLhAh7IrqhavwnRKppoFK0JRmDEXKjRrgJHaeZxmHvrUnQhXVAcQGLKdvrusjeg3qZp84d2
3yJceM/hfdnc7oT6Zmu5PSdnLhVw6I/2MGPNhA5nWofUdG0kDSflss0S5n6Tq+PyfDth8IcwVRD2
qBBOQNSewFUmusv2vRt7/6aN2Zl15xvNiixyiNwMmNTYnrWPxPv1KpbW4PlsGhQo4DRNM218rWdf
xupMMSUJilshn8TdILCvZlLMWXaHVXHb6c4XrC6A7fuQLiKwkn7eDJnHTKhKSjb5oHEEydu9UN4O
Bl9U8RoDzeOrJmvulLMauOd8uVNB6riPpyG70ZqZQTZgMa9HxZb+7c8ouAXJBSXF9c0Ouwlq+se9
HvKatJ0UOm0lkn3fS1z5uZyKVZ1LJGzza9wFtgElGkOl6sXxP+qLysJmN9zo1pvIPYUTH9hMv8Nh
yv/2oStZaYpTh3SvvbG55UG3zQo7O87ZokkrJIZnyh6KYXSMt/X755z57btDHTRLx+qAOxWiIX2x
iOC/2sRJoNlDGN9WSL1e9k/qmvS27vKhj8UUrK3ZxluU2njk9LwidCYe8p/0o+No70nu01W08gPI
oidiX4u4Imu16LUybVE4XEGtgYpXLt3LBaDrhFbYZ3ShC5V5QRNe8z5G2m0wTwc96UCs0lgnpdCT
M2MjRRMRL529xC7EyYUq130UTH6KxXcD6mForodVD4mC5mJ0VAOPdx48XiwrreyG5vrbl/UaktWQ
0tKPsVKWKHxTaogc00/KLlOtc85MnmN7IlOVo18zaFfXcqpdDWOR/ioFRyJVl762bETNtDACE5KD
Lf9V/1SzuHmbXKKS7I6xggqxjWd4puPtOf32+pm10UdvKi31AeNcBHksP5c9YrBkSIVpInyPu3/u
N09NIwI4Yr6WBL7FTkAqet3gHFcKd3DtsnIkT2mDM3zd+DZnPdq/ZY+YrLjGz6sxFXV2MJ8WMoB7
TEXe4o6k9qm0DC51KkKEBPs8uogqsE+5RgD1Mb0VSfFphjW270zLRlXf/JmSe0vqaBraPEzeR8bL
ZpeUFuCeVMEpWxCeuTixxMbOcpUjgQM2vcQ46QYGet/5HzGBndakLNUwFsiEudT3bVNs3O4wIHiv
Ol5qYo5Q0wKvuFbiuL7Ca4f2XMfU6OIwpAbkX/+Gvc75PrzdmTpWJ3dNXnYmJSYB17O+yDOvUQYS
28zu1dxe1JU4dA9knOy2PU9gpDQJ+S1gj1bz1/xG8XLdXini6OMC97/xZc5MqofSrXR7HyQXfPt3
b8zyM5ZNgt+DJjeeP9sLqBLBarFWDiFqXQUe347UstcgEYkW19U+Wg0iI+eKCrba67YoxZPwYBNC
2gwBSbN85bxmVdCrVKZlSzN7A+MexsfzGmZtt+FBhbaUcINN8h69U6NJ3oviXbTBsvf/Yz91HQp3
H9MjoDBhgQQLmvMeAqLTDsU/r8QqZf67SZww/tYQodpKR3VDG1awDx1W3uJbroPDr8Qc2OkdcioA
ykGN0JeNStRe/lDO0qBAGkOScrDN/RMH7ROsQll5mbWiMQH3ysxbt0Sn+zp/DPrq4T79NnGIFvAq
ljejc14cLmd5FgGbhmJG/A3h7svaZuF/Ceyl26Qgmx4gEI9hxBs84cCJMIewmFBKY6x7fHhzPBeG
n9Eex4Qymc5NJt/Bc5Q4t1t0WL1zXMOzj8JhhLyhiQ/eshzxYeg1xqg5Eifh1eAjzquyx2nkMtz/
R0SE2RW6Chel/6uivZnRTubbOXN/DfcyVIN5ZPl/T62X98KjuCyoLYXY06SzP9Ky3ghyY8eHVMYR
5irxwucJc+ddr91vFgho2JclKiuKQrtBp/Kt7uu21l1BOWAOgt54iY+tIJQcv0MOn0v4OE3w11BU
5MHZXuBAOAwUUlWhxNrMyEne+tw63drBFilO7JPAjb7M6gc4f5AA1obWDad3o/J326o0L8UHN3f/
T8SfVyB7ZGrteA688Vq/JWJYJK3CITks6GYnPRmLcM5oqUXnTOi4XHxfFWKmby9FbPzrWh6vQkXU
tCROZHJhEQ9E0M9IeSovJUwJ4yHEf5Be20jEAYpCzTmpS+fYz6w1WeOFI+nn/uTRUYgeqdJei+DW
0s/iemeSGYu2Lzr9UT8RoU5845vgDJ6c16RaSSz0VjKayfQHFcTGxTZXKJW1FRejurxj11mPsbU+
ESLn29+bmKIdblh7LcRJJZLjc3rOLjPWiDegbrJvVOAaQeQuSFKWTt2xzvB936o41zNRB1cgwGtc
o6YSDDnT1sCChIeO1kHAzM391MM3qHh7N89P/BsKv1Foqe1FfGUSeSLzoBpaNEiZm7a0J8oEA98Q
aEQIsjF5erPvbCasxWs+LiW8vqeKCmzrE4MR5jlBIIpC1swK3IO1Mae3FHQpiVl06d5CoIBOyxjo
gx9JnTyaBvC/zCFw+N0NkXCdvkZCKVQIb6rKjizhzckuOoWCNGJYLsDtQFzx5yy9g6F40mHzX0VL
cQO4/2lSebZaVLsvrUKUHqUcmkpK8f6oPROUKVTr1axK1ivMU4kouaQMYAspHWTC8/6/KgmNA9tf
787rkJhkFAHYmDpcqWplDcEikP4NiO+r6V9AM8zcrFqjJJqUz21A0XATfMWoPj4QL8lsvOBMaRxI
lWQi8IqVQajwC9D5msbh1q1iQzA6LA48JtAVFHJSBx9BgHty12yxBlIIpDwJynpFDExvbr2wXyZl
ITsgCAUy6HOhfgkasi+VtkGmkhFQ/3hSV+HTbK0W278+XG5KsyoTLibRObvty09zs7+SCkDrNAZX
kX+SEEOa6w53HpPo7AV2QazvF094Pv+siSSjVWJji9OGXIeJ0h1rNANoZy3FekOuOpXDW4AilvCG
Eccwrzr3HEg3Dql80HLhmIqRn1M0Pleu2WXe3zT3vi9D6TUAd2YG42m4j+x3XecyjP2rL6M5IR0v
vE4bHrGlmoLa/K3UEpVfdAKGQ3C/F/uMwJnmN6N+jsI5t33f0O8hEmByFvn91opgAXd/bDfkFFAD
7miYfer3CZedH5kfR+NPgwFHwxsFpl65bC105n6J2CFal1CdBKgwmiju5w6xi6c4+tYnD1zjCyoD
ozOrO6GZbihg4N18Gz6KSUPbzT8cAI4PDtmZt9D+X/Gt4iXhHJ/3rwk8G4NTuvOxNGzi/Lmnzd4u
lwemHPFoaVTfL32fx0uJvRyuklKD/0s/snUS+yrL0EtmX6caH/PO9MzVWbsXnDWwdaaMnh+gzifr
WnKq/zmVwJ/aj4693/5D4drjLLgp1m29J6iwtQ2wW2wF9+7M7nQC2khFGgCys8LCpghMjIZ+nzr4
LyoKYUzVJM7f1oILnfY4Nuu/jNFNT0Rct4ICKlCQklCy1V7x01mbUhjGQt5IqjPc2Etdho7Hu1KG
bfihQGA11+OinWKLhc7n4ufIKCMq8ZPTI8WVYhUgW2qV+RYd2bLXslphNoPSdJ2vdaK0ZxIiCIGR
lL381E+wHONlMjIfmmHO5thoDPRprUC3HEO01LD4mcp2592MBZhKAYPzPgY+zcFmiIazC/ynmWmx
9b3+ae1UgiBB7AwasKwwPXnF3lEv3W7i6FoX2Qv53eg6Vq+Hj0dsvtVkGfc22Mx8KTTpFIAjzxF8
UHbtqGfdjX2/SXpWaaynP2tmkJ3xUsW/zj2b4aJr/nPPVkTttxVUkHQuBavVy9bxeUKfsWGckMuz
+g+43m/9jG1a0pA5tYtnz4KdgKluLniY1384nMG/i2Tx5kroPpxYUkRwPrFAj5Dr7qt9kcvdq9Lz
rVgKdwclAPCJkJ4E054EJt7Y3trezT7m1TzOFs/zYD0YwT0P9Bg8uJ4gPJ7ZtG1J2IKWHxXPTPL5
wRRDJTr8cH0P/4ccgmUxVmYGXA9j4Ym+14vcrTMR0tp+yccDdHG+13r6O8fRqZi5+dg9nIbp1X5p
QG28iqrXR+nUYbCGq/+M/KNVJiR9l60orhpPW6rH6r5ZQ0fXgKRCnL4AWfSRXAv0UHziPvBWzUEt
M/aaxfkP1wH0Rfj/stiC34noTNi2RYxQ6mnEsfFqg5bTQOQCLhCyDHpdcCGF82Bvx3qRad0rMn7X
jOFVoNoRtEAiI5JN/ZVG7WRIPGXCQv0uJc5nBhnkssoHqllMCdJUSSRzeLwfpYRcjRwqF+J70qcR
haYXDFObfyEdWPo7w1jjN321R9oI0YLSFCA8+XnVkwvfkC/FizoyXAuazcRHGrV8UAwkrAwFZ1Mu
IHxZ2LsqFvV2RQl//8nqHekXgCrwGHY1f0jLdV5h07bGQcCn7CL3FJor+lOM4mvAJgybk8UPLh4Z
M9SdQY5u4ntF1ZGBsSdDXZjANl0lTJWWHVqrnuS1Z8dqFniuSFY0v6hHBifEnvSa3x8/FCekidq8
uH3nU93gjZh1hVwPRqWAZk6fjOSyiQIWO7T8OYPD2zaRjI1einhl5S333kViBXAjXqrZycvofTGt
7Y36eqgCi9MNZbt6kBzVbZ2oyssQC3qq49orYcsPl5+qG35rR0on4t84cGoA3s3OAFjYriqmhGf4
7w4pbynTKyH7Uja/AfCurYNn9j1RxGc++XriCwn/PijtIhZRC70URXZbCgLPc60Wz2vu4oVsWX54
T4gJS6BAgnQ5HoJIAgi5vhF2F43qGwZ+1o98WWDYi3+wbslEkLm0SPH8y73jxLCDx9L3FQmFkWK2
Qx8Ah0BG1ogzczuwXEVXd3aULmEL7nGmVn0U9WE4YWB3LQTQSe45WLmUuTP3Vo1gH6aDCOGgYUoB
6l46vTdF5MruJrwUwFsSZVxw95v1XPDA66zNNJA3dcoNUggImNhqLWu9tfHVBjbtH/hB5Hr4d65z
6oVCq/7ifyqAbkL1J3Ov9JUI/D4uqMsf5+UwwLAz+SOY+weHMI6qtVZ3cAwVDOYlsjTJJAmEfOK6
RQnkuqMrERkPepeFJTJcsVZDuiZ7PgfUZOd+qc9foCCLle5mzZ+5mLu97rhlsE0hXLCzUtRzIuuP
dMgFw/KgDmWdajLcH4i1EBG60Du8FC7dAP+4jG0xx40VbU6H6SGcEn6C8oFsIFX+H+uFVV8p80he
YALWe4zrcS69tFxrJC0RVfmiibWDd+Ldxlz9iHD012OMSOb7H4gDOUTj5votUWA2m1yqSN9R0AIt
29zcD1IHO7nJUAJTEVtOQMw32sTqt8ysSOf+gSwcUImf3AEDrQRKfVz41DeLJGrq+CcN2s7929lY
R8PK/iBv38LX/iJarqirUwDD6D3YeTle9M6cbSvdC6LWpwOJcvnxwgUN7YcFKJwST7dEZShgYvyC
a1cyh0KqTkp7zZTCB4glNVf9LQX97KwvZIazwsd6swBadDMwQWdeMIr0R9GaAhWpEI23Z69PlR8W
x1iI2Ut/ZpC9Llu8Rd0pRjnYgkJ0oh5Y6Q99+elL3UZBBGWPHwMwpteGLAZmcAeOJ9WX17ekz+Tj
6e7AaYzpSy2LYfFIT9IKAdtC+fmMxdM/Jjg/zcX4dyaCHNFw5rmbu+QeZTPmJ5zuvxbgzA+lz1V1
DLxrgmd0X4ax9asRbjVRMfJ1noAZ3PBU++MrgKvYDXy8Qg+FxdHJnLgJS6cxALhcP4/uXGU49Tbi
Gh5K/V8JqNfVGN+tE7fgyOhGae9DR8i6PwYSxsOVGbmtm5VUgtyFM/zIFLEi6O+HnYuv4sroNDVC
XRDGVt41GrPxy9F2GAESS0FI5TuhduHL2rdW6wpvXcP3WIFZxw+WeaE0qvsUOzO/GsCGhyF/Da9x
BcCDddq+R0V9T0rDyrZIeLGueTkCtkvCWE4QRuxRgatsmtvQ4Hm7uMURH74q5+Z0XMvYdJjX0Ht5
EG7h4nOCDabINIDCQru2ZA6w2doJY3S0pA6es6HrOrOa4BBKFGNxF9+rvu4jZdwNq0szcH+1wlm3
fTlPoxFnrJiWKlWsaBRXel1P0YApnYVB4mUA9NuR7RSLkVu6yAyHGTYvxj5V9HtpwQcxWU/xczAy
q33mAhdEgOuTqd0Lh6cBsRiHKkgFE0XEGYWCQCgdr5/eKV6UzIr7lK+bK/TsPckFOTGmyt3ogn35
JXnLwdz9oiJ7ZAxunY1fPLrBqwqIITLdEmFbzoapDeFsFi+Pp00nunMg93pBMSirrh5y/L2z/5Wy
GmtV8rT3NZFFE+sO6F80pFVNXIfMEHMzPy7Jp59lQZ0ToJqLBKFPAsvS9uydXcdpLnFDFJq+a5gW
LOWCV0E/K2g0XkXcRgYC5Wn2H8Mlfk+t2F1ye0zqDbcMg+FXsurlSTNvthTDMAri/lg85WK2Epan
I4AbpayzBuMDokCg/NkibdXv0il5rg4RKhrHEaszkR97yjOHrWPwIpG6kPanuz2fgaOD2SMeYV5m
J0vaaSKcOta7BokVV2Hl1dVtDPc1CSyFNodbDCYpc0U2bIHxWw9RDbuZY9b7uT1wMS5o7FBBxH4b
JiYEj5rALihFBA6wpbpRwOChzZcl+swiAb6Kounw9u3gdQ9pCLEH0cTAnFtFGVo3nz0z74Npfw9s
VCEXhPJfTYeNaR16WlAUB4V4vjVQr1Yk4KsPkQ/yA4+0mx01BxSN3L8xl1/OCjEwdCIuIh/jbZid
tz/E0RBGdQpaK/AP72AEUfJ58lg6O17plBYuQu5o2G3aPVGdVKKmauvyrlDnmJOJIG3TygcJIq2l
EexPG5LcVkVrWZ9h/4tmlbCLKzj5LyOHw/hB3XA2mHwxv7HDWC5+SIQ3Uuvo3C9e+CysjnJ0j65Q
DMomLcP0imHJm/gzNcqDrr6VT+too+Rrg8b8I2ZDXl1XVBgEf7Pjpqo7giGlwd21FbvA0omc8BhZ
DizYrn0rrkPiOLNf1oomG16ejjhOD4LuH/V28U/p28QzS4RPPb6yZawLagzbqzNJM2b1mB6585hr
Wb9O4P5N8Zej8eV1RAzfdLt4BOdk+AlzGFednirudBRD6AMrAfXHNKWL4z3DRiu25fE6X9SEyfzO
ScfOFiA1BNUkISH2U9riPDsOJ8y4zbGMFiuW95mJgujLq3ZHTbP7c8xTSB2tF7k6bRYbdmved6b3
s00e2UMFQKTlbR6/pvkDrArcqlWwFjivDT4cmZtZFKRxPSvvW+YbI82oH+FMWm/XTonve6BMuNAq
h/egF6aH1nf8CagdernDxWhktFEvvcdrjffXLtTKgC2S4Tp5xoaCbO9MfDc26RQ69b+NR3yrPx1V
j/YGbnMkYrKyiygflp963s8vzyqzIoh8lqpnzf/wr6v75FUFbQAZi24dRTQZg3eh0EC54EwIyl56
HYTMYLLsMrEjZuJKZQjEL0D25oP4c3GWHaFuYBE4tJLDBc9Ow7aXzfFYWlZnBUnA3kWFExVQSvxc
UliKyQMEuuwFY99I821EXlZLgdNEE518KjQD3C7RBpN3Upqk8e2iQyJA5Vhec0iPeSbwo5DVCgzu
lzu4zVmEcfaQvDxSkjokJaX3wxxGm2tqSjYv2RcgTz6Io0sIRkJrJ/ZBNms4S5r8Pr3IIY1fxyl/
BdGNUSgqU9d4npDzIR0UEINTfo/L/TWyYXMjHH41EtJC15KT92Fn18L7sVhw5CPJyuvXgf5QXsQ4
xEnxn8UbRCVyCaUgPepR1yyGbpgCPGZ4GJqI6RHBjZHcKzQzhjVBURI4qpcfRWj8VfNvzboE06Lw
GvLctkNnIvB4RTAJG4gi90Wmw1bYAabdXeyYps2sInhfHf5pDMoJ6kFm4Pyg1bMZBewXWjfeIIlZ
FlfPb5wh2m9O0ClTpWIsvw9iKhcHLdZG/Il91TZv0cPeHbdaXTy+Mq2Y7gnUb9+cXfeClJlXKOZE
+XNmef10T308aVBID1oaDYb75SfwqYuv861DTm956bA1TmVbz4Ukk2J+0yiK9MKhgP8jKdxOKP5d
ldJshtWUkDqLEuDCXj/LenkSTazvJzGOiT0BsdwFuUgYB6KeuAA7LK6YYW7Y8A4PNm4p5WecCw+T
CkDxWI36dLgHDEL390TyPiWkiAczslATdHoWv55S8qdv/aipxdGYjHKhRZO69YWIsML0r2acn1Up
CJHiPEVP+RCzBKQggL/TJroj5B1ceO+ebXujIJyoauAEk6ZGpcA2nGHnSVUzpVPhzPjwtTH7d+CN
MgSvyENm/oin6OyIM8fV6D5w2yK4jV3uWMrMDXEwyiFXx3rvGhjapwg4VoPmAQv8O0smuGnk2xCl
Pugkm7odrRz8SpPmVAzo1QlPOlp37iAglQWCVG+Vu0S3ssTLGm7IAobPshFQEaSMdqnmEah3k/2P
Is9mLqEnInXeMRFmrMaePhq2zWc6QmhSfXgLI2ew/8WQVl75GIBJdVhT7JzYencr0c3KezDcYw/p
A3YWLyCUklKVQ5oLz4EqJP/nG3+mxSd7YxF5e6m9wyTQqc/+dd/8Nfkfyg48aIsmMb5t3pF5IkI8
Fh8JaF+UTG5e6OJCOMft9q6pXLYi35BXySLgB4bWydDulpNKvlBs9q4Y0+ajMkrX1VytRbBUvdQR
VHWPtE7hDRbO3C0F1RZ2nnS7hPJMFwz56tLbZpB+M8A2TE2r9MO/gRrktr2FBIFR1OgVRPxMtpMZ
wjQG1fehlm2LqAJt0qtX2wOCfGnpflPU228henXeQq+GEtadoP+4dKpe4eVmMH5WtJIn+2YCikBw
XVgl2mXJJMuvqcS0aGHtlapbhv+JjcoyMKivWGzH+xZLSv+BKmBpwYOaAnwN08aZfJNphNIGfN6o
jP0+Ou3HefWn2rKpWelC1iGDyA95TUIDfTfdgY9SzXoiJOlFdg5MfGoxaJFugXebJDA0PCUmWU2Y
rk6+HIKU5i4BOw+k5m+yH4LZaOSIoIzoBaNq1hiSZRzn1fIdTALyiuBW/BXFTqG9AYeocIvvV56F
D/Joh4DUm5wEX+OivtpN0EzOhYRNsW/BEPzTrZWcn/hLMA5wRkrU5trVGd2DSMPtCfeYPMIyHTm+
BOKxHX4mKNizMVgY/MWisbIffKtjRYgZk92VRdqaarwQlJxyD57/X5XRgT00I7w5y4/eIYvmi3SG
Nd4/e0SexjB9Rk9l8cvNWnrf2fLG4ug7mZOqgRld76eq8TxbIdWvlIM1TNSE9NKo74TRWZ9KwjD3
D0MOkb/E8RJDyohqqcFw2DQdo3dxJH+9RO64b5danB680c0XfiZtfpxaklm9i9grAO00tr9M189k
mT1fiee1fI+oWp0JeHciWALhV9iRM+Z7nZP9TVKRIW/Q0/Gksf6ZUB3UC/Bs8XTcQJGL5SleKe8w
lfE9EeFNU0rkOVgi9P+W6uXdNfx5pxXM2B0FuW8BnwPsVIzS54wgDhIAtuKKCf+l6rfqZPs8yNrO
3h3XFqTc2BQS1AX0ogSW6Je4BeNb3SrkWOFpAVIdg5USx+k3lf7fGdpaUaA/E6oBHXLUFbhkqPur
AkxL8lacevi9dGHp/iV7UeIdwRUN1hUpVSEic0JSalfbnOBvKVbYSBHfrtZQMhxLjEnpj9sTxmzL
FqyO9cXJMMUxNtESGoBiAbYPgfsttExiVtALAzUUUm7Ai2G6wMwDSuUUBoql3Cn69TRTWglVP63b
0ScgZa5IAhb9eFzOwUguqQHfRKEJEykg56WjmBirWGadPSfRb+MLg4MDmlTw5FNbaNhDqZNyvRIQ
KrXjcxXbzGZOo4XXSoyoupGD3Bh+A0IVlBm09fMDmlg2VeBVBEuqySC2z7Xc5WEfMkNhICLWmPx4
XkBgSmbmc9jSJascBuPvkoCQ9CCnm4olQmej3WAwM5YKClYGYsdtgi+lwaV6wK3k6ViA28ZBKLVu
KGDqBXr/thBdFg0ikVw66Y4VbAGigqU3F+t+NBvYgpCS+7VUcrxE7rZM6HyDcyd+o+bB9hF78KwU
TNk3kLyWuTrhZ6ShA3+u/FD2uAZPebCdp9s9Rinn4y2DRcR7v7qvsD2wy9wCJapw5c6M408Z1A2O
nG7Tgo1glvLwrckS/devAJ+9Y0viSrNN7GoM0td0yFeKAYcw55foVHxzOcr801/1ChLKfOl25LPk
CpQy9wHJaiAYXsVdlXxA0QzrFHSSgqwT8nk22PiGWbKH4zXBPbIxJD5lfA1w7BNvZ1xcxSWSpg0K
CLhQwJSeZCrXnaDiSntkrzN9ZlcgT+bddPFS83X2rMHJQ7oT6E+ZWsV+AVD2U8lccSMwR4AM+Jbo
wIWxbk5SuGgeI74UdYy/DHJY2j2GUYPeoEtRfyWInRtT60MpTYAUGLe2W99vH6urG/f0+7nAkJfH
DgDtoTrHBJnHWSz2H11Rpnhp65HmMBF7CQt61QblUYMvb3oyEgby+bh78Fqc1szzABhO29UOG8e7
JV4F1UUB9xsxhKGVj5fTcRh/NhnbMsu2QqA/PNbs9+/Yctz4WQNv0mnaeHp7nZmZRcBWlzzdJSYS
5nR03yPKGq+MpY+uYUlBRjiso5kBWK3YPvtU8/uM42zcUHOVHpqX0lSg0W6hjOPWj5+VKSGpa0I4
uZ4DVURvUeCgf5eQ9YW42fi2hciw6qetuI4cdWH4MCaq3+SsSMULygD20tKG5e0nPmyLHPwT2PAU
Hs14XmTvJaqzOnPqrk4LsL4oJmPcj7v6owqfldvGLXygGp8ThON8HcNXCpQg9EaLQj0QiV1U6Rsu
afDH2uWBCI7abMjD5P6X4J8srde0hAGO4h3E4yyZuUXjaJsMmMRpb23DJIX/kDPq67updjwAChnz
rvT1WpvqKCaAu2C9odPyNDzuhbfFyYZEGboJsRBhJgplPmG1ulZqa+jfdbxPiBdGVKlH1vDjYbXY
OiPoZFnli2pGxzu0M4MdH+zVsR7p3Cr/RIv+PLyydbYisQd60T1UpsXKkQvH8gBZQ+1DsnCB6BGl
cAekh9SU/R1ZdEKMDRTpHYO3KqsgIrSNANQyl4lZemtlxGoQjN1DWgqAVYphuGydm/EpfmNfDL+p
e05kmdC7uZAtGKn3O+qRcfqaK2PbG7XUgjQDNy9Q++puyS9RNbbJr4RdJdMVNaZbRQdhxGF4g7YP
Gd3tGbRtsxZmCt0IXutNeE3sMG1qmOW5QzUdPXHzwydSdIdG2bs4O2vfPli9PzXFT0GEnfBmAzcf
1VajHpZqnvQvw6BN+4sYKem7HfUm2Bk1ks7UrY6NqLpSkahE49jRQqEZ1+Hs/YfaJA8zq9g5ap/i
j/B0U1nCz2Sv+USGpD8QjGTgTQICEwL+HaZNVq7QX2BVHqhBJLflZjEwmCSqBrHApO4iSKNQNaay
cQxT0LI8pY/in+QBNik6GwlBAIeKRdtPYBNfjyo7TgVfuOHFDFLHgD88c1a3w65pStLSBOb+gwmv
AQkk010p1qzdFrwAtATseWEpR7NE9d5NgCK76Zhl7VVhJUAVoM9P6+OxqJxI0XA+wpgkkZWZEpV5
hCD9ODnO7kFkeqDnfSUkXu6ZSt3haOyhYLSrXZ8T3xqeTITu4fUauk0qq5AKp6cVTV/NualjPgwY
kP/lIC+bZjfLC+teJovXzqLem1RJnmZNKooB1KMIB0zqXO7g35cM1o3W/r/FdOrSXjDJsm/FdRQU
UEwrDkCqex7yO0vRWxjtmlKlH0wOTNHlXXfJnSiOv38ZSx4lbc+WH4NMckpDx2dZIqb8HBWAaQYp
FAY0TJO7l3QcT57cpCFPzlgIjQYiyCJlPXdZAdmlsPaqZ7p2v/MURs48hxNM5x5AY73BQaVJoAKz
zxZ5PTrzjqWcBu6V8MR1vaER3SqJI9Tb3d1D5jh/JDV3dTveuorKZod+yk7O8rxaMoqkhJNtVv1y
t1jdWuRnw77FzkP58MhhA75Z6XadihK2nNAXjfNV6PlIHIxXS6XQ6VW4C6EdqsBL2EfUlJv4gedu
GHbEtkjoyqfOT+zCq63N+bUdZ3uJX3GrUbvgFWeO2h82re4+7/njJ0BT9jLgh9bbBp2qBliSRn31
QH4Nu4JUcrdXWxKfsN7P2dE8sU5fTYYb3dhld3DtSA86RPWVLipf7w590X4i4TCfSNcYNlhfzSzy
ONh+NuqnAMQQRyrgeYSj54yOuGNqEvuGtKNxrBcwpZUOTNY7xms6RTGJQDeyBD3iJS4eR8MDDNhQ
65oFUNiu67wUDrDisoSw0+QLklBCNHHj456c4GBdBAZB9JkJWjpb57NFb7u0MQ+oeHrBk0ywjW5D
HsNURFJXulqYpPnIhmw0YTAum6Au+LHpMXwgMnNNqRB/ujDzINl+N/WGSxmGxVvgMjxVaAYsX14/
EoglS5k682fUbYvZhN8D8F/PhRRwDKgWXed3mTakll0+rPvTpTOXYWdaL5Oj3NP2SfRkqxGe2x8f
j0Kp5sk5CfYxQnIa+ME2jHvxlwv5ffbKSJ9r/fEW44nHspkm03Kz2HtOZY+oIydaIJB8XP1Hekno
kEEM5xEWpMjqCG31L69oQrgUsvHWIJ7h+kkSRueCGZ8QjZyv4eYQ3R5caSgWARouJ4/ovHDJZ9oW
BOyKKrMXFovsnslGH9bZIjG3W2/SGJRMVeurggFUcnQNFweklRYT8yQomCCqZaeUNM1oIqgBE/cn
m0xVL9Q4f/PhJ+MMYw4hbQxzUxqha83daKG9SER8Xd+6ETwK+2EGcHaRk7axbfR/o7DzirPb1ddM
fTVKsbPEoE6Iyo9SM4TrgOJ/TGmdlDmPB6LP+ADo7wxnbv5hqGFVKcLoVySFoe9DXA2MPQuy1Yiu
D0jyATZnh9vKhQXXfZ8k5/4N5GGFn7QdXYX/dfulH85sAi8EVsaD158Q5hiIcAfjX5Qi4I194RsQ
E4lgR3WlN0ALVwrNqMsq+81t3cIHjcrWC3jLuj+QCmubwQ2g4yVf3jCARI7O6SPdCJCTe3L/2Oj7
A6tP/p5gOABFFJC52wBA9+eTUBHRRh8bGBq5SLD1GneYaFiGwvd4E+RdQT3zxVnv0SprwTaYDSM5
2iDs/imXH3uInIAavY4L7zI+zyb5wOqi6P7MDN33cjba4Xkd/PpmsQhDTPoERyFcWkRm65UJ2BSo
A/voyqwTukWhSqVxw3iD5JEA+NcCgpJVpu1ThUXylr5vkfWbrHag54InsTRLbuXRo9XeSEVMk8KR
dGR4WfBHwvRmN+6KD92JLUuL8N9JFg8qUpqJ9v5EIA3Usaf1xd6qYqnU2jMaA/knvqsTdCH8Hfxx
6iv2MCrSAQAKgb054T5z8FFFq5J5dqmzEIK6eZDb3BIxGEBwndXqLHB3gmSGYiG1SkpC3ieldPh6
bgSHLTwzVt0SEQOwJyFhS8B7negkDGBtV0fg3k3Ao32ENMEEBUODbIW48arLJkVuxwBr4TzjQLeu
+rb+ZZ+Uf7aT8tjKDY24fa8hcfUqEHX+V/otFs8qIn8djI7Z5yrw0rdrYmPCZ2EgGlJx/hwdDCNn
Ox1HMffNd63fyXzVt8pltVKLleF7bgyObCnpBc3DjBChSW9n/vOy3zXhC6r71Ths/elzyx3wMc0L
rSZxjFjAKCgZX70xQ+VYqGJk1YLep/ZTPuJXa2KKvyr17j/Cj6Ac1xcPO3ABScuPsnFLM3s4XyDO
uyfMSkjFD6jzdiNlNDeQxoQ2pJVI9RYlXmGeSdIXadVVHj2EamY4PqfGfb4AiD4wZE10ExXwdGSW
DhuNC2R/QxoiTo61DuFqE2DALTV7QLgTdGXGJUg7IG479rUGBBPrNbBDIuZA+5hGMoI67V5iJb2z
nURExVAqpN9H55Y7geEKBDS1a/33ne00ENZ3exUiXctfyvS59SFVEjDqmeXnFDV/aVlgquvodhLv
PifkGlNusx1Ks9dDRK9HbKcmxzoLL8NLfPx6xa5roq+enyCa4KdZhxJ823lBPTC56nG/8unhKqjM
hwUDQWYhjLJCBHDAIQzkvno+YUCp2lvYsT1gv0h/pSSZjV8H9uCI8jH87zX71jzDHoOVEZz6qGgn
zFmn9K4NMkGYhNsk7LOgGrPKdJUQ8OEThrg9dLnVnuPATto0DlwzcJs5U3EfgN8cusjT2ToKxu+3
mH816mRF94sNf7O3Vc4guk8vXgJt6ap2JWKTLL7+bKLW+BWQUxRGNiughM7cSTG/xhbdekCyV/J6
aS4lvDZXOaLJcRbzCKW4omWHPMQrKVwvZMHmLw8juXJdCz2OtlDXRuQT1wBE0ezj5d5DqMIXgG1Y
WCEHRFlfDrSdIj9aHi0ih8hsPsTVFQsaYGu70URAc+XCfTKs2Jzu9YSEOV3mBaGRBO6eGESAQTKJ
M1TVHxwUEi++rIujzZjsZX41A/BFNrdGm+CnJlSgG0PCbOrVszpLtGub+5if2OHPVlmRk5tdAZ54
58tD/k0JK3ou0LBbKWLqxBu8jYy50ApzdY8BVCEjguogd/+46QqZwSk5bluXS8G6THFeJN5nP5C1
vP0S1SRKLnIrU41FyHLsCXZkzElFGsrDkCsiCXJXNm+bwRzePZiRZRQz2PRyxMQcgjVPweSCFFd4
83BrOjdOvo/YrqLiimPNZBx+Cs+E6fr8fSGu1WMrPNKO6SwmspG6VrqfHIPqCROU0ywfAgiBPx6U
v0amc45d/Eq3OsCO/Qr9QFmjlV5pKEJLPk/9S7BpvCSukglWOzW6U2oELXMkqjbbZoHRtPoMBK8B
WDkwIoYpxLj79GV/Dj8TIwa2L9yEEcE6XvbdCXNZ8Shj8yPUHvR+INvZ7sWXS497sMoJlzOVftEX
yAM7dXpUAcJWZ8jXQiXLDd8AF9Gu/hPhU6Y88mw7Fumosf9iCTTJQlJwRZhiyGKHltDitiwO3axt
hL1HEmxscAiMaDCugCUC3UorqUim5mWYYy7L2KfhE/sxjQpEu3v4yxsQYg8DYCkAratYffp1Wef9
ypVo/eQ/Sz3FHuOkTor15ojLq8ulwpoIxc15/Kz+1+ckBiX8k832YYy9EV6llipAWsnwf6AjQE2L
sBh3IVtoHEHZID8ldiQu6AdFS3uwWNmqnMco6JGcLsmfXrPpNpbfsPx/a3q/6cB/fOu28M55ySt4
iv0MDQqlLz7IAzNRA9jkkIPkDD3nw9VvK/wdHnj440+cOoWxfiYJzDa5KZO8XtynDcDYm1CdymPj
MuwjBSM65dpTqOjLhhpexXW+p5OV/GvuSh1cACxOkYm77y5tjOANKXrI4yCRgTzuyTHCnm/C6dWY
sY56fXRaZLJHYEzkqJs5wUwAPQdq3V6Wb083xy76ESvNISnC1rcgt7C6GYNEQiLXQoZ7y87WXfzP
P9YSKhSuu9Zfn8dULQOQEYFtlV1Z+JlqJN4daNoML3Rqp92ZsEEdU++Phdx+EiFi4k5o1cTGLeh2
C3dzP6QQlXn25zucQNs48mqP+crb0ieOR8wMm0aLuRioGgOTdZHWFQQxJAhOJ0M7p1unnuYYueCY
ngSEBnu4CD6+wsafNL3cX9EP+JTueqE7rYB3OnhrTluW+8p61rL80UXCDj1fqrAGqwDMlH4AMOsb
eqglOtRe1p20TK5HTcxJ1NZLS+SNNpn6uuOfbEy19fMeh8sh5qCa66syRLL6y3fDmX8IvZuGN/hC
DN+/AYKQThAvVoFiX74C2bkPIyCGs5sMJ27HVAHGAWa8Tz6lHpiV/kCKq7LDAejpgJ9BLD4/oc/c
5/iFUF0RO8pb/q0gdOTvNoluOtM+4edI6Cn1kxOKn6Pce/XqXNs5Qx9pBBKxiVZXFalO0sjpw+LE
Kn6kjg/dlscmB2d64+sW/siwpzbAPVqsqmyEPws6m5ujCiOQerc8iQ5kvYCp1eFoxLnjSLRdBT7K
6M3jSQQsDBBN577Ck2eW/tpIvHttUB8V0pd0js8YA48PTzRVydV7u5+leq87sZClj04T5w2b1acY
8h0kEMGcppOPfbrYF0KJe9io6KsilkboNVPv9jKiZoriCH0blB1uYGfvx/Zr3fvrHeroqJK0YyGY
WbpQ83l23cbbOEOgKqkqi+HFugRdGa7innDGSQvNvYOmZXS5wg4Zfz7YpAIbbFxkdNXpp0qczsZy
WsIVTtdVsJUQpyh8gPzj3iK6ImuYL7F0DW64lEIa2J09NH/rLZfG7Pj+hHGjz24GAanFgDOILmxz
NqZA4yQG3Xq2Xw0DlfcsKgtSVJaUlVGt22xSB9FX14+Ps/d0WBqOdsW/hWKWSAI/TdLTc8MkALmK
HpBTuL5p5MAPBlMHM23H4Y7oJEbbpIfQZ2Si1PwQyfQFh75UB4fF87rNyCsLHI34qZeid41jzXqL
fw50nhpkhV9GzCIrbPFT1im8cddDgFaMibLwtgtAjHqWLnSOzpTT2lbh8wuSoKG2INLFM2IS0peT
73Ce8L9j8UbSvSg4tgSV2mDJlzY6cib8cjfV0dZZ4R4ictUbu+KTFIGHx3krgQ78oTW/Up354DZY
Zfg2tYt9JrQfW3UNqO+ezzskpyIEzQKsWJbKkCzd1+wS7Y4zR2YeV9iynRNrPbcj2n7q+1CRexLq
OXDrEbfvcmj9XD6pB+fA7JhcjD/crZV9qYLs5QXDpXdkRUjaZSuzeL0DohdctrOJJI49rX1TAWss
RTbDaPPw5Y8r5KorX4b0vjGYzAT7qhGd4nLFGG4XuE592gwPwk2wzmTGeiiNHMNJPWLyDlA/cZbq
5QXqrFMrW8pIl6SFrrmCYYN11zpl4/et0DxdvGLqLo+qPy8WPsEd6FNHqQSXNaV6SEBh0UhB9doL
L4+mbYU4UWdjBZdUpvnw3fS+fddSrL5TMHIdtrI5shPOy4gKR2B60wn5nplCQIjFhMakJuPVEZ/A
Cgy5z/Bgn+fZHPfDOPJxpEk7a74Ox/tJCnfyJ5q/ubzA0eKi9lLddaIg2Xo6kMjGVilhdp+OYVx/
NxI2fH21ZK3YPNuuqs2r2KLau9fSjnOrMrAmXmxkm/4djDlHByLvcZxvld5RSGoUcUCS6kJm9iVS
1QDe8hA95FHZAOkJTaLwKCZtl8j9dlbqykWuEyWGQl0Zg0a6NmETtyw9AnxFheebybGcPyBP/puv
9CDKcXfeZaf/6GaH/FmHwhZytbd4hWR+N6e57qBGQDaiWEHjMdRl0oBXU1VCmGodptX/mmSCJRtW
OzoM0QBsvUj1M2c0cplUG6nefYgBHdZXgQJQivifPVXJGsuM7rf7Ev95S3Y4uieDC7oQrFHrwsYM
liQfNSfWe3IgnWeFqgC9WwcxJQif2pQLBJdLO09LSkUzjnDs9t6QlBl8832Sjd9ckd2is3IoaZI3
UNo3RQ+bYI+Niv8Kk7COGARF53dADUzcQr3xvpugqYI1fx4cXBLY/4fW17N7g0gLV5s58SYQNNrk
aS6J1GZSUksLCgsS/HVhPLkXt5RWH+znWKDpHQDDfGp4HZotoqW7fXNJZ/NyOiGMJuFXht1lR9VU
bsmY3gptqNoXlVuPmoAuHbmg+4/nMzV6JFCa0Qh6BdpzMGi8JmTkXEnLbm7KecxhcrBRy9mWb8iE
oPb5mPhxHPgaoCg/l1R4gYgB4MNnDTDk0hBVj5yMCQcWusAkziKsYttLfg0YWbYRvmwPrBnHt9sw
QkPEiRVXrLieV4zW0i58Grl5jYbwPs6jCZSQqU6wxn9byIgJmzLIJ5sDmduhMgnm9VZW4v337O8w
3yrZi2HHOfqw/dAjYgS1BILRYVWoEy25xxMhHcl7y+BDh1Od6NQRjNZLzkaR4gabSV423HehFQ4G
gAlB35Lt+D+jylBvIk5bPMaobdktZUoXfiTvfkDLZU+wll6fdRYM3fxYdoQqZTApyxOPSp4DGnBT
eeAenqeWLo8gTQkkJmHspc9Wny2zsF0lQ06m34DxEecNYP5F+GnHDhd4n1z+YGQwIgC0Y8N1mEkf
ZrT6iFVNsvhnyZwsXue4FtRFLG9b9VlQDaDWUjl9R7GKPoDVEpU1a9aNmtVvo9n82lJPQerW9LF/
1VbH2ZicgpXj/EwT+U/ytxuI0pXoHQKOqysR5bMRN583dVWENzY9+MzQt6meVr0CUc4fu9+VNL5J
ZOzbG2bS+aC++k6M/ldfVXTQW9h/UrRDTuVj/TOgfk5W5JH3HiE0m7RBs7iBLcOdCDgKNb4zapyw
bzvjoHzbuwc9CuPgJnvmnGm1JmyoIEminbgVwAAFG91kvQNz2icUgpZ2kLW9/aUxzzR9OsBk39/s
52XP7q6xtXrFQS/NZChGdeicTWi3D7DgdqzUIGm2t0fUlq5mL2a9+7rwbJaehzPGviZGt0VZBq2b
/RvQlXwvH+WPtU+02+mi8s3WE+uK3RxzM09fXPYGqEp+ceVApv0jCSOhXgoSZinqzd9waSoxS9Hf
0ZZgG2neiwFeIHPFR7dU4fZbXqhCNa0as9GC1qdE6+ldjh72laf7YWWJY/ze3yy+MU3L/sN6myBq
bRuoUHLy5A3T6kkm+PxbD7FqCTUXlBlMx9EdwPajyRJ+Y3yo0Yklq1/v2mNctNc8I9ryR5bO4tVC
NgQNyrBZzdjlb1TifpfePZ5o7geG6PN07yWps7KqgMASDJw6hRbJTUZ6WwfuZhb9vqGxBs79LoJb
vvHpzR45UJCrq8AsEP5E5b5Nn7sEDkpNvd8zZ5tzGTZZ6TK3chF19LULdtiKfsgqI7xGyxRS+Ayk
qk8CXVxS2vdVpU5uXhKlNycjwfcGT7QscFUJ1Jg6xBHoWLef/oSP3wXAA1XshEsUxHumYDeRWWP+
fprzrdHCMxL14zrtCQ891Erdqjw9q8YdiknwBZwv1tu/vNfD5NTVATIQaXsq/lGS4TJtkxUwhzI1
RSSB3wD1ZmDv6dBf+OSyfUFYmftnIWyuVKwrEcCS9UIxncWkC0WTAPt0MIHCdhMl3PDNjqlr3l1P
goLCMvq6yicaAcCcJioQMaXXM0r9ufwTU2dTFT3nilzi1c6kb2zci675d1SyWLsaAhBrgvFwjI9o
KpwUnjg8YvtIvEtcsGtSnD+bcbWflkhgzXnOHB4mJ4F+pBpx5ZxrSypBfY6JLUF0wXQQ7gkyheNT
jxtbZmf3nW7e4UWL/4TjvKvxQltSQdkkkFIkLenEl/b2pMPQuj4uwZLAnazks0NJV16n5EgxM4jh
LJ6i4glIpKxbLEdTXbYmuSa8Ls2AfB9d+bPTPUVdbBDLxC9QwqsQRRsIdEtbDNLybZ28HsJd0NcA
HxdHt893gijTzqHBmExHpXAv4MQmpFLj0png33LuVfEezlfGetz4en+I1AQPI8H/SI1QbqN3BI7t
jt1UghicOmBlNn3xjrlDg6pEgiFwkTVmAgmetfS342j8o05Txscmb6PQkPz324sIKy/KAqcVOsOq
xRuwxkxDyobSr0L5WKVlQGaU3nRVYpF/SMa3BrdekPaNVYSD9DTW44HbBMRWnq0vBobJRnx0joUI
aGt4VvKrbFv8kC1ZzDoCqXicL45JGARNGaDH3vjF2oe2zm0RDS1y/u83xRhdUxPhY+YecbhXzHbe
toVxSr8JF4mQYQbY/Rl8j+9M7YesQBHo2KAv5obU0hCssxW2YQoxwMQvMJ+bkWurdtIAcALDz+ex
JNqNXzsDhsx0zN3fT9nkv9+e0CQc9f4Ac+WCPJBXttgnNl1yeIEbeKmL0crYAz/4jjbXT2MnRJCk
DOh9Yzj3jJEpBm7094L0h7fjoMtL3s3nydTH07GJ1Et9mUyakQF7TrT/JWyv9dYhDpHNOMgcRJtL
+lvTpHmel3754jygdeQtREBNPXkmoD7dNus3wl9F+XM0X0+fJ3RBcRtZkAHTaV9vr/6KpAULEeeA
EYdqpd+/xPLhtY24dyNF9NZ6Qw1MccAAtm7vF6nQtcqaIR1/ia49cRrnn2Kgyvb3plsT9Zj6Y5lc
y5IQ9wTBpGdPh4AlTALrnxDYwveU1FY5/4NfLDOOy/SOeWSUKmmHWCAq9rU0lxEVOc249bkoGDk5
ImcQtaMxbVNWLQfLrvJQjn3qzc8RH3B9fiKNf/SlltJgIj9/+seQ/a7CGAumvJ+UIzr1gAIpBZoB
0Mcey+JrJ955ifErvsuSkbcNvvs/43nRU2iTeGlW/SonztYMh/Sp/1pkazH1rdaGN8UOcpwr6lwS
rqMuWx2Cz3XxJYch1OqptoSxD2mAZYOO1yCex8hAqqH/0d+uzTeVzjduSucCLcxeSyc+yOb5ztDk
qwTkWOuX3xQ4Rt/dX+j8htrXsjU+7zdwVQmMP4NSKAa3JjjYZVnf3xdqAfOI+GU52+JW8dHrBnvy
eLpkFD87CtZbM1XjAGncjoypUG1ake86KWjecH3pbLaNFGm2pu+8G8zxtlL7vI8oYWqyZGlWxTrB
+l+brLGVNr3EMRt3YFsDRHyGyJ+aArVkUBh4FaNsqcGUaMKHx/NlO8Gc0mQod5NKTwbRR1bskka0
r97Xupru8aFVTFjV9mRTb8TM6oacez+OYwALwSdBwBmzj6cc0l/8x7RjHJUjP0jpPWM/Swa+vSV+
7cHB0aed/vhGlPZrLSrxiwlH8g9PLRAHylIuonzfsUqSQ0tu4XfeQNoAsA/Qicq2QRIfcia7pf1D
j+kfDJ6UpeJEqujHyKAsr2b95MpuROHXuTlG7NtbKO49HKW8iynjmkDq4hFaCjdY4sQTTWpSJqYk
4h5KZvXSoMzWKOJ6cA2s75gCIvwymwKQC8RaSd4e9hDsJkkudH9jZ8iPK+JmF9i0jsxQaTOheHb/
NI4eQ1B9OZBfG1E20ffTgyp+M1nm1hGqwg1R76l/762ShSkx2iy0q9w0WeZuYzjx5J7nvulIPXEb
886hlBL50b3+sjwu+UUp94u93egetEb46j2y5vXRTUOFNuFYyybkRqeKPTPBEYEFPy+7dePxArTr
A3ifVXWaQvd0boe7Fpf9jT7177WDuY7gWSwdvCcGuGznpOTxbTc7TEro/L49WrmzQvRyeqhnefp9
qYLUNUdN/P6m8XRsYv/XYOPiYQ/ULU7Tl4wxC6DS9cPzb3wY/NDX8zF1EdwJfyVuPPMxsPonSAnW
bh/i8O6CBMTQKWT5rEoEIE0ss8xSqt9OrzGtx7evnfLHszmCNNHOWmPhc+fFIxl3T28qN9OKiHhw
L0DldPdxGkEcEsmzLXPi0YSZIO83WUfjfJKhE85ppbHvpZyooCO5yZdW9Lgz4vevm53MkOFrSTH8
a/MX8wZQTMqBk2nO2sv26HEzdTHR3FRFWv/gCiDV+/FQcK8jsySt1fHLVYn4/cUYvtpLPbpjKLDA
sGdbSJ9jXuVDPGkDV+Qv+NUA0sj+5E9dsw2UDU8enxsiOosxeos+XskUtCx1LBsP+r2+K1IraQ3j
Niv1/nOa804gwkw1CT07FTeEhC5a0iEaURmsMLGw4jA2x/QwAnE5WeO1LR0rHOxwz8Ctg+wpkqtq
6wvxZABThSR9+onf/W3ial9Qz/rngu6pOyxzj0ITfaO9B+3vrnmqn3RF0ijS4eQuLbT1pzBQhqoT
CTO2O7sZ8GjA1yAMjFDEnq2SiEOf5puMGJHhNF086eWIpcw5Y9aDGmKWZtzyHh6uzJy/23Aia78T
3Xea+bczKqs1P8Dbv5Viie/mX260i7NuspWlCFsj2Lv7spQbGn0fgkvbotQHl93jRKvOgR95WTNF
BFR0pMYxVbZZM4rtilLQZzTuabTHyzOEF4oQzAEVZJ4r7z039yTmhoue1tzpRUptxR1ygWhzgOfn
u3R14GnWaga7zAn0f9a9SqsJCsoc/55lhRTAi+wIEqqDWQrqkHzVCsFOCcTSVQ6NuWlOMNuBc7ZL
oh6Lxulqnt9FgvqW4s9PPXcYYFG2s5/n5wg3HZns6y1MqbLAHlr4Hg6Gio4IL1e1tO8S3LtCqGjC
Tyfhcww77tD0Bi92gmKDRaqOqyVR7v1lxnNdGsbSKVETm3nWBJSjbsKC0CA19GMvIKFdUe+IMOh3
stp2AnHgPzbwC4DeGI9oCBQE3uDcml0OdypZJ1rv3LUAax9xAPSa+J3ed9qapTBDySaXkTWVa9sJ
nmkckzQAjpumpUKzr82e9cO6MFiwUOpInCk7FB9k4YJGrje2EfOV68DTEtLS56mT+dja99gSpIsB
2Ehs/mzEbmIgFGv3vubhXtDR3jbhpmn+0rlFANcPcpRa401ndn5JLXwQ3BFGFCrMRWQGc1cvtyCA
dEQdP+rgGVVGKiH1FwgdWG2h5wrkCaGYfMGE/RibI471ge1Yt6tAvIZZYA1IVI5yJi97L7+ACiZ1
S0MvQfjhw8UbYIfw1iXUTuM9hanlJ17Cmbs8TW7dT6rbm6x5Pkf7nVfcQDcG35Gjjz3eWieT3yMA
cfoseAD3QvOojnYn1jJYlQa9vAlU8upghjbKZsPSNBDhuAgdr0ECCVFXLWV5qGWJszccOHOUt4Cr
2DA2xiSgD1VxDapLQbodgHtBr7xT3mgJfFjfBehoZnWeayDjGo9QPSvHpq4kNIdTMNRYJ1GnRsFF
cztqVt9zAJOJYBwjdKeByi1MVvImQxQc3FkO3WOt3LMC1h35EEs9du+X9fB1Zz/TH9a4TjR4da04
1cf+r1eVAp2OZtru8qiTqTn54qH7bdBXgnNPB1DqLL45Egn9K3/c1LtE+T3SxFk36JoWQOUw09EC
pgK/kNiVr1v1MopEWRblzOD2rMNMOnMrfy99V2FYNjesaV50Gx9GCDRbkshKGCwl1Ge/56+DGlgG
68FoxC4iEjBuonv3Sj0yCEHwvnD/78Bsd2doARBE/ymNA1KwGtzTR7BP2cxvisHX5BtQO7z3hU6j
Jf3Pq221efG/3Rg0gDYxfUAFba3b2vBo72Znp5zPGBcFsCE5uU1ei4RYA6dGu2Rbqon8n0A83nlh
eL6BIQJjsZ31C4TErQsHtIvI7Z/E/PnZpW1+zG4rORvIyLCBf11hSfYPI2TFg3XlEnIDgP+EhTYI
4A6r0a+7DwtqIE1xg6UDFmdijS4DkSSx/Dj3m8y551tcQjiXVQH2O695fut3TngBQIk++VGf/b6B
Of8PXqQjlAlfeLmAhbABDg5bMHPd51rxzPa+UnYva3piqLUhXp4nfiJUVuf5QFjs21WfU55uGQAQ
/1hvCtfUEYPhJ50v9Oskshnx8frqeUHaY0H3c7cpOqVqyvrtfUtPfsTn1uCJUrFC7jFSTFDN0hE2
iF8wx9/8DuwCmL99hif0P0Y5DKyYNoIUeSDhrunjn48YUNsyp4ixVJicAOWOpuDc6hUScBQI2qrK
aXhfNE6wHHIwCLx2JkXxrA5O64G9xsEh7Ecuio/w44hNGhddyMzJbcIMXCETGDpCQHm4L89NmCz3
5rlaRo6xbnb28crHRZhPJbwrtzU+ToCM8XEIlMMrYANN+MZHdMKlDbhQyNxBCB57zR2TpDsXt/hD
xpDdEsUOJraAzEgW5ir/Nbfc7guRygRdjAaS4CXKkf3H3xch7Ac5OcLCQuM8zaCsWDrRa+sVaoNg
kbCwS3lHqc+t/j4FPLfKvphmuYVGGWSRyVCPOga0deUUu2dmxXCIhXUGxuOIe9uwW3vYxRlv4lzq
mR09hDRROcAF/2pgQ6pFhq3T3ij73bvtJWfh3oBdT+teOqaCujD0Z9sItfQUh5iCICTWuMS+uplJ
zvA7XFH8C1170e5/Ux6wNA+ym+I9jSaAa6MpICr/mEUeq+Z/3TIUlZThXIXJgu4I+IWGPirrnGtm
2xm71mV/O/QNxLAg580KWtE9mFioBAHm7IVTrVtWTZq/AZOx+9cH0mEOHnq4cCKO/1HvMYebkl2N
ewXilXO4s/GT0leG5b2PVf0BP/OTCDmKdaM6OqDifHhG3IdwkQok0QKWXnS2Rwp9BTsi+L2a62rx
gpTdWHTEN1wUf4B2iUBhKHjb7OqErZHpt4172K+eiiEFYbL52/nA9W5hMs0zjKLwNtVt3vT/O45B
4OkV21lWZd+cfiQ4t3AKq1QtcVZj4loN5qKTty+4msMxeMo0Zp3b0BFwWxhNFKBLj6PPFKbhPkX5
dnj660/Xqrp640Ip2d6fCH8UdY4stT79B1N/c/N6+dVtYeLww5KtnHkZ3BXtmCGB5oi4A3p/N8vh
1wgD5DWoNgq7oFUMNvpuJOCwYB5Dq36YfdnrRl2Y0YTkrNde3cMl1dt1JcizJSIS3gHiFHFYv6CB
MxxP1m2gz1NwaGPo9DBfsn4jL2mwjlIxOsVY/m1jufpC0N2ds1a2p61co7XWA/rvvPzwsx+SAk8x
i73+eKB0IND4+WClOuf+QqLWYIo+gVvXaBcpRxe5S/ezgBZxfIpMs+YLIRr4iCe38f3yeOkriPeg
Ad6d1FwAupdEuvyg1DXDzhRX91bYrT6y886STgpsnRqcVuFs1lMGy0Il6dV8cz4pgRTF9yieXXaU
LXVa1vfkdrEa0dtjxZ6uQ99e/CduQdROI3nqqyVuLPGViBnhyVeV02Mo0qDYs3VCE+ywJ3pQn1A9
Mnq+vVY+NGp14PTndCZjdwaX3wW+5iTvd0Rc+fsd3b66oklecOlQY/qMt11/mNZEzYfH/Y5coDY1
EHLNwfeVF05CxzMlwSkBnTAIXnYpGXdd79NTdrmdJajFQlCmrF6+dR19UgHL4+pY+RwWImigQB8S
r3grIkHyV1f8hTgdAtU/q2YwmZvBA+0AyLKQHaCvOyQVgha0t24eOxQJYd2SXrW97xKYw6NXjHr+
ySkOYMujIzb38wM+5q68Z5mpQtTargdGbE6F8xcDlga7NyEAW0s+vVstaViKcRayINklKNm6EKPp
yJFLWCntulzRA8T019EgPBmrKg03Ks1duFSB5xacEJYZNQnSoTZIqXQsGYoGnFcl8Dc1k4QA2Ohz
Fin0vaDPuQ/n59rocqOE67PM7AdA3vxi4o9k5jJjJHDOtTEk0K6CTmoNfGSECjVNgIREZY+qBK8W
Z1UpGTH9BptSAtPnjPr2VYKvDAvh4Mi9ZFoCLQP+/5iAZbxzIdIoRWtW1IrB2xbjGjhsvH30jxaX
iC8gMecPrY+0p9wQ8zMNEyIxNmMXQXXmltdeRJ402N39Ul5HXeg2cFceOx9ygIyXiuRQ61qXg2ot
v7TZS4s6t1/0jiSlwObWFqc4DE509cxXHTBAupU9L044CTa+axzB4B4ncOKfz3j6tX2Xo9m+y5Vp
7Ac5kT6jADjSklzMja6ZNvHaP5V9kyy6OKFA9Tmp+036hXLnb2dekpkkl/rEs/miDkbmmBSW+JlN
8NjWnLALJfRdtq6tcKSqJjcwv2hwjY9Wncp5DVk4tvtrqL9Cvk8I13LRv7CxqmGqG/8fSaNgw2IU
38ciF3TTMUR7cf0GPzYvH/yv0exDaKlkR7XpX5W6e1NYH/++Dy75NKSvXUlBAP812NY0fG+q+q+H
joVw4C3/bQRro+EJ+S8wTo8/mQSw14idliTdM94kzMbvgvwg0j6Ow6Bn/Er95WKCji5144Ebigwy
I27cJxNjV8+62cp2jl4NNjoU7bQGEgNf3tjPl3kR4tLRgC7KdJlQD3Ot49qKOLZOCU+Zie/UhSsi
Xo0nNgIBTGU8Nq2M7tGpeV3zXOL+olIMK+CV0SAIR9C/UC8Qb8HQiAK544quk81glkVSHq7IPR5Q
9i0CYUfV4EPmJUgJKP2PkWv2Q6V6QIrS2P/Aso3N/zBD8K8C1zXOOvVn5yDOToEKbCzmQmzBXPJt
vbrHaOjYiM+TFRIBgWnJXPUBaMO9K+yAjjPSVsZ442ztn2o0OtrzwXU2RIuSzJHeL1Vp57JqHVSQ
GdTFLaVED8kS4Og/2xDjhIBEdwgu6HBj/28liLJPeUHDXN4ZBMfEIsjrEg9pDuTH+53loPUVQbkY
wjShQ2oz6gkygiocMquxjGfV0l9b/trldPJlmhjjXNvuJuabCRNf4jO/lD9oaGknfe+LW7QqEuiv
sMfOuuAsVRh2pkf+bZnO8Pl7mTnlj1ib43ULSEQJcjrLKBB41ukAr/TB1urPL9Wj/qT699zgQt5r
zZ7o0rzwjL8bYH3CiSkuIlQaYTcQbp2vTiS37QQ0hLtCzYXfwBhvfUKP/HLjQiKGYjsJjkLnjF3g
N65milzj5Xsu/+zbEx+07HzCv99cD6EMVR4/UyyWQege3nL5MV+7VJuXa+K6/TCz7kxMBnhZlsCb
4N5WQzNs03gJtTHEqDVKOJ+OoMs1Xv7npgQwNZ6KX1Bc9ta4wEL2SH9E47LpiCDQ2HBFF6nCi7c8
ntlssOaksoGZ5XAlY2T93RqWgJRr6b9snIAzwvckiKRJAr7hGIwp1MLjSivZVQ//hbYFf+P1AfSF
FVAUU6ZRPNRB5dJVAFTtaaGpOiMcH+kvJ7eYaYQ5Sbx9qFtp3VA3GfCwyNoxHMRRYlRCNzZLyLlb
t4i32ujGXEr253n9l0Q8LWIuQDhvk3GQfRLqOjW8JQswk36LmhIK15e1avcHmspJoVFY3HwGYzM2
xdJC+QXRPnphvB2onF7SzAwS47OC1cZru5XoXArxz1JHukDTeFQwf8FS9qp51XV3BWqBsMqrA2a7
uMaVSNMRw1ParQfg5xDr4Nvc3RYSjF+LVsdczHayImJuFp3X7DkZcziQsATVDXU2zw8c+xhIiPhg
eVkgFQoseS2p3J0R1crCY0atE5utzHXg2Dr5laO3Z8cQ1ph5JPsgqKsBXu2dDc8/h+m3CAiy7sfb
76U9eLKFmqUTU72BV7civDXWo4YBInnGXfPteeg7bZ2JSHdc6jmY1SR1m/f7VY6RsEvnVzDKdukv
v/g5nkddsm8hCo1yGbNlhxIE4fmMY3GRK/wfboNUt3rf0yGCxH2lIap1HTqu2D3nLd8M+ZbhJ1Na
YCMEcpSzbbFEIdPo8WynyPO5U1M1Gz2tStlzkJj95XuQxZwz/rDgFWKTnfHwOV+V0fRhEfM7XNgy
HuiOebs99fH6RHTRgg4UDiETSe+7WEP79rvfD/HVC0eciZWRhLqR/XXf8bGElRM4Ydjaw1jgZr8u
91zl6p0KjdnPSLizdWYbQoO7dFnonqcF+INtRy8HSHQyJtaXgsxxPVWnB/XGs4FjpoIU4C/URSvs
ycFK9yJspFizMP/y39tS4fvwsRaxOggBit8F6qEcSKbnyb4oABgiPgFggFZFsuqyG5bUdl906PyY
bfK1SuL4H4yjxwFhGr5O0hhdul2UHoOauqrra6yCIxTg/0qU7Tq3nOQzq9GyqIxYU2pLh1O/jO8K
dyJA/KJbPgjFwG1TRn7A9zTLvr9iQZmffkH4dIi9sofouU5Z2N0CSSdY9R1To3THHVIzEFSMtVfZ
c3BPNQPCF3vwUgVrhpaA+rg8P0I+sldEl9BjkuhwlMVUiVmsnwmWBa+8q+zMBCYd2XoFhpfoFVfg
ib44C+W32m9ypGy6s4njcThT/73mKpKtjD+R9JAu9g7zQ1W+l1WdceeYGgVMvM7a3gzrBeOb9uUF
Lu2cM2vDUNJnbaQlN+EqAiWJ6FbzqyAYbrRbBVm/YQ9ANcLMzKGOqONiyJ94ldJGID2/37Uzu1Ik
/TKldYSABPb1o8cWbVM4ew0Z+Dt5XsJn1IF6cpbsSyYFJ1qeeUkaCCtX1bg19UcPjDZONiKmxoqn
L/rL/UBAnvVDez+SxUrI+rV+umZ53VGTHt5THoKErYHams3dt2Zjk8ysLobVdwOaw1cw+AVWkVCe
VqXIAtDYMcAtdshBX3WBtDJ1sW0gj4g+H+O+RCqCmyC1U8VX7Qy/4QTDz5ZlNqA5ar71ixLFo/7v
hOwSpuEi4lHRGjMekzE0HTt9VRM2DUANXFIQ75vB+mHzTbeUcRksei/EUnwMPyLe6iCYhYWsttoZ
COGHNZ/a9YUWM7T2T7ERzPCKh2itkJU2Bz5FyCFbChHELcMfP+PfwMn8qsKfP7/mIuwUJkMentij
Ndlk0DjrRo+lagk6054DbooqU0J0WEMdYm1vrKcTZY4YOQJNpXgIs4gwMOSF3Lk4IF+r6G0yIRos
RhZ7SjwFvAGqmJI9hnrpX3HbzGcOcT1ACoMlv2Jl5YISJ+55G1iw6feemjIQKM4B3Q9Qq4LDrJqy
irBXnkgrtrBaKfrykcishAarJhVfhDHY83LPtO4fLKvFOxf+FnKbKZ7J87tUBpXtqijjM49BCRYD
WsFeMTKbbNM2Gnr30NpAt/C6RbnIb2LBlFfYhKfitlskleEoc88C3j2XcG8HXXDG9CrjAw8NFS17
JJ/C73yZ71nA5tqYovv2Hgm87PZdICiuiNL4WB+HRxUwrhxDxA9Ztl7VzV5FkP7da37zrJ9wpQpX
yATfIE9wtgt4S9ObmD02dz8+ZD5Hs+IqgQC4B72v5EYOBwnDcWQD8JFX09/sRLew7Q0V7jiNlCt6
g6ik7/tEY2eP8ni2C/1/2EDrayiGvE++xig+umVL088f11sqIGvrodaYD5IcjKWvUbtusZZyHK6F
+Ir6NceD0xhesYfd6dJ3ae5YVd8GpbEAFsxcLNM5aRs+plX7H01Su4URF8a04sI6LKFGc+5gKwwF
basqxOHntRhJSb+skZ+sC924/uovIGMLGNz5Xgb2dJ24JD0GM0lig/1iGv+DHikMUd6oopbG72Ro
W4iSo870ZIrOWig6jDtW634K2yb03Kq+yIFBR52rY5+FhFrDsBKLiJISn5wmy+uyOyh07N3AxfZ4
s/bwWeEYt+23JCBZZVr6ayoSYrBsykVoEf0ywy2LD2gCzRmzldjfaeyC5P8iYZYUfvRm4paFHyOx
NnbcTogJIsDU6CrYe/v5uTEBi1548EoJo8uAw2OKfIF166hv94SkNRQ4z1m06SzJoonHX8DzuuhC
XhrYXVAaoOLJxo10SOYBR/x4pyk5jNvhda2hoOZiT4R1+NkihPSzW8vdsFLPEpHsrn/NR/qHTqNL
zgvl2tQvktefKRe8BmOuvZHh+ifmsr2AONhirP5r6AKA5SFOqyd1OznpF3gpGjvaHEbL5jGCbkxP
7NajbMKHt67VPGeA2aVVlr9AvWdrtG1WS3DEWau61ltxpcAMKutKErUEFvwYzqn0mSKXtIMF1hTk
Bt1bKCm4fP4/fYbdQwR6R7qvnJ/3ILmQztheY8JhspTJ34Rymlrxeseaifh8BYUUC0QL6b+GL6Ir
KpAqcJvv9G/4d/syZfluaJwzHm70eYizcMbCwj0X/dVE872RAPG0yZ0WlTdoMBE1y5QD9ULZ+mhD
eCr21vEoiBV1hj7P0QqdR83Pnnz/p1oUPgrgMx+AxN6fVO5wz5zxksoES/CjcOZjZyWLcISb5JNC
0xJccRWi3zE0O5Esf+P5hSuPnJOBAUxxZq26mQArpdXmV+yEO7BLWhhtvLNorEn5rlsg8TAffH0Z
fdLe3BvhGM2mT3RDQ1SGMnjAxoqBZBvNjldpgNs2bF9E9ss99PHrbe+66UBG0cO6mi2Bx8UIb6jf
B9bUGeAkSDgKzuhgJV7J11Fx3maFDKeeEnil5oVy35xQWdHq573CSjUyJSkgNB7vpO7Is/6FnOuF
VRKhzozRf5cyYo5ud5Bn+eX1riyi7uM1DKDoWFA8xVZQJzSKLO3veTe+qjnbPzXTBBlsP2CIA9ep
Gj4cMMwHwMbQk3hWrswKZClAdv4T3iM81R6oLd+yarlHjER2YgDr7xEPrt1tqT6fgWqR0tHr5kYk
zOPSDzhEhlwr6da2wGDVyK9epyMa/4XpaLu+jtK4tHPutcs256njOolDlk54I3cSscaLGy8JkO9Z
bz8/YPGo8EdY0DLEYLy0MebK0YjIqko0ghiVu4hiut6AGK+4ch9yGz+adt+RxV9gyn5VT3tVMgPR
3i6/Xw/NEL5cejjwCE6QkxYhgpEx3JcD3rDjCsgb3V4llCKbIKVluyc+EnVlvGVbB6hNAKJTlJJI
CDh3aSkJh9BrkxRiVMr3cjH0qzfCNVKTl1oZFk9+MwBYq0bLxUO6YSOKrGGv8mI9k6pSHtPMnkGI
6bL2yhOQFegKQ+5leIqb0fEXo13GXZL5wE3xprDL2T2MuzIGHQvFGlJKIxaezYN7BpNXddy67tOD
CQiypf8A7HWX0FHtaAmqEb0FXrdbyR0jneiJ9Kxgd7CyjU3eI199C8mtVXVwEdbanl9U0lwWnVyt
u1QQR++ZbwPh+fdDQG8ghKAMgUSvJNb1pQ5CVpeneGBmnTPIaZm8NA8ve58fc6B9XRMINm7s/EVl
SVD/dl6Lp7zPQQRXp5DC9+Cx1nVzkBjKW/yJunhL6Nox3CNZ6lpd9HrFl0YDOCuNUkVyg5e8mbLS
i9E2VdWqorukUOBgU3jr4IGH65r5mI3tFAfgPwuiQNfdO3Jw5hc3OfS3ZSO0y6ECx/uJvwOXPTCK
zJACdUseUR9DbGoH8PDLd6iq1/dELDY3QtOA74zFuS+6ytKdl2oKp0WZCYPHZcFb4d7/DOrW96jZ
2MYDdQ4Us3tC27Vrk++WzLSNw15XsODf3kZOuNWc1rH9se8NWZqyoQctUDuavNEDrlc2Y0hpYBw2
q36K8wiYMCZm/5H6Y5JGar6UcqhuPdFfFzTX296ChudWoRLJvxq8m9gy0WxXEDkX6ucEtXuC9XuW
7hOypKQu7Sf40MMBHprBtkkAccTLnjAJZ/PAwUaFKziJ7i4ywb0myxA8IHZIl+xDrPhTW5GnL0EY
O2lfNjIHk2ER+rF4ruaYjg03NqAfPGEgcDvN4iEEvKn9vGgCYpz7gMapiVivGWHeQLPF8+YLNfdN
TXzDe6leKsqxHnjnQDYcGtqymyQSF1yC6S/CCOLwrSy9EhscQUhQFHrwkSGY6GUhGw0FIHMNKRXM
1E93Gfr/j3s6ocNYN+bEZ1owlcAphXy5qRiOwCXKBy3XIGcrPbNyIhWSs/PkMnC3dtZM/rEEr6wr
W4zmZKYgQ7k/muLDuJP6et96Vqt3ix2D6cAjImVzpwYnbTb4pkd9Cw7ueuLeOVjLAVankai/v4Kw
ZoD58iQCY4RfH+UTFywWOVWwUt6qadQ5Z/TWn/VOOMVmeCoFPTGp1lsW6XeRRuedeT+imBpaWL2q
pO9y4xMwBUvNxc2Gp3lgZvqyP2qLeXNr9G3QjtjgdRwz19mVDXqTYBo1r4ygrh4BW14fuRptf1tA
aWe1YQaIi/vTVIzjYBUMsIizrjE2pivUTDUNM6EaZ52Q8+6F6ghy1neW4SiU/5XQ02ihyPa+VMF0
LttterKR7gcphhcBiY/Kpu21rXdcVFsXh+n2LXlh5dw6+FU/H3DrO4Z+0U1NFS0OSPSJPjiycnbp
Zmk39P86caYWGiXLjsVrT/6zzZLxTxkz3vYfkYne8sLMdTmsmOdo3X38DEwJU6llET3n+zgMPr/q
bTwYHnYjskiTYjmpjXVtlivrlet6yrLEZ6RC5cJuUaLNJz2gvOr5iPzlS1vKk0kdKFYn57ZqImNy
vz4S2S1urCBmS/20pO8d5FVzu+nkpqH31oncpMlRKwrUOWuMf3/jMU9JcBmEvwybGWF4XRHN5NuU
8GUB/Qsx6kTg9iT2bV+y8jP9upmBu9wPyolmwKxXMqyL3iWSRIFmqtr5JL9UrefMZL21xcoeIO03
zAVdM8KO/t2pDPJceMrGlQIotZI892R6R/OOGcVLyCPl1nKT5CXwHl9ZV6ltLmCPtOKkNqj0ThG6
fqO82TjlUB9pkDGMZRM9xXwQQlmX2MsawSQlCU2Nq0+psKiDHpeweWBqChMbGynTPTwCEEaEuiHA
bhF9D5e0vDbQ7iXnZt1keeQ68ceeIniFRzG+lyJ65iYMpWH7Hw+ub0t2vPM+OtalOJfbg07ByD7+
CcFW1Ky1go6mNLiZ3DFqvMUTNi2pVCqJZRDU/BQ0+4jLDDH6fRLpLFkcq8vdACe3xwrmWXlD5shh
lnqbNhExHxIo3Gd9PY1ETKyps7Iq3qjD6aXgWJjUYUAC+zaeoCMaiYgwY8Gl5vOrlBp7hS9u+aC8
eM+qFgVXAyQuM1wiJOpnEElGPq7NGNki6ArYLHY67aKJowP3kwBlYjvwf50XETFw/dL2+303yZOs
6E3cJm+AR5wW9x2b0l498SDl3P6f0ENnySDekhX/BSbmKc+6FHUO9I9C892k9ifwF1ZuyfLhmhTV
g1rlLZ3ifgNuTsb72+DoaL9py+cmJRDeGna/GTWE880lUVhfL8vjKwrwE+vD2poA3dU1zhXc8k6a
f6bFkgLb6WCnjiyrGyrCyT8q9xwwUzfCsS+atZ5p1ra/oMjny6O/cT3p5nw/Geod5EY/ywgFELPc
Qz1WEoxBTGRwtypZM4fNXrdrmaBnyKx+2Z4vDhW8zJqM6F2+jw1vSUM92MWbfn0lH8gvi02TwUEe
hqvYAgHF64FB9gRn7SRAVGS5llUABWaeO4ZUVjh0EUvFjTKv3ijf0KgvTJfoWPnPf5WB3G5FhevD
4fl6VKOV2bzSf8h+LDjRETbOBAwCGw2v0VzWqXyy8picPBkmcdqSBAD5b+HfZYHcPIDHU60stxBA
OHJjPYVwA6qRcU2ohTW9WevyQAalRydwTbiaJX4osS0Z9LUDpx0bMCNiP9d8ofntVDHU3MP4Nqh2
zml+R3MFHQOBgakrPYsSAcCLP11wirmd2ZjT1HRd4RpOSAgMWbiViGVlf6/YD5tj88d5xLXwJh33
4sNI1HzYBSjBuDi8sjzHtiYYGIVj/nAYAr+gqRpePXDOeuzzJWokfQ+HZDhTGp3KoKP3OlhKb6cu
b+LddRMghgxJz8x5B0LsaLykmssS1DEeSympf9EF5TdC2LYye1TxHJLkKmJOQx6ax5IREW8ki5pC
C/O7PxVGLWtaHXVt1jY7PxPbOOYwZgg73sDXPLmjbJczFwotyPrMJ0whj21jl+Qfm18xxcNL7+RJ
m70saeLypww1bnlo2yHzTcsGyO5B+p35zOittS05bAsAb5fr/DNDPxQ9RwrMwTyj66nSN4nk8GSo
83k/Yxc+6TLFlxpZBTbzSq4mF7atCP8Y5PiREVdmdEoygj+W75koyafC0YiJntVUaloASAboTf0W
mJsgJt5m4qq/XYY7tjHSy4iJPYC952eqJpoRbtoyNVFSI8l3MTo43JmSDtLcbk+eoRR7mMMq7iCs
6KnVxWdn1fZUQ6X/C/fYButsGjnQxG2v/NsUZrabX50pUbkGmWibXv6+1XnCVfK3sSlthQWEbodB
pIaPcWESomfRs0pQaIR0BksemkNxaamZ5y7oOO7/ScyF29uD1v58MWh2mDsArJ+NgkdJGAoN+ixk
/7/nzDxTuJac2QoRRyq73QKy5hFEjsNjGZizXjqXI1Fpkv2pg8bJ4tjPb2hpNl7Pu3ghm82/wpVk
2vd4eIVIbUAJdMLjmpZFVSfMaYwGWjrAlXcB/tyKVdgwgU32Vtfd2Jp04ooFnBVZxd086ZHmILzH
JUego+PAK9BXmCJD2IRx7o557Tjwr2v4cPmpexoXz3egiy6V31fC4SGQBoN3B2hJ//U6Opgk26b5
p/52DeYME1st4UpSOWOGxZVCluHRp1dASQpddobIBzyq2zgGW+1UNFn9Q/POe6bs0Yqt07+u2QCd
Spp86VX41hSgitY75Hl6uv4YOm2ixi/ZS9cDOLfcUOF7PhI27rePRlIf36Wl2JsB+1JLJRs7fVEE
D8sTc/DUwB79Ejvt065PM4/gnAC8uHo2lEDm2uOtb4/el0q93UYKGIef9LhQMItRAw4GAUbKloNr
I8DtTBcJVpMrmgyRqtT6SOSozGJKlO9tQQ7HklrTh7vJOSj7BLl9rv/TRJokZGoIug6XbiV0+qiz
AFWCwGXT92gU/LicBXBXBfuyoGym+v40ZuO+yMjNqL3/iQvLUs6jYu/qJ+sz0Rsg+0uoqEZVoQig
6PcA6VI1iNDmd3LE+1qf9bxqW4BpSTn/W518sEBAVS+B/5XEPzZvrR3WXEEHRVcn79EDfMGuBDbW
n4QZFSGRfz21fBmiGPc3M+pt56iAM84yIgZgX4hPSQT84Zpv1tubQapUaRprUqEh1JN2WxKmeOpD
kKvcAXkpteFGHQvQEo/d4yF0udDBKaf/eYs15QlggcGrL5Jg5JMo9EJxH2hMUi5mKuyR6AbNYlce
Ndz8uMgKPfCj1mIdbzHmWShdR5SF0KW7SH/RGe9bUnUq0BcxKYyS98l+RjO80HI3nlMemmeTXZQG
JZWYWlyitCpe3xU622h/ValOxbsMBzrFAi7TuuyIewnQ4BDoJ2mRHGS6xkfrH279cHevKILVuCnZ
0WUQkx36mwLjWqOxTDrto3P9NlaizpxiOvZlb4b2y3WxVWAsDWvaGgR6eF+PpLMLb3mja4H8wKdI
JJelvhqSwcn2X/W3BzXxGzu920JY3NEhJvdYqyFwUQSaydWgdfITMAtnvry5680aucZyAauT0VR7
iCJSUded8xMqKliI1taYyLKJAok5dwyQrSmK0RbNmq9HN6BLWr5tC94ni9fG2nb1FvtpKdkQeP9O
abJHvdTma1+R44BjkdxSBF56E8zH92W7rgzTAJNv0LLBbMuvF52qjQGGBqJ4nTWuGIP2WWC0BDIF
GNagaqqaKHdKvAM5mkh36wQB8Da3W/A6ax4V/2IlwrVlSZ4gKc1yydnu7OL8PtuTBXqIvqv7epvq
zp6p/gJKHjOatz+2zt6Bny4R3tReNmMqjHeSRFe4dynGbzFPZ1CCr7WagOgnkp1jv/lKoyqAVcVM
Z2D8iN//0TD5q52G601CclHGjSE2x2TtDTnzbtq6pw7Q5oXSmsTLJeN3WHXCJGSARnXePiNI+0B/
WGCUbXMkeNxgTExQxC+lLG3Ssx8A1SknLIVhIiZ47OBekNVHA6608ajTGkkFs7VSZ9Mc5lofcoCY
v5LiXg7EiVDnU2EXJAhZlnp9S7lWif9Vfm9T8LE2O/6pw9+NmXk8X1081qLiCILOBhmH1stly+7E
fnB5CmuzOziWWcjs7Nbr+7h1sq7AJLedobyvaHNvN6DWif8gd/UD5nrAjREza51k5X4hwptnZsLo
ZCRYBmBkh5SUr9W59NZhzeSF2E8y9ELqUB1jwXPlYDRGdWY948Xc193wsaqKRQ6Wse6hnN9XkvRW
w0uj5SYjvkbBzZZqcl22jWw+uEQG1kb2Wu5WGHhSWxuGCyK2TTpknINuY0k7lHxddrkDQ/BmLzCI
m8MPMxST/MOkB/2mU4+gBvNlMnCDNuWSPk+tiKpwBt53FRVj1JVYiUE3oRo5B6kCMzdOCZuQHPSd
Gc+BWZWYjrHNdAOwaxgZptxrolzUum3dw/+/nAoh/Xcm/GsOEmBzQqWOCZUeMR6R0w+2pSaFOqJC
x0adabM+tywsDyQZkdaFtDlS1HPUqh631TKunpiCZkZVKrJuThXmEMwDQcwMrRUu8IgwNt1BDION
gDlaFEYksIKmbBWkFVgrc1ySzpQIB4DWcplhZhEJaeQmiEF+nvlcdOzYS5XTlxjyR9Nw4EDnIrCJ
mVFR14ye7GieOy2Bt9DAkFLwQS8qfLyE/b1Sy6ZKOdps3y6FeMK1TyNcNkMOIWUsl5TCDSGSgZEs
m1WL/ab1gsGywo0y6zen83Obi+QcOG5qYQ4jAuj+BibsQfvyrm1JaYVC8GwoKgAaiZS6WOMqhysa
9rwOqa7KUjMeq71ik3+wJk8UQ9dzhCt1kfmDC4UXRfKB7+YlIWrVpDyhxItIfH8Vmq0Gxv7Nj8XX
ACGg1EmbJWlDsSVLQg6rv+NfZ/Xzd2VTkfgfwBFLn0OrWZGHGmU5rpl6t09XxhvuDdrPHa24xIE/
bSV6T7tytLV0fqiDbXvVfH00f3zNMwr6V7zThVTmgZCtGo91MU9dUaZDEJiybELQOc0Bto7C5Qj+
kYiCl4rwpn1InMt+uyjEkwbs3Gkbw8igBwl7BDI82j2xjX0EZDgk/YsiRRMCwDxl8auJsZU9JU/h
h25aY9XfC01lOONAOPTHTjtpS1tD9ipr1w387XFvFabF0hjipn5zFfTTCcOiH1AamACvrYeVksVj
s+dMIqAc1+uOr6Wc7GPc3YZbj5cpwFBoPcl6hDjCIVl+O+znAH88P56flO3dOJbCShViPop7D54A
VOzgqvIzW5ptoApTJO4rKNwkWJtqNEiMwqQMLogbPTD79Nixh/28xyfZQahzRfzZbFyslyGa35RY
nChcRgI1c43Fly4nCA7eeDvNATCHIWXDZXHLrlYS0wz1LWNqz+uD35CnS3tY8LMZLcc3Oc6Mqq/p
e834WjYqmhTQEDd8e+hF+Jy+FdpXKKsr6DLkUfYvvKmalCRJHRU5mJzLjJ5V17nQXh6Y0246Qi7M
DqbABjt33zZWoP8jv6bm4udw2MD/GyXS+nQYzQfwFN2ZXftSwVwb7a5wSf+wu3SadfmcRQ5NFsf6
O7qsEP0sNHGgqmtj3m9RACeQbIBjOS0ylIS0mB9nOhWsnigA3vfQ71yVVkS5DApMXx/grE64lGpH
PT0Vbbe2LlufB4+hFYQcUT66/wwefmYnC5fH07v6NnH7jnpXapRBQh5uleujTTWSDG/cz2lka0Hx
XANDi+eyGzgXUH7EFedmTi5HyatjIC26oxBxwPe1KJ3jlKnbbJaySrcL25fZ0QKvXC7S7wD9oUu4
bscdqnzW1UGR3EoMoEsKuCDE4+Sl+XnxAHiT6GXnSkHnXHjXpR71I4rea585BjVrQRZLZCbNWM5C
2b0ih0aXbmaxevHUuIR7PXKlEqdJxTI6RJCxM0JtIHntC2L444VeFYi8nJlJPm5eSzkHYnaoFloh
3qWpVxvs0s43G9MoUqQBpJxYfEO8Yng9Ik9aQv9zjjK9CA+57XHER9UtICNlbY197/pmU5lEpcI+
4+IwX/M5Xvuu+Fi00jkKWHafEYaRY7FKMPODX/Sj7HxIrMkJgk7V1MUULGP3BnlR5JpIREbJdcsH
XIHhM/vob+KN3OAreJPYZigd46Bv5EJwjLNpJInkwR+AEM0FkPBr84htjkTERJNzVZYbNQgdtBn4
wrhYJtEkkZePgbvABO5WKfoyj5ibKnlKAx+beQJq4Efq1vFMUyXPuWHBAxl30L+9IDodBAULmQS/
0CEquiea9aj6iub9ZLQDyScXVyOrBdJbU7x0zQV3tixzqxTOEsyVJ46jZ9QrMIZ7TDyFbpSnyOES
fEYKbxj6bGE5/ycy5jxFukcqVEpnrmqnsh7+eZuMPGm3UejNj4P6OBcCzC8gYzLDWyvKT2/IKJos
GUQDmcH6bAtQOOZDisAyv2tW/8lthgdG4OfxcczXnHOgJs2DkX2FAA9twTH0ZvFwdaJRDwRv7tWQ
l3Eu9wy9tcRSbJGOOumWhr5IhQCek92O9gUj5jWEbQulDjyBRSelpcfOArcxeZ0mbtGxq+Fp2+Ea
q+Z0z2LHwpBHXih4JKprO5giuSsDt7H2iWImjHEswiEs933vQApzoiFbSIlyswjV/9zcrXlprKwu
s7ll1WMgrCSHCb9GZVLC5WSAyP76nYrxYMx1a4YtEuI2AkncvECDmZFMUVj3Xec6pN52rS8XQCM2
r0nPD3yw+l134f0I8Z6w38pDS+cyExEN59TeKkd7b1tWmldOd7lCRBdzTKmfZ77pe36X3cSnoY+p
1wzsnYh1YWJKWR+p3b41KZJ/8QBeVvgbkmwFfzblSr9C4QbNiBuJmiL5CGV2KFyjeJQfoD3vr7AU
AzjEJbx9FsUQQt2YteInODJaOmuf8wF0GFd/oSAokJcGurvwuBNIRZUFcQzyIVzEPjroHu/DiD06
SGkCCrVws4kLTty65pv0n9N2xC3STk8w+04+4BGhs4k+lr/Eh9H1kGF4RkdY0Hl6aTk/eDmhMUpW
4lXFJSRMQZlo+uunHOKGTFWQTkuP83t59KIS/49LwvybnxyyFd3KPJsKv7IqHnN6kCuKAVf/z80Z
2gwI7QbHa+HmJGNh2wrjM0wErMVUrJ3JK8KeTPAyxcNfs0eV3r+HyAUHq0URfKGpmJQFYIk/i3D9
4ZQ4OlqONfwQZYZiirToytnW3OiA5BQ6IykkQRQOmSfe/2gx1f4nMvRsIx21bD9FzOBMhJOdGZov
mxQtZTj4Lk3AHRKjcV6tgKJKHPfTfDXTBrr8fkUCCMIWdob/ww6Rz2wPSl+SICx1NVmESuFEhfx4
Qkw09Bzpjjs8TSTB/rXa34VjFUp4KbZWegFDwJYKPJnNoAZRqbwX1sE/NcS9QjqVyy6fdd9FG5OF
1y4M/1vipLOggsOqpjq3+M/oPYV2glN78wP69JEL3lazfijQitVcRq+q60MNnG5Hw4yl6cSZO/TZ
H5SKknVo/zpsUSQ/MXtR6v1/QwpMDmMICVGUM0EN+eetdfY9+7Eg0hcBCG+yYYM39AvLMzNJ67Cb
HYmtAbH6uJRcF/OCMjPg+UuFkAKCJdwkkbXHKpSDHcy65Z3Cls4JY54C7SeUC8d1G1DiHOxIGXOC
I+Rve98v/2kgcbw9EQ2N58inTJjWOYJtQPzvIGGQ6z4uqRmQJLi7/1hbdNjYM18B2FKK09RzcEo5
q0geutT607L0SA7Br/apmlGb1nBzWYgyCDGAMqdIT3/rtkaha16ZxXbzTAftRIxXcpV9wVhNMWlM
+d12n6iXar6CUJkBXO1q851ISTNqp7xrS8VZnCXtXt6KjTlz75hjuRN+jzgjHVPAbbp93aU14a9I
VNWR+hJccfz8KMuSVEjanoj8N+M0Cng+49nqZqvq3TO2eJhb4ypfgrVYyB368FjmaMnuSzEMdFie
Cb9GSVSZcLHnCxANFaP6w+Uy9Wrl7fTvA+6uFZaZtetskdtgzV6Uo6j+bCWQLpQmGU9FYBQPeWml
kcFTOoQo9ju5j++Jb0nI05aS2rfsIONA/5DkiqeJwSvOxtGQacVXEijeaXjF0tp5wPlHnjv43jwR
PA/gtAvGM1QsSE/77kj8KjZPLWuOCoHIvq94+PGtQyH8ahLlDfY7EoPMhnejZrjpqYsSDBKGtB0r
4PjklV9HLOVdvKNCcS3Ckm4+iv5VR9WQxZZZ9ZBeygbj56r///+X8c3NbPu3yOU8ioYknWb7fhyf
vxwMuQW1cYeI79KDzdORAMVM/wKFwOKQDcn/c0gxObUqA1noDTZppZiJV8ahm3URQq/r1EmBoThW
VJ3UzBdhH7rY5EkcSfg/DvUrrJZN16eJq0W777sYmLy34Q71pHot5vz28m7308+OV8+sYbD0EGw1
MC9zJ4JwLy8D/TpfWps/lZIdoNGx4nfGqSbdgOyl6RUDrI+Abw5Ff5IfHjX15cDhg/UDWLT8z4KE
RmZVGg1jh1k7bWQLCb0Zri1vuGZ8sErXkwjjMiDKF37Rog9cr9wluk0ScLFek+2UOpVwY9vXBMmP
+7hRFbyqHgXANibTbvrjyGq/CqcJ7FqP5BqRBCJgVKZzAvLRwstLOrWk1SnIpMd3K4P6x8x1vI1h
dPgWJC4nxyu5+k2PObSB9amHHcvTo0JEa9jMSjhNOBAg1v7l0DiCxCxJz0AzzQmDQES+9xNo+XXG
zmlr+mw2VGuj7/d3vyh3KV+Vqd7pkzsoP3j1HkBglJsmPsar2e64IWBlVXo76fb8U2dGiAfheHPl
xRz9gQ78ua4iqPcDWVUfD0vmz3hXCtoMaLgFXMLRcxiJqcc9ZyKhqfdRuMsGjZC6upa+1eVdMwwP
6yUcYyUZQgjticr3Vn9IBOOGvTrYmQwuHVHAT9BnPFshuOtW/I3mWDBNW8ALamX+TsTsXUgpwrpg
ELPx/Kw30F/6njfkQ70LXXjRT15XsS7q/ElEuy6bk6uI7qvC5SDchyMsK9UCUNiazgFCVMn5b+rV
IQW7LbnRKIC3vtL38YCLZqkaZs6xIbmNCd434Aw9dBswOGU4v8gbiubjCTVpYh4JvI18Jq5ZgsTT
d1ZmWuno/WQ/D2oRTb2cRU3qzeF9OTjhZ43DPMgRk+INA9UMfOF6J1cE3Qrf3bR6FoGYOsswtjaG
qBgLCjI6d1mHB/QjRnbaUrAjEFwsU1JgiKTkicNgek2hEuMpYr7qnIaMPddYc8epGjQ987ULNwWc
HQPNTm6Ih4fevthstzV56/e2VnWYvqcXsjTKydXvySo2GmAZt1Uf+zMQTRelS4EDBlBJ7OEwL7wV
aLc3SuVa9bXDDMMvRg2PZGUV9raboMqEhOxq1pgCaserBgfhcDc9kwpZEkvgmOacZY7G33MXfLJ2
dVmgjp0qKSU68+WIXXRecasMJYttn/XF8BevRi+Q1uyT1TIb3DCqUrPVH5m+t/m53NPXADO6iqEU
g6sai5rqeVGWWseqg+rdOqgWofTtCwjtbxpCh9rLOsSaifmtpyfyALZLUNKk8mbSzxbAM7OXL12S
9JggiegKUA6yp9aGqDH057MmBJ+vU0bzD/us2jCcD02m7qsJv9xYQrLWsth0qGMvubduw1NaBlri
H3zuHIJM/PEdhGhN27YWJ/iRDdLNmeZ+b2P4DhSGoBF0nuCnlVjm1GB22SWAQOCbhuq4PE+dk66T
1PoU3d4zAUhZPiQc4IG31ln2aWuVhIdt0lGRlia9IbcHN8aI7FRKm66JpjXPCNtmZFgQgE/p9AY9
ylIl6MQyLSeT0aQbISL+HESKzYSBXi56uxtbLJ+WftvOAELfXNsElit+hO/gVAIfVjhTqsDgrS7q
V6IpRIYtFI2x/kRg9+ufy/esbnBKuUn4sFZJif7Nm2IvEoEugh71bKDAd1g8+vjpo7vTqycTwSqJ
CIbcWOTohMG98Muukbg3nT93m55a1A3TusfB0iMYkq4gAEtWirRccmP/9bl9fFli4jqoTkBwYprR
L+oUtPYnBu22NQx6WAjiwJwW4qktNpuX1xVMS1zdACyXP9zyvfko5QYACB2oV8cR2ZPvwT5+um9B
Y2TLicv7BieLl3EAgnSSlT70sUb+e2TzdfE1/rIYmNwxnBNbkX6Gh8GEb5XNHbBS/4SImei90MlO
xYdoF+0aYXfKAIkKh103h5AG1md008x3tlNtQEoz1uBodQ6gzJqvTmrUX0zmyyhiIg4L2003Ar27
zDmzeJYh4JYehmsNYVzhG2wgxxMBJNiCDMCkH3m2xwQ9H85TVGYTL4THu0zN6Yn2kn42836OaqbV
GKv1YagDHpJ6KTrwjGNTIkN6QiKoS4pLGCPMfi9rm1Gkgk3HeOLDzzz+Hyf+sUW6S1rPcTBNSiup
DDdBql26fxOLJWCL1RTsruWdt8ulUu8QamgSTJu0EfB5Vzade7RAMu+isBsbLyj4j9toeavKSJqx
gPMPn8SvmyuBza/i0ZcnoofrlYiAACHT9c7Is5J3cQJAQly4nefn8IUJiO0njHlx4PfRse00MA8J
xOJoVl2sPHC4+NxIL/Wd/e4C2RDEDLlLyMv8FnK8c2ZsXtk3dtV5X9Ka8kTQGIhEiiXMFNFbNPLZ
vmL4tanvvDyE3aM1kuspskpusOF0MkmDLurXOOFUZWf7DSS8Dc+vDk2wQcZxCrA7FCp893G9Oimj
fgbHVXkesxqAZROhLYpy67kFPriE9blgFiv0+Bay8Nz+FFBsDrFmEqsAxAPv5zWfL3JmsD9WRcWX
f58zgaud8QY+NhNoHMcRdBAB6yRV6u94TfCbsaY7I5uRsqjjKxGWrcD8jGTmhwhNSs+Qs1gmhi2C
jDTGeKroTa5dUtj11tRJ8tyHUCoLIxZevA9PNsXVyRAKe9P3m8573mt7xHA8qRm+ySLfxbxoNkYW
NbcPZgqvH/Md4eZYx/lq3soBYqyMmZOC/lblznSHIomiZbc+EnkcUINyAnZlPZ2Zplqbx3p3dxPU
JE9IIf5fRYKOn4B39fvQ2Ud2n0nZ2qcrhUbfj27F31AB8X8pw/9Ta6YIkAzs2pdFvhZ/iiEoBbiS
bTRamy+nzLP0p3MAWc5e2y6ZRv66tE4hjPWeEX65bMLFQSz/SjgD+rkGcPi6xhiUBme0S8hrZA/J
SkQBRPs4JoxX+Sxsv1yy1g5qNNxU5GVtpS39GUTsBaLf8rhJisTQoa04eE0AzT2mL1fAobIzVwJ+
LvfjCim0NTiTmgQkP3YabAsPzyCVnOrfwA+D4tAQr4dHmiFkdYzXdtDPv2GxBnkd/baNXMLFm58a
Otu0OvP+SaRj+Gaa7elfUBG4crUZ8U6L/cTdZ9OrVGJ4z++tutQ5aVcfO4LiOQGiOjS/PMusv4aE
JHP2Q9wx3TScNElsWhYYz+cjgJ1pJyqfCoISVdlBfbdZWaAYPFuYKB4ok7Rm49TpGgsK1x7SxCao
BUBXrHYE0hxnDp5Aze4weYe69+c7j4BHFGtu0QXkSC/N1eAB6fIeDk2DMeb+lr+5v4S3d7QpbnNp
JaKxDGFQFKMLJLp5JT3bELmUc9vudW9SDK/S/8oGwP8JpCrlIS2ihwteaUQQ5o33fc8WwKJXA/Qg
cA0qpwGu3BYsikv0qc4NpqDlMgPicMc0epgqVGyecFe6VeXM+sJ2Z2X3vOxBPO2Mdm6EnEQ4Ua+D
n2PmGpmYnm5sSpFD3mYnTntg7nDSwjPiNKlgMIrta6Chitn+tMAG5j/tva9qaIJ9PRcI5Nqh86HW
yzyiZ+C0UE78Avbzw4gzpn/11av/QkOWgg9NSQHAWdCGQ3Bx0kcooHfpbg991vP/Wu2X8FQyCq0y
++rjh2WlX7+aEthGvpE2BCosSUaF2lNxBjJo/x/pJ5h8EWBZ7VAYEljJyjVCyp3BUV02koHTAsAC
flPTDMEUVb/hpQjezk4DA/aBbm/k6cQ2AFtItj4QALN+q4nzzABakE+klo511wXXq3RdykI/qpH5
G+GPYaznwhIzAQPpWT2SYNHDb9cG3PVqcLwwBB/HpBqwnZyhnp+c6YorXuOE/WzatD+Thd5ir/M1
u+e/W2JVYZeZTT45XN/ZBRFVeYS4oUo3VfDob6PZUGH8x3Jx+0cOf9A8R7tcSoQf9se46T/X7A8P
mfA1WJ8AjAyMYjl1TwV+L46TZG3xJMEd+ifPHlgUzqBisd0Cr5l4A/vzlc9RCf7C2hhiAEc4sjAO
uClDkwJnHUa79fAvrVaWzMtoSmRXHT8RNXr+yC5h3bpCJc4Fr+oT+PsM6qs8neFz+zbCGt0jQlfn
0ddpCWlCb78xZdhki6Pl44CY5yuub1NBGXE7fn2bd6V+CqVqE++55XYaKGbDvrvfS1b/VC0HjxY7
aXAN+45RWKMoYdm0f4uTZqdsHc+zizhUstxAGP2srnRWi2l7FfnjqhJqfGt8+cxQIrc9qO7Zrldb
7eVnmE5/pAAxlIYJojHrua8kZBH6kSe2tABRroTsso2n0adhmgI1mWLPJbJY2p47OeUO0GZ2IEe+
rjLM/eymVozkKL+x2kg364nszni2hr+nTH/UcY91+N288ulq8dvGd0ZRbC3h5NrJ1uKbYKFe3mdy
AzafuqOAAX6zBO8CqG/qt3avg9vyPifrOXWrHknLN/LvzcjjMR01Nyz0PNQdbhc+GnQOjpHvDXKs
KJYcnGNC9nHahWY4nsW1e6JfnlD/Oik9sOyqG3Ya/WJQ9e+AGe+82qazYzhHBvR/t7Yq67Z+Nn/m
r6z94lUm4rSiGK5l1za3A7wwycktM+sfMtUm0T7lQNzTEW+Ppumxx0IKKs9pITrM8FrovGdlmAdM
/9CVTqDckvzYvl5NV1jj2tSd7B4S85USnkaIXJOf8rucnMqMNeCCcud7ttHZSASg/FOdcdEFIdO1
kdG2OOT0sDfxl4Z3jSYNScCXqBbQJaMserGFKXwxcggd7NdTzO5mnkmXzrKgdcnc+6POki2zOpN6
naCWnzhb6hhueEVxEWI+8EOLyJP6nwzVz8HDIxdZqpc4MKDMFg4QGPr8xTEqYOLmRY8auK/GySv9
PH7M/gEQbyMDEQtdk1LoIss9Bk1GlY/bDB4zNAJr1L9+wUjdnBTw1NXqSjB/wgwo9Ky1nxWt34Xf
bJA22AkCd8gWUOGkrEQ5xsWQkp/ncPPpi0Ge4+OxH4KstdXVAAdjs3ki3het1dJLvyUFb+DKzr5b
d9D5dkdZPmsWgeZaEkepv6GRNMgS1sVCP1h3GL+sLMjQW5N6c2XzxMwM5Pte5XqJNxNC8fk19SXy
aApOnthiBlyoElhWIVcAgXP1Y7pueiUvSI1RSkUWUmcbsh/2XmZB6zLIbYHOebTfQ8tceA6L/etl
ThS2uBrp1RcS8HXAnsNkv520zEV5RvnslfLwMa8MFhAiCDMVUW5duoJ6HRCktPFbLgI5Xj0yk0eh
TEVncxczrCTVWPXmpAFslXogHv8hMGTpEJglssqnJl+gNCFpXYHBf4VSunMj4aLJBuYRrIxDjtym
5daJ7b/H83ghYEL5+MCYxRIedZ9tLryfsmTjb83/cBxuBFtUgJthGktbdnoEaESwzYZz5y3v3elP
DaXmpcSSi5mefWX7yYCijQOV+Nc5PfKI7ptxZxyBBXl1uHITTQTrTbyQQVBE6I6dI5DTnPXz1PrP
v0aBQu2SdQJsVbqT4Z2wJ7oXqXrASfk0rGZEmcgWbFAU2aVEpn0YvY0Y9Luvz2wDTqXEvL0Kllsw
+GWckQNd8cISHkDkDdIDkKOMxaMJFaseefQXPpy35gC+AbF5+gD7y18HojDT3cRFFg1joTeMDNSM
WfmG0PwoFqAmqgqEyJM8rEQVF+CpNtGxYJHUY3Brxt1KLXUb+JJ97UocOyJcJS3qxUeoGcmO3acx
/S3wgRkXnDgzkVS4YkCtssjKw6Y10PFVtP5aio2A+fglZ9obBFJBGPBRD5Gyngy5Ky0NZn6apPDA
cjsyYTW035+39w2bABQ0Mu1ca8jVSjtHQk46N0zab3JYk1cIfg69BaEzajpck49dgEyR8WYMCSwE
qcnK9iDjKwLXN89S57OCUkceqYBDZ9mOWEzcYfL3suYS+v3AstBCIWUgrPTJ45/VDgcO1vvPEEX5
+1gYtiyh7FADk5mK1pvt/JGE92p2BoCwtcWjKOMMcOKJlTxyb9WTp+xtqNlMA3TwlqYCIlh3st20
2Pq2fv/wB+PtB3Nya11Wy5+wDa8kT6jbl7ies7L9btHpm959BPdAZY+Mve0dochk9+FI1ohtKFp+
aedIgCTfo3R979UrAm6XM8AQVOJYrJ3lmlUNK6YITDC6j+Gke0rZNFfTl7Av9YIDQ15O+L9bRqem
t0ZyOzXNhkUEjgFpCe/vMB0ranFxLhowMX6RICWm00FxeM3sbnzvoGBOKNK7yPZmjyotZ+aMKaZw
ejJ3WXYXiJ3BpPIMndhvwQC8wPsueJ4tJWTilApq7fZhDjS2+feMS1jhD2r+IkJJ9eADJUnkaiUp
zjvdgeE33dfHpV2AUry5Uk7Kl+f9zQxBBOByj8G0Jfqodi/rYesKSezTSuzACwKF7yBQh/zWMPIo
aCIFzifYyQsXsBVw8zDLeUSkwruUy3/YSWXCUrgXgqDd4pfSujUW/s3nF+aeTm+DCihQfNzb2Gb5
TSSpzGC6nswxpRCNe28ypjGrDNtbNkG9hEVAGbLf2jRJXZ9kXYtWmm906XOFMy+4QNhSoRPxECZK
RJJzUxT+GC5ewEf5Ih8wtLQzjlAVGCOBR4ZpgBSpu0tNzDsT+rQRROdv6STrhRLWql+oxofeXfgl
1OLrwGxrV/fX4uQ+uKl3p99I/VTuWEaoV4NNoQeTiQK7Gb+hVi89jifXieyzu7pNpHlaFolRQvHG
+Ax5qNuhvchGSdprvdBKdjujk0rsqLfH8taoZTPcGhlX081KIg9KKknf0oMH60jNv5js/ZwEWw1U
ubD1PpR+h4Pe/SFQmgBt5gww+m1hScJoyCG7KxN7ASobdl5SpBIN+BDBEOPd8ItO9WtBLRUyAVQu
SgHLbjLvQz5S8YZO2eddLJ2PPkV+dhR7Z84NCDKthv+ds4xBl3/vP/BEQP8K5XCj7uQDDI3fb1Vb
8xM0OuVnPjwm2vYNxaNCVuBB0nc3GFJjkc8aFAhZni6QuCKUy3VO9VXSU5WXNCVeAGq0O9dd3w5z
oduazliuWss0sxhVvuoqxYGQKHT5QC0dcI3/7sCdWYqBjcW7mS2KuKEgVzNn/CdHWBeaorSzzsUi
xdyptY4/JkHrFyHKXIKA8Hgc1OKF1Qd+VYahzARqQ3iWmIxDko5GEbcZdmdkKzJhTmmVKyFbyWyI
YPvplefPRI6PnFtMI/gpkCP+DjB9mwpVmxY2ReNUyxd6WcUHABSOfV/af1eJMwU65HM78EB9333H
7OxJViy6yUGolNnQzn9a5b5QHCcRjV30fDdvINhmUbNvJ9DBvfofwLtSELqGIcWVTMjdf0RM+pGK
wlNMqXknGRHnfg/Kww+soJ0o9KY/8w/UQp8ZVxRzL7aDu2KtV/dRg8B+Xdpxht0asixh9g1auWvA
FjToBeGCaWI4tFVralxpPloJ7ooQWal36oZynkKNEHE86bL8rRco+UZwgmyQo6o4DgVibN++ov8l
7AbnmdaMvjBIPIBz6WwpgXhade6XRz1J3M9yeEiKuUkCQug5h/jY1/SGmpPb/NMcnQOQfSHAoR3R
MXbN7M3YkSf4oDA6firNqlSjxuEhLXbhuu/BVBGSwQiqirYAVKfVRMldGTzjuz09z4zoNWO/qe/X
Z3HfHbn9OZBCAkeIrVde+rtb4BHMNX/rMpchAczv5sVMVDv21K2J6Zm6f7ARSpZyd/BCNwP4cjsr
LmRKduQ0hk0Sl0jnZQgg34wmY4wVTH7Ki3/JqRGPXRYKFi+iFNIEJ4Dr/WzIQY0NGAhIakJ81kRI
tjQOSPPwBiqu59/T1q0zWwHHiEhdB4DfEUgBmztix7y3I4TSmPTlLJYz7b3bHFHTLO4zyfWNsCpr
1lajZnVjq9q98X3C4OiCcZPUb5BcHDaXqDhq0wfzsSSdvF/+cldIhj969hQHtivhLAhRFeTY637Z
e47N5eGWwd8VykT1U082gEujdsG3JEG9uLhetWHZ5pb5jL+vnjry9yd0LltQrRVpQkF0cowfzTTf
uX7piS/lzpf94uOHbMdfnSX4BrmTh7vnA9gADgoQJ6VHJpK757Nf6WC9Kr8Ee8rW+xqi3sF3zywS
w9tm13K8kGW6G6ZTQHQY+fpKLj6inXRBcLGjwCE7Earw0WqEod5eg0Y/gsr0z4NiYbj68qjhekt1
uh7CI98ZBQIyro3L224jcxdYgLm9LLBGCQIMVKHZU7F0j+pQ5FqtaRIGGxM7rQ2nU+GtxrSOVD5P
ymocHnOtyAAyoE3jLahfqV88HzunxjGsZQbMesmHNOFyVGhOYhY6tz4bN0E33xXJfg4uu+yTHKrK
rLZfdNzMPaUmWsBjwrEk2SnqfOe66lTDFKTbX7NcY+0n0tCgPLk18/2Jiz6gbDCY8SzAHfz+vcdG
bu/G9VQ0CDDMqhDE36jr9Qhz6680Je/KZyj268z/pMmn9ir03B8qAbA2brDGKngmbSg1WyAgmZS1
lLGZ0V5XI5paoKdnjVTo67fY9RpQqYjrXGfAVKYqo/gQTFfR6rSGuK6/6zPHEwzB4V26SsAuCqJB
N+26VcuG8T7qPBsF/PCTaPE1rauQxtiWwC5ThpSTA1NM0kebgEfOtppiiTxrzRCO1Te2n/OXT+f7
zPrzFqrw+b3cCP0K232+u+uT/AgtPZhWgLxiextIgeqFwa8I9Fys0UKMm3QmgkCKteFzvDUpjviP
n3gOHUMdC1sCztiU7QIBEie2EiOKfFVHQ6PoIDD8Sk//wNxnbw9nk65zyM00/6vd60PzDWHdVQnz
fmeHhrn+NvuBEhYKtNTeWgURMQWw7C+lOKZvZ3A2cpD7s6MJkiBdNX2ToTWsJ4sWtz+y6uKy+9uA
30ChW8dyGLQFeHU6VSNT8EM0BP3OGr+UAay/Xdp6M3YZnn5O/qk1ukKajKL2AiIIx0qJHHaxuaVl
3zDA/ZaTTkdd69y3JoFfRGo5IvO6NoNBDjehU26C2zvSYbzFwe0PEIbPaUb6t36F4cu6WwadBEHM
tOWYVP+GjNBI2EaZO9so2IkbbTmfTUMceFSAReFtQ2aO7ZxhBYIHHDVDSMMDJlnHDmBRWD1C3mWA
8eB+69MYSD4qXN2gxnHdm7cWYMGXRz4t296CSzRlOSIYZ2aKWC4nw9/gsHSnI6VUKRmJg/VMQ/QR
XTxYMCg+hCcmZnOKpiSkVlkahJwpbQc2tib39hnoUhK2ahvjC1ey1NtbUUiFU6NgnuTC9OuS9nBV
Dt3tm4FD2wiqU2bGtcoDEpr/Zq90FdTRo1UqWDVThJsK7rvLhpKbFNavDKSLwrJLiwyPBM+/bYR/
u8/ymd08FdIIXQ+WlbsdR02P/R3X+1xZtAoVvm+uDgUHG+LWBu1PrTbk/qu49xjB/W25ViGJXmPu
iDknmDs4lqj8mn1hPpB1CoIMnGw/+0ICnLF2bRe1VC1ocFxdBryIDU6eGrBpvl/smyLs+ZNRxE4l
OpNa69dChpCUk2wvFKnGMS8UuttWrIOfqYx99wVaaFSVj+gpT14KAvaVUoysAugOVgXNT+1uhh2C
is/Jus5A2nuUYCB0L8hS+M0gfUgs1pwYZq+OGRGX0X/a3yqk6f411w7gdaRWy+M7JjCS5N3XNzyA
sf0S/p0ujh750aG0vCO3ibn+cVMPeYNoetb+CJ4t76etUfXSMQDE6JQcHlTKkQtKm+jAQ2nqbRHv
8A1KQog5o9wM9/Bu89wcqLvlZdVBS7hQBlZAE+vMiBFOYKLF7CUo/F1SR37kmneVH3AtUs0Lhtm6
u/YST3cggN/rm2+ngDY2mBmEkn00oht4q2tQMTFXjRjCHpSrPZY0hySaQdVC0dvHvANss671WrTr
QzcfyzDymDn96TiSHjD9JYMkHtzDZp7SArepUaUZHyG2IsCa+KA9j//OR5wwkThSOevWGcbWs2c5
hsadRmaJS0ffzlRZHojKt0Vxd0Bj1UFNG39CJ8lr7y2PbfEs9U0GQeCrnh9+4cItlVhy6y0k7QL3
/T8fEW+fYQwPZb8RpDazI5wLwdOCXHSwI/7SqF7WNa9QMuohu7kGl2tljIbJHTFcxHhcXNngEe+3
RLJC63VWdbqeReP9pAb/pYMx1T6hA7Wci2PzLdx6MOjK61C+8au2soJq2v0kYoO/WgTSUIcmR5Hx
31UJdFF9VNa/iWvux+VWyMYfRvqW3Eajw0VVOGDwU0JlC0VBmNWu0QkrcaEo++tqMFnwGp9J6NK3
+lln3QcqYjtuUnCY5IDqFGvYHmgeRLyeaRzbkXz7sPA/QzM9NiU1+sP11iiW007KQOKQ7tzYpLvT
x0jYFQ+6iLEBRK9kbGrDshdN+SZpjgcxzAzPkT0WSnMCpah9QTv8Zq8p3oFcdksTEGJEHZ63XVE9
NlIcR51zmkXhhobg03YFXuNyNcGcakRqv5pwM+FRLaaG6ThRWTq9dR438p/rpwzJp0A1As002t1J
NXyQTdlntG0oBaqgNJDkwETfeqxObjlMKt/XzbHdP1KXpDi/wqzymCJ7+3hwcOj8qW2mKMUsUXKV
DmbiSksCFuc2d0EfVC2XLJ8sJfY6SUpN6xZgSINot91zeuq/Uys/A8nRrKnJIlkA3l5l4Q5mbgSp
xaqdfzRePU1FJFz3BpGsRQx6enrjBUz3gRycXOXZdNoXgHtyZRhRBcwjgzr/R9VlCV5D3XP7QsVr
zMZtkgMFhK2AHw8OzVh834nnlkIPTLwsF+wcdt5OHJ4whSbm0fF7xrc3SqLB9OpL4hz+9wUiSMsy
8PK516RqvW7NFFkiH4+0vsvsR+W+rl365YdeUVg72R+7feA9lADU6goh4b5WbUK1IEdBWf76IM9f
CiZ/CrCatpqc+bmFztszLuyTq/faeKD4jDZx3JUs3EqGp8M0uIg5jzDQkS1YmQbgiwfBDyunG/+7
K8KzPJw1FY+wMnjsTKs6yYKatGsP8ExQnGbAg30XsOdldJ1r42whBmZvZ7MDNbQD5nF/XpaRh7c+
qzrJ2E6lKgvQX4Csa6ka6QuC+DJ/hSURwVXQ56Y/GgIsp/C7iogGl/sctuPdfcxQ9DItPsh6P65u
KwpA/0Dskd5CCYxAKcDaYYza7Z/M4A4pxYxkMXYNJv6qK5rSlMUK5g3NCuW50f91oe841/tL7ub2
gQW4cBB1rIfUHjuku8S9OuXcAloY/DA8QHu73MaZiehdfo0rx8WdRExOcCebV5cscekWNi+oU/v6
v6iNeyar4xKFOjEYxmka1kFsYNJHtL34eG35zD2JT9K0HBg63Hu7K75h7qXcJ0m8wZqPh0vzu1fb
SDNPk6v6UtLwnCYJNufI2K0qB1eyRosFw0uVeoAyBuabdpa9ovgBHFCksJbJlqkKM5kOLCQvfsAP
eGVkxyL5KFXAMisdvicdNrRf/2ocWLQ5u7BYMXgkjToRxcYtswkvsmhdQ3EzNxEM0TvZvY+xKwCh
UN/3oB9Lk5zjX6ZpXaxkuXaVIPzKnyJPTaBDJGR3H240RVrX9G7gFpNtbVeuEr9KwUeEWIhFUQSq
tEHiH9NovvMIAi5H1c22HUPsPP3jen19Y4jLM5aGArJVJn/7emmlOAfXy9snndjtkJnDaJGuB8GV
CI1oa5hOkSxueu++ZW2bgjR0ka0ehI/WWJUwJWOkKIXZR+HgSzomGesCken4WnUavUjHFWz28yVb
MCMsC2BAU94T6YLvwRx0V4sg6ZwDXdlh2t2Hgj9EmGMRkrEtClIF1DuwHXK7IcRRirS/bklxpB9L
B+jolEYtwMTWHOm/deIW6R+sdYMOiZFcWoG2YvjEBnRmpWjJFeVGMhtipUdq4pPJevpk8UuY+Elf
gdgwUTaUtIX6qY4YpyZHhfpwhqxi84YghT42OhlPaJeixMCrsCsgHI+35irfGD/kXsatfnQbnPwP
RwkyG3etTRoZIsWu2c81XFl4w2qyZSSdsp7CWBvHosbeCpj40Dcf97O8xMsvReUvb23dd9PcYbz5
GPOlrrcjA9r5/WVvbbs/LCATTKdELIN5VzvyrAqLqYu5S9mXQ1MsxSq9girMHF4pl3Z4iSIQeZx2
otgfFaU+4sap7yiZgc2Q94LVL19i8UBhFFkT+rmfSo9RzwiIZo+jx9nEHuwm2cLCldMuKyBENB/A
HwBztxB5SfLq9tp1+06j/G8G411YcJUUNRpF0kIazWifAKHzj7mSZ4HZrEKf8y6XwlTZIWX64+br
NADpcTFuvur+9+PVboetMxpwjOhnEV3Avyf+TEJ0CMv5ygYlPLFc/vp3yYCeSU0T8H8357Q48sBa
YlTB5sPcHDScWVzUgjmE61Sk7XmT509zPhX87yTJenpz2uZCbMXm/Wpb0+yWjustreW0TrcfZIPb
/fRgylqxRFsb0/kXHk35NPS1BD0eg5t034aRTD+CLATqHipBaxp0/Pz4isCZK8f/Jgfcx0vC6T+M
VypDbAJ2Fcay7m2sGrQb2dF0w2Hut/Ew5sHl5lo4QgjkuvCXgceyiMNvdyrvgILC/0IAnazsGbyf
m8HX4iqKaN7jUJbSCtxZc51hr5WsdZz+DNlwIZ5GOvjA7/z2wbLyBJ6Uyy8FR6DiMP+RfmGWjtGT
NYqxU7r/YgQAcVYYBaNNQXyXOzdpTxD76QTB99TKjuORJgswtJEZ7u52y4oKe2WjRdy+9L1E1ZbM
lae35Rxm4PV+rlBMWCdd/LD6z4tBoDc9RTwSOnQxnh5Hb6bjRNS/5QVnL+9495axQF4Td3KWrnQV
3hLdeGmXzUhXFtLvngocxKpVmrJA8kunQMM4K5NVh8MzNS3hdXyzMs3Qs3MhZdBy0of2DUQmR8Pj
Zhi0de5EOUOkSV1Cz8zpHmfOzfmEICqnMm8/+1jhiDAcqPyW6lCe71ZGNZy7tBDH5qkEunBUjgfb
7TopfTTyJzBU8FLjZMu8n2Hv/+3gkDqFOM50Cf4taHxF/EozUX1TUJHELW4GM7a1xr+7Y07iU1zD
NQH2mKAmGZZKf4t26OlqRyrNyylzVjR6jHUGZXxyJWJusjfsLykw8aJAbJsYaQ1cy4coQKJiP9Aq
5WHlAb0zH/osGGVl3a35mZ1Fb3v7pAz52YNpJZsUjOPC8wlytMnbjjD5xVks/rxjHnaQI3Yo4kaP
a+ij4jgDmFZbK5gprzEXncBJuvSohewXxF/Gddeze/U5ZxGV7JlroQayz4sYTvdRboN+yH/VBaC5
J7rc+eQwPIdqCEp9iUAlWeOmONdWHrADs6kayZ5a5/XnA45Lekh6kGYCDPa1O6ouMaIwpSqzGS11
1C+XKll/PNySr8DPLwZwA6YU2oTDVwowtOx449aFlRzcOToNoRrFahcuEHn4ifEI7EdgoiFcSKxg
27A4qWvpwGeUus5SYylHq20cE80XWgbE1TuojgaYf6sW4KjqO6YSuI7Ty0u8cA3njTeqWnaUsi/b
UfKPwBNh4rY9iyd8D2hqm0mvvAHlx5zpiumoIHGrZJwnVjv3g6TJRBU2KGqPS8vUa2OPFziAw1DV
ZdO+vTHqLy5Iw5F1l0DziwrfdGLiagCJXKyNgrtbrFR5Oi3+yYX3UC8JSdnSPovitq5A025SGKnV
Ed2zhqQYfiFfhxgWYSaiZbLX0ytRc7PM3miqy27ZoJqftoeJa/z1JLj+1GoQIFIrNc0IEhAbf2cY
LcB1sVL47RiYARpFD9XMZgmMyT0GF5slOP4aIKeXFm5D12dKGVrtg+Y74gxtlq3qiJ2NDNRQaBTR
3gelLqbQ5rRE0EGSsiy+JQIai6aHxv/u6FV8U78FHzN1ze2/lb3bGvbJDE/xIK34PU1Y5i5MtVlq
VHS5TaP5KY2o9iQM9XO1Gh81w3FoGYn39oA1JWGXuQDV4NhxETlgp6ymionneFVHSIbFr4uXg6e6
1kMiREViHqG/rUfcTq/JBkY2bEWLnPwFvpcXwg2D3jX8uhCClaARutivI18clb53BKF0sCYOvKkr
tfjiIacHZHgKjzr9VM8nvfobiNLacoydqUJAj97usK/jK9VCgITfsLHMjiiRkmcndnSWJ4k/1+TC
a6ku7wkbJRAtTXRqY20anQxJgIknTG5C6cMQYAzzFB07hTXjzRL0Xu8AHzlmeHQjyk3t5zt69YE2
tfOsyPvHmsB2rYrz7yFQhwaIDmA4pOYX6f0ExwyxzFXHVuC98SJFtdsZ1zQtmOiVkrSMC4bGJtv5
OvGJpgnoJEC/x9wiqKzRQPd8N9Ws/6pHUX5Q+EqvqTI8DFjbFEu7T053pOCzzLg63aKw7V6MRb/Y
us+SggSFUbRsB8BNUn+dTpvJDqFSDN1ZhcgdUN9madJ9NU6kb4O9oOzOIACac2BgAVB0iZYsjbZD
g3KzdimLavqcZtNKMwMt9BOtT5eFHpnguKOaRCbpr9dG2wRniS+srj+peyX6YlxCrE2ELnZhmAzG
Th5P6FwDXdSIIWertSKAx/tzctkjb1ysr7ShgcGECcdBPiWdRYi+5yfI0ssRDGvS3XeaNuxa2fQz
RkgNmw2KI7aRKOUSZgD1FRtUyRKXGXso3n/5lnogajPeIKB9s/g77C+ve3YVaruaAFsKza60YW3w
Kz6hKd3cPBPGbG058A5vZ7I54hl7JjLkhv0Wzo0xg8COSNHrXD084NIPFdjFPoInXncK1xr5UnPc
VYVGXgAil7Iu3x/w0ww8eHaS3RDskfYIN0j7xy6oGb9rnOCt4P6Lcfj+JXjkBcFzGpZQMHJC6JMP
E3cyPHGXfZGgjwND+HYQpUFcPHDDOzoxfL+iXG1FO/ShzHYqcGANZ+hDhwEGgY7vzpP0R2dn7udD
4pXUdMX1DsSzexNcEOu/X7+g/XbZ1Yxu3ZNylhs8M1k+mQqqYniNI1xVAirOfloiXvsN56CQn6Yq
Zf2YrIt6bbhjtI4ygtf6Yn14WfvmkvZfjWI+KVedF8Gg5oFKKJEe+Zzdinm0QAqokUy+MR/hhOsc
mN52vl3Sa0TVaJ+qfuVo0VuI258wok9pIYlYMlQ31n+Kp2R3v7iNY2hFjmedOgQEcyK/KvcOsFO7
iHLADoO3z3hHvs9azVTo67pzxiyk34S0u0iTHXpYt+CeKdW2dKjZESptIjf5uqT4FukfnmrZeMcL
M4YRsMkldUkZ63ADTECE6WsnqSh8SFWn1urJxurjwc5EGawDe+XTQDBmVSfTSZjp5YtFsJboSjLu
APTQt9nWIozzlk5MRpUbsFCTmadIDugc3lKMx6fusmTIkuvLgsJwLK4mRlY50RpCfAvjePyH3+rX
nbJp+Z8mRtUN9ZMni117tzQeMeHO1VHsjbdwL0H5VWUUi9Df73+Y8pquEDKJmc2lnD4NluWArNKg
KkHueMVU7ocUr7SQtPqp5589Avoe65pR2fCsN3ybKROgqRK35iMVUY/xZ4542CL6PX89VV1WxPjy
A8xev61Ux98Phwg/ChYE5freJFwryvWnrRbS3HbIgXDhdGMGZzH13FjHxQKqmaYXL+OMOpDXj5x9
/569BObYsvvemkW0VwS4BCIOsWD0G4v79SjTgdNaE6WHAST3vsL554sBMISrRI5rM0H1+abmAJHc
URsNqjzczwgxlQLVaJ24V9IzpLBh8poeyHESB9G+BZr/nhcrgdBOOlDi6+NJLqcG6kMDuAlzM+Nl
9ceQpD32XyNal83xEktg9qDdvGRrr03l5Y2H2eBzztqCtrNe/C23VMGNWfy99SV4kkgxc6rXhF5c
1Y8T8sjuJJb0e3XdKzLC8iMzqY3LUZqwE1yEizgYPTByA9pNUgkAR/H++4CjOcWeac/ewbcnLfdI
iFTX/aBOWLeeZLxX9kSbrx81VwhQRHUbJQt2B+2UTUALHSUv5AFdICSZj+j7PwLkUGmK1FyKvKjW
LaXMdUgd8cVi0PtU5dY4cJ/JoFPHG63iXz33/2hrNXKplD/fK4p0W67WD9WK2ivYJvbsx7FOCe9S
xb/Sb55+JWIQdE/1oMP7Am4lKzo8ogVZwmqisyaluXXI1qQMVMqTKskm3zhhOmuSlgDYZ3q2kqoD
6+/iC5svJE48cawbReLqkBLsL0Nv72QseuvhahLSJRo6hR0GZuZqvQTAG0lXDgDEZYxHL2NbFpGn
oN0Bf0XoBBFViN6oY5rFZ7vWx6nUmLkWFrdAf6cP53GAxfEJ3bsKx/hTJSioMHKt0JgRqMXfM3ol
mMIgYyEMRMR+vBYawizFnz8/vGZI2PFOZOIgEMaBST8kSKgASxtasrWA7Ct7de64n9aZ0Pi+GJGj
75yBpLUtacts8C+Bnzhw4cmaI2+mAHaQTrWnHmNRR2+h9coOr5Bl0zo7gVvVGYInuogfhLyBv3VH
nLPzpfP2zzI4Lls13b5lebyq7OTzlA+sqMt37ySXonSeXYpqAxjSvMjL4p1w0+d3XSIWy3NcE3fq
P6hvLB1jJqFcalxJH7IrRWTsMh81BlOE9oA5QAad6avY4XPaLf9YuurJOQDJA3X+E+iWPE1GKDW8
ab05kTQTXwUd4seDPrWqsetDbgs/AFHgGVbcd/YHrBwtlJsaQ7ha0AtqK4EvrDFiWJNfw3mmIiVC
E4o04c2Ul3+vG7i93/+kqaXJdXiaaJu3uIGw3RoZEjNi6cC4ZAHXd8BLk9YGUXkDW7NuF4b5lS4f
2m5J/R0bUW1GccsJx5aupNhkJcNyXJjqDBO/Sqz2+31tqXl3b2xDA8J4NX006Ialrgw7+bxmmNfL
aX2l+cld3stoEINJsK5nAUBfO3aLcA3TotNXaBsABHgBiXpJUY+oILp/7a+X95bpwdzL7tcMNgVf
PaxeuZEFmWNl1aohuuA4sktvzHlDWYZX9jHH6ata3ZXefrpmXHKljc7T6BBLthLjbRXncLiGSbbf
Va7d/cePi+T8OEzKInS8H6qISyR32UybFLZvWL9LjesufANk7GseXDwHEjnAy2XGsKz5L9VEShjW
W7l8QKOJJow9JVCgJueUtAClI6bgg8VbWkOL9b3GWGaL9ZxKfKy29/E+ZCjPQGrM02GSMMYH8V/a
kFIcdzHL8s1v8hfUw1qL3WeSsnNOsZmn98NHcK4Y+eI+CJsxqSEOX65ufzJ2M1go4ZmZJ5Oq3NFF
J2YOkYYreyOvfiOsQ7LSXOjJiJQf2J3dmnwnIPmxCFm5z92slVQxVuBHmuwu1NTuG951RoGqMF/l
7nI0IbfdDwEgoNBqK9UE9pXk6eQjsOwvw3qkYJtRcxPluIkEFy0rWzaCiWR9dgF0mzp5sn7fKI07
PHA6GUsfqNliTndXu73VGGteXVp+ryMMfQswoqptp1Hd0sphSC0oYFVESR+dqZ5V9gYs5w62i5CX
rV5dmWevCjcvbl0tCwSO8P5tHVX5EbcQCL4UoRhkoRVKRDL1ke+0DSFOa+806Lc0g5HX/1IQ4Ce5
DmLVkabmPHCeJWNpq5BL/QErZSZj+4HseoY8TfsM5gvNxK8J89pQox6Y3CcFpjHlZRJG5VOixyUH
ibQYdr52VZ6YeAxg1rdSRdVxuUOowXEHCNFV8HnGAFZwqeKjyJUgIC4WOMkSiMvSBUcJOkX6lL0R
p2GIJYImRi4J4k58xflWCqddUQWJ7D00iZqwTkSj3YLsOytFVwOuLtuqwGJfItcY42EqErgzHTMK
vVjC5wf9Id4Xo9qYqoi1rCPsUr97g+Qu8K5pduAChCfdk39lkHyJMjPSfA8NpTew7FQEjC85C9FX
EJQIIhgAZq0NVms+kA+9n2wyGsyJgcdr/keAI0xs7w2WF8m0E0FYXIEjV5QanzRIYthcYUn5vzha
cBMnyQe8OUmIDCnALMDZHmKqoX0XfX2sI3YLkjEQN19lCD2wtMVzGjgCoiAoiNlRLjzFDz4XqP6U
Ugf/3gbWHKAdr+mBlVZOoG2B2KCPgHa9oGXeAmvvL2EhVpWOOvem2XQcvp413874QvXRKT7NaAyx
iOtCaapKQHJF/D2o6AZiZpDg+lZxbb5bIAsmU/unwGLc6wu4RpMc7Ia56An5wwRgGU+COmGFWNgp
AJKnGsspDKUvXa/4bDKRFL3Q6ERgoCGxjFytvRpA/HdH9DI4oflz5+bIZ2nlC9dxMyLpcG/qmgEm
w6S1uRSJeVdWh8ehXb6r0qZTuvZ7/22H6Vbai9x+M0doLppOh48NHgvpKpimsJcTLNO7KWSXxQtN
r0YqxldmxVWwx4TW5TrlYq94uujfGG++Pswp2kecbpQDZn5v5aGHnuKaiBdroGt039ioZ3r6R5QJ
apPMo5OB9WJTUYD+D4WHAwJYPSIDjue9qznxCPGPHSZxS+/puZMPOmHoyn9Zcske8dTje8z/yf+e
7HHo8eYAuQB/vehCodhU7Ion2naaWcbDpMU0fXbNtOIMrK+hRFCyKRIpH8MzfFYVQdH8tYX85m70
+3hPTerUedt99iuAtaVjllCT4SF404DIhQ4BdbVRpmNTdr3/88dDdUHuYPEkwux8TkyZXJCAKNO0
nzMJ2BwphQ+nM8e28WTFgsRc1EMgWnOY73eEkjnh1gTV4af4tisQTEXK+Rwz8HeM10t1yxvGzP1y
Bbk285DShA20QJaCvpMDnkOigwpFAvBzoOd0pqw7YXF9s4tOj0LbEDlJNE1ngzYfjhToq4hbXK9x
X7q5lOLIS4NWP8JjtnpBfr8pdVATpEOaWjEOBki0TR9EVxu2o1WvWWLP4IEzNwUmUjDTCcZa1mhr
qvSJhYmz83Zy760k9Q0ZONTav5RreqPste+CtWOBBFK1xpG0thO+CwXQ5bQ8LBtCRoQS4Z17lPMx
f/6NcwkujBiLqGksX8qxtJyjd+ZssoFq/ou8MSQCMOKaysfoR5AE3nB4OHZSxgeV4HsLgkkFY1sR
YF76wB3BtYRWyEyZVuHWvTGf58oS7z3fetkTJh4bXNdvhpBK7AvW+EfXhVoHMeF3py+93/KyxPUu
IQr2XW1mpDIWhk2CYyZ+W2RBt/mWUs0hrI8a+QkXg6PfxIhfVKMPXolyrhceU85Fn7/1rbpenDXP
GL79FtsGtAwBe2fy42KCXe6Z04a0w9ZxQMB7oyb2FnfkeIDE6OnQxqzwDHWU4LHCXZuosxrQje61
pD5Th0ee1iZU9q4PBWMxuDVvkH0siOd18DqIufo3VDK2Fpe1KEosV8HCa3p1Ur6puQXO6aFsN+2c
tdKPA/LMIezOr5WXEXo0v1uFVQ1RB25XKAgDKA6kntp56lj6FCHvrV6gml8vMrZoE9td0bjO2Drr
KBURaJmeoSGHfP/nfpFx2CtyVsO1qQh44gwB+fR/F4TDpD1sLub94uQUTfWmTUpWq5TGpEzqbosS
ad5qZVrsYi4pfQtSW2PPWX8u9U0p0c2beYishGW2O3qClZXB6/qB7S3F+K0gL0/DDfFBImuOvcgS
umEzm8I6NnmSQ4iCRbXNJgB5XJyyrnbkuwc/qYGnUn0lY0nm+wgDH91LxEd/2zVA+eM4/oqviqzz
Eufe9PTBaONzIlpLVvtDUSqVm5ib5illy3vwXBCq6q5IR8VRCGt4tj+L9u0YftPR6QLdk/XK4WiA
Bw1pYiagFCHBmENXMZ9sezkn3JLgp63Tkoq0MEI5Bpaxr78/0PGtrf2VhINmUmhFULk+YZvlGMAc
XuKBXdLVbvRXJdph6wTnKC8TtqR7eNnDTaF6i99sEwoaFkhnPbn3Z5BDiLYVEpK+N29W6FzsFTYj
xMCEFNkTcHVGik452y9bwYvyekDZmi8116Mfbp2Vf1TEsedUvsJdWo7iVwxjDf+bbjlrRRasy/AZ
xtuPPEMP2ZZWZ0ugFw0uIr8XXmRgXQMtdCevelUJjy5eN/DhiXSZBs0pLECMUEP66ip2KWXPQEEc
cgIsP7c3bscJTQErK0U0mqlTx4rID+uMeoYUlpbOVr9cYKQZF2bn0Hjkod+mUatf5HdPiFeIwhF/
vvjGhnMEI9a4btARBbT2xBjtdmfWDioW8B2jk3GvjEerp7sM5a0ieAcXIGLbfKIk0tCPIfv/an8f
p+NMf+uFcB0+CrlhybGZ/pF3PryxUYQj+9BMMJoyD15Pt0rTNdbUIFJNV/3C5diUcdtIpMxlN9w5
HkJR9JB743KjB2b8y3p+5GadTUWn9ft8Yj9pA8gg795mwsJrIGcBWUyvXVEwZQQFV/J5T24SwQ2o
MiR7pQJGmAZgzXhtX9nKJr27Py3z+rzj1FpqI/wdHpkyWjYtmpGCJg8KeBJV+QmomB/WvJioV2Eg
ZbE6gZTxD/BnAXD9TudHKhBdwsCpWfLa8ExTsIqHudQRbbZpaz8kZ/35azt8/4tBc6AJwtEiKjlh
TFe9U79BldC6SVTp0pq54JAPji94n4VjmmjVFSIEelI74PzQ/FS/tx7o5eWT3PQtfloyIf1jhHUY
xBPmd7iTppht/0Q5bLEOedlJOyT+4EW7Hel4yDZi8h1CBdjssyPGfX7V+XN/9vB3+wJ/vELT4tV9
lufy6Y+uHeNe55B70NwAysKBDnt23BZCQ85D3Bi/bVP9UETyTKiveISHl1sbKYQpWVsGuggeP3Md
JI13LSlWBI1AcVPV4aAsX7Cs311NC5smj+DGs9dHZoTsnd7WTs1umxM9QX510J4yaqAQHkx3Akyo
zMV02xmNfexGbUNyy3n/92hytxACqCeWShrj8O6oJuVclb75D73mQn+p+EwFPGXp+XLfRMjCpCvT
I9Quw28hPR7rjR5l98bTNwJBbwvkpUkJvaEYdQkWfGAblnU5VzuuhSPa/ZeNcdr+QvmjgQ3umrqn
CUxy6B2ZGnJZIX20Bpw43sxWMAnHDyuMjbrfyWlQwkCYd7rKBaextVnp0a2KYUH0ECo7XCAe1fmD
tw1ppJJrF+T83B5QySrKYni25R2WVuvIMhfI81qRC/lTLLI0ANuxN+tS7ECHZavs094aTPsPAWFQ
2OoGgBbakEQ9Xuy3ksgZ8gmDtWvd1X4Jmz8st7xBayaNqnBU9ZtQUc0qqJiJOI3rFifNGXxWcM2A
otk01H3xIiUa3kqlc8jlCEoHMq5HGw/o6ot3UfLtZpKNkKL3aAqSYd9g9SB3+KQY4M4pBzvjBnri
VZgZ5mUM72WhzUOCv0fcsJaNVeOoS5tbpVgfAPegFTBQE16PsnnXpbzRh+73c+xMre1e8eZEhr6G
bpr8T2EV6rf+504aU0shxfnIYLSQZJN7OdkVCzgFNFqW4gCnxaiCA+Mvzcbe+D33YLOMJwXTgc0d
PK/B/MPhw+83koMFwyHrkWVP376+qo1GaChAur5PziDUowCEYbQqj8EXKNrXYt77/Tc5DE0cwymn
gL5jjZ0Rdi9ZHvm3dtCN6xTPNKMBNLJ2x1B0mMN+ncb5LG3oIAva5/EXdHJwPDbv6C3FpJaS4Tnu
SiRZ+gp3CsD5RiSJsTJgbm9pmJi2wuX3Qahu/DRh23nCGHYGkab4i+WxxAtmo5/yFNPE7LgHsitr
I+K1NSTrjlm27dbj8GwF+DgI7F3oKppaYIX6t+gRXPe/jD7E8o2rCm4RdVXgyPatDVsxEveVTqSL
9H1jvCSMRFGycrP8l+sHNVulo0/T2BFcEpjIPySLiCCJg5lBzheBCWxVO85DSzbkOGopM+L4VZ4K
TbUtcZ37/5A1QOFUO/GgYSkqyMe7sedWT0opb/zDzYeN+5au/tlHWbEEh/rVMpKOv9jGGJJ+1cBo
xZU/JfpHBhrqHpq7Rq6fVXs3SW7jk96PaMDTFtHcynB7vMkpQ9AIeY952JY18BK1Vx/Jir8EnoUl
SsfeyKItyr3BFdqa6JaGxlcq4b7kgaKA0QrQW2rkBSNijT57Cdh2a4zLX7dVZt9nCpKb3lBZTPxh
emxQYSSpTcjVb4e44P4hmAa/E0oSikF9xEH6f6Ovk/MoLJLf/zCSJ54kRB4f/2HO/adbnpaLTwXa
ctKp5+EDP2HYg50CJQ0KwTkeUK7+19yBm4xj44eVwNfELBw9B81a86NjJ/Uy0P130l6ZeZ97o9aW
DY3cJiJOrBK7ANNCZr9b/rywY5H6ab3PQ5R6+L0tp8tJa422RBKnPOCaGlnDf8H2+pJHvB9rtRuN
Db3ftz4Le/Q53b1IeG0Ay1qTgMVvAL82WBPdf0pgyBajqYrZOja0ikSYzY9mh1wptj6z5CxrQK1O
ewqDn2uRXMbw8NU+LLZrhOVCgc+RxWdE8V++gzgl9tbbPpCkAlgCZveuUilsw0I0WxyvHbTm8sJq
NdjhRYzUlNnrYChoNCNW6HpiIhJNhSutv/+QhahBdYURnPyCrbeaMiPmQ2CENR72fWOdXszb2IEq
c+ZCeXqDEje+U5SDzFyG+l5tpCCixZ4ZL0EoBtqlXYnnBHXve6VWNAMdfxk+78Ib81qn5ffqdt/1
gXKwkTpbn7+6HgPSuR8ayZf5EnlLqfA81u8yNq1z4jCI4gkkDeZzYnWs6hEmfJG8X1WOXq1jTSBm
Qn0k28aLIZjWLvtGUrh7un0zRECW70Grn9sfeiJ4Dl18NawHzYe1SwnoiV84jTMYJXC842CtAQgP
X4geNfuHO0SNwrkxRzpFHFGigowG/QN89NNMwaZwObClhU65kw84kEe9lxaAzi/TP9IAoHE6YQCL
7FdLbTAA4fM9t7dfBiBQFhGlNTDhbbUUdaL+F+ckDqKj4iu8YQOKPlbhEdN2p17AVuZ1qvk/xeMS
Pzj6dVQEeSaJPQEOOiujrr0h/7HBivM333B3eALtTI9DfUEGrrKlbi5YeIwGK7SFnrJuuTkEeFoy
tbOgTnkHTvG4XECfj87AXRO08KGXo1PVSIEwk+Q+BF5xDCdaV18tVc9OUKLYCvntXjwtwbvQcCGy
0X+g2NRAyi4TEaZcdWcqf31C26MQitwgp21JK81p4Pf6MlK7b6ylP5dy/G7iWKN+d6dzrYR3PfKV
nN689ebhYRMlEmgP83IarOYJ88l+EiFMevrzqcXVxuJpBfS2Z4lSCZDMdxmwOjp4ndWa+dCtGzu0
0g/PGnsYqJ8FbvCW9gKuWDD5D7t8dc1YXXXYPcriXnvuRtDbIZDbX94LNQGJDlu2XC0FTH2Y8fQM
08WV3RjbHH4hQtNgXJd/cnfjEuhCVlsJfSur8G5L3KXfy3izpVlIKnkQUTJGTZMnUnk/7PXFGonN
5rQ8dq4osFqR+urF0FwZFQLnFjCY3Hh7D7GFQaORAmGHDWFdj8kNa6mMCV93xWvy9v57ttxYmIc9
DHBlzYnrhscxf7d2thJuO41f0CQfaoTvQOCLPN/Pvo4rEMrkhYoqZ8YGuBcCPiJnvnKUhvUoVetx
DKHsxz6lnBzZeIC6vAs6SU+0QjlNbEKMT5dGL7/U8H0FRTAlfLXxI4O2jp564HWQcCSwYD4RVfem
0f5SC1N0nMWTx6/gA0yDk3/gD/YCLmZyaEdwZQQpIS17+14OJsW2gatts+s4UHh5TMbuyNNwubws
S1YeqwMfBJtm+4/1zXxTIu+tog9H7x9GiWqbaLVERleJ5p/fRB+/qJZLnLq2fKSDNBIDpcSoTnbb
H1ORupwdbQ64ZnyuHpTYbHuwB+hhdVAV4oNazED6mENM9yyXOf+1myJNNeL6y/1KMnSnMKe9T3VV
MvSdxHEyHgGkkRBddY7okZKvL8zW9eUuJPAXZhcZVGfrFIKZOe2edyKrSV/xbPmJxrFYrxvH4qPW
YuAusKXCatM/OAvY/itDr3Esz7dePY9kIb7r6IcbklPTH2DHrW+EP5PmmlBVP1wzdASYHGoz0iqA
jhSf7mHXpDg8ZEeUwaplKWTnyLlFyvsF2RCQjwDt045Np+MLEEw69iaFk0VZNBUS6S3oQkUieikA
5nWQkYbdhlsUb9YeuLMrTPhlvwigqdMlbhgre5gfHVPw9Ku1zIUH8uv3THm/2nMIoVD3P3Y+h8KM
hevgGEMxdKFaYxL3NXTUGG6wMqQGfqFDdxs2+f/S9t58L+Ux43ozyQ8mNw3yNPXJqHXyMtDm51GG
dZXiIFBs+D1tM0FLRcTz/0mB+Hs/1j2J+L/u6YDKzYTe9oEajpKvvVFe2KRw1dwJzg5h/GhDizTp
m+dmRK4pAu3x+LhoYE6lCcQt5rHsQqAN5wWk95W+dxaK+SKmF6lCLm8aXN7j9nQfYZNomE/TIRip
l4wfFEtvP8zGw+xO7/j8/vSOTcpeIeyKWWfZ0ZbcUygo3RdBHEGsSVRtX+Ji90a0snL8h3ZzcJaJ
E4mGDvVkI0npkBV556B966Qh1xs83DHyfoND3ewcfN1bctOhrSgBfv0WZ/LCgfWyeqn+C0P85jiV
j+BedNPNzcsk0xF6FHjTFbNWM62sL4xwfbx3BoM3gfqnl9xP+kBF5Jjxm9YI5Nfcjg1rqmYZMQbf
0dcszkcE24i7ZbDqZOyWAPZjNI7uYLThEm6bawbtq/N0XxfxvWShI1yxNlVn//2JKC9Dbc6P6r6C
MtXM9rx/F6lYCmCSfLm865ilZqeHEjynoutSGzf2gRMyvGo2urjSJFBTHa7t2Nhtq4RxrF4KiXoj
tYxyaavcjK0TN7ci7hLgY9As4vPxXU6/cpUvecCfwDI/+4YKx5gZ0ACHtQZ8yV+NdO2NhlQTWQcO
CjgNo1eoJDEem8hSZVSEsKQby4bELbke7GZIezWi1av7V2h1WE+i8qNVwlVj7Yuvnx3ObpzyQ4La
UvTZ4OX/hIdS/mYhmfjJMfnhm+/IGRY96mhCzldxVPDQRmFxxrAqooy1iIz8dcLdWSHUx3GznY8j
TF0yPMuqdrOQ7Q7KuoTuJIqzJAL/vkT9v3k1GHW0Z9d2UY52JyzxCCEIB5UMNXcBW/FXogKVJx3v
2sKVW/0gL2pmgk07EmvNfLuNJej/UTZEGwu7Vu9NZkPu5n4YUvjAzHB+m+XhOplq3uzFRQJ6eAnk
Qh1jlvoXzKNFwOzHtbQBnmNdx5M2XtvHnlM+6YIunLjtr2Csv7beJND+rIGbtyDwq56vjjmdaRlY
P9cMeK4ci4aUjQgmLEp95QJcyT9prm+bFUT2imWs86F3zLO9jZjFmUicXkJhlG9xoVu93GrAdlcV
oCq/L92m/tKRqkuyTd7JtawwP/cQ4Nv51sf6S648hnLab5A914AZ5+r6Tby01kYuG4lCoQTiWa0X
gHFT8Hw1htmfMTCZP18TDW0A19SqxfFDU3Ll2nfWQmTTbHUMWaS37NEU7QnFN9oROyVM3JQ4mFd6
XX1fkUVR+cOXOTBiju9mh/JNUHwjKiBHgy1zuYYiScV53MjTicBnzDu+dd3xzed2J/jwcD0GtTln
OK7DjqDu6nXi6W4tW1fOKrp1mdqCAjx+TF/tFegzNaltvn8g+758JSZFS5MqMIvPcxvxlpbcZo5r
U9LRlNdWEbr1K5+e34Wa1ZUzTZCArAkLC3uVkhQnxCFD2vG7urzulbNmo5wv5b2ExKifARBNPDo/
PjrxoNFPq0hU1YZhxnODQNvCm7pJplZbySQ5M1RkFNQDKOrhdcDxhpVSIPm8mI+lw95+Ao1C/TOu
mP/6faqh5wqzNoLA+hCxMIIoYEiR+KU9s5d38FA1PHJ6XY4Kr2AewY03qwUxEa5sCFBp6TjCXJR8
4iGrZPI9dZlKFgUC88/FMhcV2ZB5bGH2R2qr2tn99nsmvq7n6I3SByPBpEkz62w0qRNvn3z/QCvq
obM4PMwDLn+KqvsjXTrH+eKOXvOZhGxOL+OGxarXeuF0e2yiMQKJ1DDbpz13hf20R66cobY8o5K7
/dh2SsDMpf/KGFRXFfJgAfBhokkDmgqNWjzxMdKDSizEFZfpI3g9bfluoB++l/rMz4hTy5G8Z98x
YHWS0G0Ui3t26UrnqJXk/60JG2K7tKBaRKSysuoUg5hb67JznQof3h7+d0BwAlEEfMYs9RBvAZOF
/d3QGn0uEu5saNPJbLnLIETPag3BB/kbyyXI6XUpaaOxol4hJSJsn5cRdmz6/RYXz4G+X0ApF9pE
RKeA9Q8EOB22V7lqy/6EcdpHolWkLmN7yFCugICwNAkSbQoSwQdd322LC04RRqd30peBhZLammWA
BiQD7LGRmmADGKfmzP2GlbNyy9Oi2kukp0WqIBS86CKWJHcfN3nCKnvg2xoNaS/lIF65N3zZWnbN
RVP9s0IVL8jBDU7zDKrD48gj32juUn0kK30lujpPCVHhenbha0ptCQWqVsCtP03vU4OEeujhF9Jt
oN2bpLzskbdyG09Z9jFa7A/VsRZ/C0h2s8tBjU9Dgy7a9zuqO7gZak6DedPl+AlRyBTr9oZc75KE
S0UWC9JkrSu3IFVQMCILPubRHSMk3ABs9M4wvjFbt6ytyjFyPDOsxO4UL7Dyoj8VvSVI+mg7Iznu
8iqA/zswWS9ylol6XMTfZ13GdcrOehSyH37BOgPbE60X1sqoMi1ooMYdCWGOzPwKKKnTxHT7j7Po
wBmRKcEMcFdPeh2SGQaZnrFIn14JsvofXRFSrZ/wVP+OXARsArnDfLEdjgHL2OpiEBvTLdoWgcCV
ZzGQKW6DwWwoYACgD4qNHz0kcljMTTAfXZWweNm2Qfuxv9m0+ahkeu8CdAVwyV+It2ou96BIe06B
eKXUp8a4czBm3aDq/DhlhByowU4mpoJK222e49NQ6nM5Yu35+DJqtdIgiJ4Zvx+2RTWwYMZqa7pS
SD78Cjfz7V24Fiedy211ljxV9QP8kl5iPYXszXMfQaOYYjSvbrMHRoMP2OUqXfiLSnwuh2YcaxX5
XaAz7e9zGtcaYdzjFWO6TphZAJzeeaXjJJJhP3EFKaQwzhDpxziGo59ifQW2A8GG0OBhYmySg1R5
P8d6XOQphbRHtXmEGj5JSAqYXu8cKmPtYiZxwmbCOHb/1UcAApNmR+kE15Sx2wA3AVZk64kGyOWQ
wS5ZEEl84AtnmoUHLBsvFlKyugZvGF0Z4US815CmnoWhbxYhxc+GGxYPGzJo99wK2TNdowtdpsMM
DI09S0bBK7FFJ38NWXViVqMvt9cCj6/0M7khKs6fcqMSMFRJbp3sA+F37yFfDHONfq59Nmos/iuZ
ZE5sUCKf9XCF1wayWk7zsh50LLUoXsDYxJ0wvEbt2+fT+rFVYjapVOsMPZPU5QAbQvD8ou4RpGH/
8he0/Mo9o0lgpNTeO0tJPsKRYikahVHmWSpTfDZNkWVQPk/US4ZHvTQdo7blCyB/wDrCmFCATckl
QBGxTVsLdCLHRzsXtKGdHcxKd2YmSvydzi4BD5VI8bnCF4K7TQsibgVh48vTlJPcRH/6grp2Z8TP
EEx1fq4MXNiX3toXixmt4HIFyqQiEqhrIP9s9kRn6+oRaJBJmj9oMuS7YPTLabz8mq00jwtC0rwE
Wd53Gj2yGhFUzJy4SpO6Lb224IakyFQ3kejAuj2PjRGhfTIrby4QqLQoiQDc4cDOs44f8LhjvX3F
tCejfSRGKl70kr4kd/jEeZ7u9tluvH5rpzz/cq4CzWprCjDn9ALS3Q5uqqaWWp8aFqcW+o5SncAx
XSCC48+paj3npSiHlnBfPwI9MXFbL2P5AUVmd3h4ZTGXUlj/FFDSTu8QDU5XHLYYYKxD3BRa5Fgk
f08xInuDKg1KrJWeVL+WkV34t4PcZyKBlzMLx1m0sxmBDFTJvhr8GiBD6h2GUO8T931HvOSC1S3/
MVwXx/J/YEtKexIiN2AXrMBQbXVzubpYPzC5meYA5S1iXbAFBjl43bfpDFKAjSIaZ9ajBYAq/kY8
sfjcQnN5G3CDUrqZGp27ZyQ9xtYuXu6opbKoPQrCNDw2HGXON4F24FPDCzADqxIgCVmcpSEwuOis
cKsbZwPhnskuwq5CmPiQPjQDX9uoSM0YO9+kfgJVJx9+9jxOpXphUL0z5pXJ/a5cO/MHvzpndEvI
goRMr/6tzZDzAWYovnn5JTLuRorWseJMP2bmWdDzzHcEMUdWO5XvR6b2KnLAGTp8pD6jZl3LEWPI
r6g9wgeHQEv5CgPhYeNUgHENSdrS6hFH1lzCkRUTffj8iJkSfzhXuHMlF3jjT8RZhg2jhXBiJll0
q2hzBoOz00EM03Lh4DkVRtntN0uuEKsh9WBJQ/+sLwXNGUDZ1KBLAkPa/pzqdYAIy98UoNfyxFdq
jbo0SjikGYYNOK1vykjnFZnc3bGCFwsy7j/W+imvIouf9r1SqZ+WJ8jkOK0TKlvaPbT7NLKZJ8gq
t1XZjBLFuGlGwNGtCfiuysjeHxrnwOtdCPWi7CyD56D4JILiO1Wtc4Gk6epWFmELDxTdRb5NuFwu
Y9WZ+Irynsnxo6eEUuUksbqR2JebSBAWRnCuvfZ+wck+z5wxnXr1w/pA6wADCVUSzmoMET4mWPa6
cwZiICJGx6dEBYJ/IBOr8oTUpYcbzyux83jS+lWwiCEFdooeGx2vt/qD+/Sy26wHg/70F+5IgGlo
SZ/qvUbKYem8W//WDVHapwxnBitqwkEj8yw84NzQ4TLJ3xIs/CkgBSmbzv/SWf0uBMJN3pFDJFcU
X0EkP1sA3O+Eq943B1tXr7RfQ9Nzi24bLcdFJnTybDplDWmst1yahPcMC3LIgFGS4CFmqjNvURYm
sQ7nd7N0cyIfzor4COUgcNX/VPHQ8YmxvxfJX+1/z0ZskMGyntjaXnDnZKil3nYwNBVoM0W2Q6HT
YfH7quRGIaTEPl0aQE+ZQFz/lILtN9uaT5/hP7ZLiQnVPax0U9kPAEdDNSiRb2eQWpX0s2bHS5jM
CQpRSwtVKredpgPrWbdiurMwyLrXv/kVdS+JpqBcd2APRlZIuUsyBiMmMtZ8a5+cxlAJfNn42b2p
q3vHeT9MxI5slxC0/c/pupk3U3AGFBMqv7OQ4OPrWri3KyznfIkG0lnxBwjncufpudTdGdhiJE0r
EspA4cpWWAUze2XJXz/FHFtVe9+G/PpZlKYs9/e/SASJRGnWRqh8e3w9V1udi7gw+yg7zTR4VtJb
4BZE468Xtdwva2BwQCTMFzVr04ku2/4B5VAteVXQRpjbqH3a3LBuZheQ+evNjlODLXOGCmQl4Z+z
F4hgAbw3AU4HdBE8AJ2DzKBTaIxR3xA9bNoe84BgyiszIFOTnNA7BA0omQmtCLdgK7RapsTALsH3
/ZMnHW3i814pi3APPXmm6uQ1eCi3g7bLvkCcfTvljloNEFjjBqcm7UBjzfCUnVU1bui1ch1TFEc4
wFUUz2hrf829kULWCsyqGpdVnZRwR8bbV/b7qDsTimZ2gGEh/Yl7eOCat+9flIP1rm05rNlrfkuD
U84Siz6uD2Y/1f6n2HfC0fx/bqrhY6o2bJndDpSrfS5EoURc3Fyxas7XZWCHobEjr7jOPP8w8W4J
oa0GQWuj7l/urqbM1vO+SWlSYmWJbsG5Hefvggl4Ql133+0XiIEwYltxCHYt6yrHeD8UJQEMsf+1
LvwpGAoICY+0dgLOpMEKuZuSipHM/4wbQwcZOjyxMI6XX+SGkmM+A4pSFjfJQnyMUFXtYqUMmAG7
uXNoJGFjeWtQ9IuLPauzbTblWJ7oYAAvhLZTvyJMa07xKZuTT+hoJ+LUNyOuyXDjbmo7c8nNGtHx
0RCGDMvGxw1u5PPQzpBHdBip1K+KKoD45Z/YhNzeU0EWZTTLylVRW995z8VFHtPuptrTXMyU2RWm
2I8CClWTL3y8WR9Sjpxq1M/671A61GTI+Zt96hB3jjHv5bVy9xFJAeuUTqgO9EJx7FTtRV3VKEEj
SY2BFIPRYhe6zzYCZDyTjmpw0XNm+lzIqFbUPjasb2HJqU4PO5Yg3eW6fCh6ZsyW/iHj/rMW/ksT
w/ry8EzFCUhDT1SmPgLl4hJC/bBJBd2Yj6xGklnjHZ5GaPiFXnXZH9IAGA4OEsNzmHy+qcOeWx93
FTVKs2VIhEp4hRcrLF+/D/22uzLsK41GqT42n2Nnq/wcb9dxpsgftJmM/BUUHdNh23H0oDWw8kTJ
fgJWwH9iRwX4XUA1bSkdmojNVCMJx00MaZ3VxbnhR7Tyb6KKjBR36XxEVhoZPpoCEPWbU2DbnZg4
CF4lVR9HRzqSY7sPtol+wdgCVKD17LSEhseyAruVn1kErERtrc/3nyuIhDHHB6cfB1PLZM+Cc81X
xVlZN929HlReXiFHZ84+I8PBY2g/V1vHaQ+N16AWJcjYG5q2A5oci2kAiH7TtFDFeP2cV6Rut3EU
oE9hrVdMHpiZioGQu0UBq0/r8oebhec7qjV78VIqQhxbablNOloNAGuVaIG7VZb7tnSruAB8YkF1
kDt5DRug6AQuTzARLOF4XRDsqiAgO0+F+GdiGKNwAToB9xPBcO9idQv89CVvtMzQCO1Qcafkp3t2
2R0uiuAzgDld/3vM02YMzKViGPzPAA654dMiLgXDuA+GPLgiNCS1643Uxd/83wZOBAw06AjfgkMc
hw13M62I6xV3w0gB5FvKdgI9oGQakqlnwmDCas5Lucz90Xw39r2YxrRCW73GDMM/AR4fffzKC7wG
7M49cpsx3mM1DtEyzdVLqzU2e5XkufLpmA09ynQT84t2kvcKcsrwF+J4Ej90ZM9B4iQ7WsDWIHAO
5KAvGuX8sFsBn7BavV08yb8n287xPXspwsXNe7o+Gb4tV6kUewakp1hm3ECgWrtftWFzR46140ia
jRmv8HyrsPNuYBZ7NsnMhX7FCYAWonO5L/cLa1cFRqX3V2eAQUbAk+Mrvx6daG0ypw31s1fxocg/
HmENkadb4HRKOH42abVQTeJcSPsI9OhGx9IKKqqBECM0n5eGeUDP6SqdwtlQClr3UuHstREMl5fo
bVyb5qbs1idPpEFSa9CPkckP5hUb+KyNVNls6V/2B86KPeCJVq1heArHfx47UPg0lwcdqHIcvMh0
SaR46rV7R7w5IeQvCO+C1dRd1YsnmG3Tk/1wpPcUxF0Rr3NjmykmK45Qn4UAq93up/HMMSjjd7cl
fjXtb9gaQfC9St/+8rjznRbAn4EUT1VrfDI4OpEshHXqQVPN9jTVe4WitLKc+ZfR4ivvIhFTdVEc
PBl9rjNP+daijIiXA7NDnp/1dXiRBvogZ9QQbvEhL9PSUWvoyTpfj1aMqsLZn0LV0Pei3zVqZvXc
lGJpJsb3Uc/1NnmQiNLoizU6hOHS/OFipbFPHwP5asvHZaRX7/60fG6OVkI2KzJujcgSyOZHkFT+
6Fwu5xTOvRq/SeVoS3l1bDsfjsd0pXMV3nVuM6IiVB7yg4qi0iegp/8D1HyMtRV6pmeERG7iCDe7
PmDKBZ8em/KYdZ8WNFLAkgSMj3IhDKbS2zki6hOiRS1mMTSeP+aMfLcqU7eaHbu/iV7KJyGGNqcz
tX7O+8j3vsVvKrSVBdm9/8609qKnW5FrwKSY9I3SqdWptkpM5XOC3fVjo8y0A/zD8xQLTv0g4/IX
dtU9wKTIod3wvBctfQXk4135/m1bcOfaRxBxED6vG6529IDystCL8BaSZIekQagvpYNOl1G3KD9s
zxZdunAifuRfGq2fCwmY+6IiSJgNI2HpuZW2wnh7yzp+g6/JS/OqkFM7kHB+q3tmn1xXodnSXj34
a/0rThVsee55+nxnQKlgREROF6Y89UOpp3eyEdVNNfnAZswnP21L6aBDGViK4x2qhX/DjVGmwRg2
D5N6mKlEm22zqPcoviHzoy2qqMnU4vaogo3cgr22RaLnlHrF07csLe4jktQW4Ixpyqa6E/alPgb7
e+WSiKrIbBnP+SV3Fa7V0lUPjkcpyRg4ZhL3T2T25Vbe+hwQ10pVFyQPLuPYZM27pqNUKape0GEo
g71wGEJUsahkxtFogGAlr/a0rRFvshwxv5ekC/RVgUyGypGcgEEG0PFRmzuRJSiLa7rCch5ts/3k
0gLeJGIxb0hmrda/nQ41CYo7s5x294u9zWgd6UViHHB9ry5wq42nSvX/oub1zmR1ne/e6blKA64t
BCS/T6ZVvFKW6IBXoLaCRTBcitYfjTcGsTgiVOcZYEpaA0tTn7aIjbC9bKOia43MZsYvB4PCv3sg
2lOmDxvUWpzQOMnwkXZ4lN6hOr01rhthfkKDn01R+bnI+iqkFMCksz7pdlV7X4qFuluy4j9Hvcfl
cEG1Op6xdS/5vpER6Klv6p1vwrW4lA4zxAOlfXnhWCTMcwgsvMT2jNol2292V1G2pTedb7WqC6JP
K/+R4fKqJjEJi5gmGWtf78zFQ0TAiYEG1LCh/A9mfEo5TgUB7uI27MuHWzRkeN290cPyBjaHRqkb
thJWStezljF8GsvNxNjklxTLhXlTRtl9DXdZoqzoHdLGgadp2JHIwyKG6nLqnt3fVq4ySNF43L6D
hkcfJw83CM9xwwsjZjYDSOcVmRmqO5dGE9+qsuPCCTYpHUAcEQOWf5PBcKUZS8AyLus7/GOtm73S
4YUoUnMYHwI52adgXrXC+ROzGnlVDFgNp8eWvdBu8sT5Vvspb8aotzd1rc7nQ1gJ3v+lMlEUObsH
UMCV17GQS1kiizwKhnVygk4c3nZxW3zpzt81nS3VXE27nv48vHlzVEylKr/Oy+9F53pOIA+BxHeJ
PfTPRr5JZ+8bGaySZs+DLYDKouvSfjumQYBpPdARZF8KEKejNpJ40RQgdo8zUy3q3ycqLz3IwdP/
1QXDmfo1S4PKYFpryBY1aD/iZabhrijj4In5ngZtpc6YnFVeRp1Y0TPJ3YJxK4kgKzTDH+vLQNi3
lwD6l+RMXh/3MQ8o24ncCQKd7uEWoB6uPzo/6JecQpYyfxJJdI7PMP1oXnqYyJlofVPiJY8tVTX1
ySV4dTGKhoe2B4Mh3JdCqo4laS/0u0UPx4gyIMZtIsd0sZR93AU77ho8eppd3kHmGN0d3y85CPVC
ZulUWDtCvo1Nn09kPDIDOdXYJcz83I7mygVof3BW7ZebptJe1P0xhiszf6iJAUfBF3BRWRskuiLr
qyteygP8zxtohxH6kJuc/Vavwq5VFRwFo2YKAEHh70+2jvaQRG8vK9NGnBkidO02JpQRurPpFQVK
zgqgspU21nSYk3KB2SviroDdoXK0+BBep8rmruZuwZiVirgrKHnxDJAjmh5FjSWyqWdj0WuGaS6Y
jYNN85Xq5aZv1q3PflMKe3oAfOfIfgqjH8QCDrX5I7orSfvNDdnN62Nfz8falUmSK3e0sqCknPN4
6wdVpd7oNDLFJbeX+uqFH3j4XcfT/k1M0c0R7A1TXMwH/mzlMNA/vdzGw5obDQvNlkJLlY4bcK5e
R7S7Ugbx7+odE/Jsws5sXu9pLo87DtMXs6r80BlBwqHo39+CPbKLcFymLO3ze/7ghw32agDcgPp5
cRFNoKt0hAd3dz8kNI4CBCLuZiVXXjxBu0c0Mcbmcjz4nY9ryCUA/L1Cl04Ws/sPs8k+UhZMGLLj
hOHaTVtBmT7q7mWf4RtNFu0vVfw//Eu28KVz5FeGpq39lYW+F5rR6HkO0nlZYya5h9EaUMaqaA3z
Ki4UCpXWZsyYJYVT0/KeB16qF2VfPuUxX9ZlfAB2w1r512pQiZbkxNvHJg0L+m28voHIXuflGL48
/YMnSi484t92N9oZNRMlQL+Ugs9sol0WFQXc7F2De1G9+OgJ2mMMIhIW9yRfxtVWINEg430baITo
ZwCfzLod68SRux51P5Da09DL0AgBWKutKAa2pEWQUehJk7DKpBBpejmyUdQke4gipiEh8B11z/8y
tIuUG/ppsJKsoo+CKN8YK8QXf8EzuclW3FCgtxlxHgtsZ/D08gj7xlUdNdAM39PkewaAkX/TqM+d
rHqqNagcr8aX5Dwld9CULRjLnE4hWVs5O6FjuI0xRTyJDqbdNs08IGWnf59/kiPUhbX+wdmy0Uc7
2bUn12sIaEJO4J173pBBfVu0ObCKgcDwF4DzkRj/SEtz3vbzXe+uFzFLsvllxJOBDTYkFXYOk1Oo
CFpQQnh5BMorJ9YhGp7lOs7A/GJVVWU8Y9EnAdDnhLHNz93rHncq5vQYOS85Clv420w0DXUT/4/p
GE/H0JFt4r1dw+ncLo3btuoG1nYPWAbWHqgfQ6i5XNlmYvThXlrKzYge14u8ICD1d88Ub5KlqGgB
b5fTggZrFFd7gstJGk17BbDLHubBSBqRWw5Kb0NwrT9v030waNzU6nkXqHX6BwPnkHsdrO7OTNHn
l2Qb+LsRHQBy3Dt0gll8xMC7kIwjejp0FGIUvcJ3tK3Z/rrG1+jiUK8gkU/MCMxzn18MLzmHl5Ng
PEuzGHoZMhSaVyc3mxI5Ektcb7pQ+4NG6B7e/RJlA4dnF2gqIivD7tkZy45UW0hv/Z38k9sC8N2c
TkG2dGFHZE5MZsK2vVzf+uEdKPgkg3VHbtTgSZL3C3k0U0SbGZDsQrCu04vQ9CkeAKaB518Lx1fJ
jCPvdjVho355HHTGq1dkv06B4IeGWGoEczCqGMPFLPmWN+OoELjhHTSpAi1o1jSxvtVAd9vMV0gB
XTWJd/HbI77N+/pkg0kUKfaC1AUVgCuqmKeNjnUuYNgoGedI1VWoFtTtOOhA2ByCzWQcQQJGoALS
r6O5wHZcLbenfJLdpIy8bq2Pxp8taJ4CJt16NNF+nr6tnQSg0y2WskuccFTvl0IhbmYyjYpsW9V2
F6bEgTWTvfPi9qsJBOMxZx8CKstq6yv9jUKwSFtNQvlRPCjZAjqG7Uq5051PUqmOHC+nM8tMNi6l
CygcH74B1s2SHvtgP/pgJqOXs9OWIIFSJPdkfqQaRS+OCHxBsik0m+9jhCAkJbXrCSbOPYHBrsrw
jnp8Gf1fM8e5wOIg7HpatGpYz8rL4yIixnaKhsEYUnZ2k9HCs5mKlhIlk/wYAyN6GUB0T0yfh4Fp
Zbn164XbKL7TzNAnDcDPFMOGDDL+/B/nzuphorpdoCn/0I/Bt06nD8uvH2J8ZdFZ3webfa0xqTmM
/KOdaZxR/jmQElZi45X5A44qg51yPH0yfh+6anzf2K0HcQ9LBxgLK6fWm3bwv+ZbsO/NyZ502jWF
X0gqYkYgO1064dRtXGbADvw41XF0VCmOCre34S+01J9T7c9bVdQSysM4Rc7lSRLgAmLvxoSlez6z
HGyb42pFJ36XqiBPqbWcujDCU+VWukpyzBfvSPomsIZ7kbNhAvFa1cTg0RQN27md0SRQixeP6/eE
j2b/JZk1SA2MkiMxIVLFwcPxef9QyaWBnxJ2E/DIWRdaKgMmnKHwYYZbPD71FrkSKm25QJ9rvbfK
xMuBH/HMmN8H1j086v0ADeNc2WPkXQLZR+uOUVH6ywpoCnR9kyjScTPbQxhkTnrI0HDmAzWE5Tm5
vAZTMtWSjgOhDKNV+5xy4xJ1CpyoN22U/e0s+r9ERWs0OAzjqGRZ1wZjEEPScIulaE6938qI1CX/
WT8BR8K6Y3kibGpcJFBTWH7pyWU/tXlqQ0GkqlD/8wNcMsfPYdY2PAF8LzyClHPmlj09XbO2Looq
pXann+H/TwSgRnTs7w/IPHdOEaEWlO+QfBiZSy5bJoAqQodgwnbM1Z9saPTGRWRvlJxBKJX1msZS
r+I93EeXSXT8zaoj6U2FYEne5gXnQOUk9g+AXabnzeVBl2JQcM7mQp4SW/DK4qdQD3FqRBWq+iGh
t/BsTpyHOcjfSZ25NaZ1f0tc96VDZcN7uURZZrYUybF9gBSUf8Avi+7UPKthtIcvdcso2DQMoo7l
9RLdHJEr4FkpRMKmbWA1h6A8tTHlkNPfg9K1d85rZNuG6TbOzArM+oIddQCqvNgYWtiTZiRVWIcy
2SQUlQ5LjBY1EuNINZKRqZLP58aYdoVGiT1KK5cunBR/5s5O9XOpJmkIKjil/0A3nqW0qOUnAo8T
VnXuSO3FNqxtPMe5x71PcvmyM6uSU5yhfygqEqEhQ8d6vhexYNdKphcESgZfHak/dqx6UjwvSdsx
m4w5nwPKmplU5d7QcZM+CRL77FFw6/Alw/tEDh1KIgqW9Ig3ZQhQGpgphnpIRpIOB6fMLIp6nusC
POOShCkmMNVIcqEV3coAM1WzomlS9RUzkSTX+fUMwgcTnhKOB9L5oHBYSODkAq5tPTs1NZ5yitpb
hPIHlu6Wm1SZCeRRWHMAD5xViTkwVZdXRoE/A/HoTdrLE0v8FN17kH0RxZkjpf7I/SujBcN4tnSJ
OPvNeN0LwDSHw/Hlof9u52dIPJCFmOh4ZEKyv2rUxecjh7zmCH4oKqXv7FGkofkytwbS5+VIy/EC
P72X7tpXJkgceKwrKRhcKeL1za1CHf3c6j1oQQfe5Uqo1mYUA/FNqp+8e8eUCRBKlAwT2PskC/2A
mDcZ46t9FLLG/2VZeqpFTkQIUkC6BkB8LcodvQc3S0vlouLVsVYgzIeV41Mf56AZ7Si71OVnh/4I
NyumwjUNU/UN2WC+ZQHqXi4jDWG5vFTUhqrff+vHgx34iSyJmn3bR24yMD1a7aZGqbgTE0QF7VFC
Q7Y+UpW3Uy2PNwQGOLL8eISEyjBaQX0kmrgFOj1U30SFYCGFSaxfMfmRZfqtwDEHddJsWms0DXJ8
voVnV83aRofuoSwqfN/ZhG1n3nW3em5t60YEYpwktW6t2xF0rQWF/tkhMY4rOo12vMIrpx7Kpz+e
zruaHu4YiLpFd+vHnpislJ3ylvOoD2OHazYuIts817HXB3lqMuZLUSDlGEsnT3vH9D/bzvMbAYvu
bRcGTYxKY1eVrXQlL062X+j7nvfJCbv+tA1JjFNhfMgKIG9lMCbonccThmiMOlDqRzdC8CLmMBdo
9ZfoJfBKvH/Y9z8ajSsNjsR7M2qJHq8aANx05EmVWSxWnzRnn6FemQswU4I4PqFiw15/CpmBRUVG
1BW0TEwkO52NO3VX7iNvcceS0LkZoMq4P37uXI6sjGF03g3jI58envgwY1t/6t8sZeS/zrWqgUBw
OT1YqJgOoMbczPQbVH4r9V9WkqnwPbMWFqoARPeB+6gur/v9oz6tcHpl7Yd8KeDrYw00IS4/PRck
ClS5jTEPCTTKRZnRsJienNMExLCDaarS4UJ7WYErjaUo0aSp+LYVQv3v7lgQAf09BSePP8FPcSM9
SaYyqGok67mUDVu2fKDnikLqEAFXsFi0BlQawycrgUbF1g3imC5WvRM6v9njhzRpU1OVvEniL4yu
LGaQV8fO7ZOGbwYOe8TDO1DWvLeJhVMmCG7S9ygEzhQzx3RIUsc1wQql6uf+xAr//pW40slA3Pgy
K+cQCa2SyPNaH02GZ8bP8ue3POX+le67HmSPBPAHs/yxIiaSi4KxYmXavJyz0YaLdnMFPPdFpz1a
3Vzi0MqcCkPirD1/TC5MNvkXl5tdiJsumI5MH/d6uRiQ5QmRlTaCopeZ3olZjJNpMuqzHxeIKXEe
O33I56/WDKSEv3NFu5d6CA741YXLmeDUJC9gx2D3STML89c8JiA4BSPYnATIyNNsaGsx7lHYuL7q
BNeLhcmbYs52mjTACHKg4b9hLhJ0w5u8+7RExTgtnIXK1j+2vj90EAPE3uePZSx8iZM/9ULrEfbl
3iXYFbt5ray6t3oORNvnp9o/DZEuSFpVpYFyP1v+w6jxokcgoJLXWR8MIMZuBLXsloW5SwPYiEe9
f93PHNLh3Mb0IDSeE2U/erDCsb6vSbJoe9o+JKhSI76TMk2BWzvYakykldZh5v4ehOJIHBKOLPQU
GFnci0NY8tKyTHN4HlJD18qA9ADvoNoPX3y40C/LC1qhG+kj2nYQkI8ftv3Krq0uhPHHXGjOSRll
KN5upKdopdnWIHYUuY1PzhW1gFYZ8wKSXGfH7mQO+OZhTO1Rm95R8CgpIPCNLB7Gs6n+r/AvkoLu
5QokZyE2SLUGzqeCCbyl4gATkWUjDtXEuKqrAw3y7gUGR9UUflCG5ei0BBP2/e2OTWCrNXVaFqlo
Ax7V6qqEDyY+XqTPEHClMsWWFuTpfEf6HQX56DxQglRM0Y8RF3Z8+VB9uwum1XSDHzd25gpGy2/N
lMtgIbA3Y0O1fEHLw/c6eyTGpu+EkkrMQDGLiDmyIgVlhWijAtq9r+JiO72SAD8AdIEDitynYFlO
lxV4yDZz/bQSBhlHJrSrcDQck+/pk4EyXGGGdp5LqvgiWsDHkZpNCyQT08lk3K8FzN3DehSNmSht
q4z3pFbQ31SI1gQ7x7BIR6VLhzLEmhSx7bjU1XEAx0PDxDL+x//EcU8WZIjqhVjGtpwQeCJrbuvw
g8Ay8DJUvx7PwSnFaXzeOP0xXUUVyVtdpXSwj/ZwDj/Xq9S5xiihbrUTyOjMROKyQdG4OP9ksXJZ
4WOitaT4Mp4GT8Eq07C/SQBuPjpAlq9ytscJQ02uNi2nvh2stVMCjqQ8j6N9imA2rUeF+oNhLt8E
xhfERBBEYSVPv+kykCbn8iLJ7heDR4ZQs8WQYFeusYDl3S2ypjH/0a+WHCKtWsgQUqwGBYOtPVKO
pNct9bv+rR11ndJbZrwHocVIlzT0h7ivtoLHmiV0JnPaI+ihuRWRx4O0r0TpBECjo+v5YaZGk9c8
M7166e4ePpBD0TyQ1LqvzAJM8eY26wOuzqDqOvTOx8+Alu2IlLPF+auBDbx6f6W0Yznb8+j9ESUw
TGvMtBxK8isWLi3aAOvp4M6jIlXFbCJLaC8gzuYV4gqWhVgHJORKAYTyXhNL/ru9AjmSMgQ14xLa
/7HtHN4nPg0n5lLwB9BcobgIthjATivc7L27uo8FkL6S2/kYFZXcdRfJ7nJTTutA2+mofVzBrJw9
QVtedIv0alUXwAbFWK9PMxSPMIqQ3p6fp1oWNBhoULqjkiym41uJutQMrJvgPMQaD3vXrhXK0N+Z
Z390RjhRe+uqxMQaxLGBFkQCqvoASAJ+XlqvcpwYZdB5H4wwFA9vE0muk6Y/VgAi+kX+2rIaIuFB
D5yAZjpSxZIlP4uiMM2h9xgAcZuhfbNNBDZv1l14P5EAELQ4QO9WOg9b8djpX0e+SZQc/qSx8+L6
ULUaa5l+ZDbEcR6qsu/gJbveoU32FypfJcsCTXM0N4sfeBVoL6ziI1ShngK1YpIwhHJFRrXWJTOE
0jY0re9Gv0qkIdsSKoGn1e88UMDqJJQuZ13xZ06ZN1Xz4isaFGK9r8SQ9Qv4iTPWsAx5b6InDi/t
npL53mz1xvlGD9bBa7jBQ9yQc2LBUPbTJz/G/HlQqkKlnIHUH/LigQf2M6n/hmOD7Htj2j5zF/ef
adRHuanGHptel/1sOhtAiIDY9anQ9QJub/sGz/8M49UdFpvdw9bb/GeLBIJYQMHYGBOTomezfHQp
/jyRbitoWgjBTqnW8EGsSV1tIiURRu7+cc6Jdqm6Oqps6/9a6TSeU2FgLiH7+d+PUYHKFaqGi60l
DW743N870/G+EAez+GtwX9il5uoU/DRpepmuS57nhv0iM1dgbS+W+lDbevtT+Oi2hTzVMStmua1a
uKztCqhDh0IE8GAn1ohhCNQ1U9FfSqlZoFb0yzPN1n+8v/JnmcMS71QH0qU3jKqCoHnvW2uAwGFu
g0ehfox9X8N2iwbNbkC5I4BLnwdrS0nsdJT3KAdz4UCHRqmoqNpoTfDbEhoWK2XWpLRYCsWfD4+1
bg2Ge36ZnymJuupOMiCaMbeJEeryoCkwei5cSEwRZpq34L6hFiVCrSOpn/D7ATnB8yjgm9zQ9BCp
ozmJEli545rOvGcM7bRJc/c148fkm1ZOW2ZbC0nBMvmsLlhCLTmnqUQ3P5KmlmkpfiVjWtkjZxcx
r8QlPujf/5OAVW6G/y7UCCD5HSFj/HyU/KPe2A3oIAHCzylP84G8Pb5IjZXlA83NWk5o0S3GubBX
TM7QPWLyNMkmzY0SGx8G4UP5ZLZKEZph/HPTN3pG2mLXZaFe24e79uHGVy6HAuOa7XnFAJUJMK5r
dQdxbeLErjaf7SLmS68O2cvheAaVMCcjGym5Pi5EqCtdIOCarnr4QyKKI03tNq3nV9J+ijA7rlEg
z33wrloK2lvRldUzqytJi6BJPGUvJyDTmYDVNttPekU/s5sXUBBqzMyoV560VdSU+t4h7Fw54/HH
J8At8UUlUO8nZzd26kHqftUNO/GumQzS8MuvzBIM+ayDOX2tMb5gb+eCLFaGajNmutMxGt0AG/6s
kDxR26kg7g7uA4Nj3TjaRGdTg5FixK5JwROYTjNOoHMMLtIHrk9fU/M2cNh1HEWHEJyOiDySn8OG
vbblwh/T/ya/uUOoMP/ebYBgafUB8n6O+c+88FPNtq9Woa1urU0nec2VHaOcB9E2W+dzGHg0ZoFJ
8GN/c3RaYoT+ycpgO7guL3nB8ZxFST1SHeWEId9OAXo8zU/dPPlGGeTSRbpaYSpMvvSigiPS17L3
WfQ2D2Y/UHUMSri1ILZY0v5sDVJIsmlewrnhvwDPPs1zQSbBBAiCVFBTd7u1K5PB2gjJ1wcYiK18
qCzLAJJmsFav1l8e1Ua3FxyyyYsshjvVseoYXHiLw1oojsq9t066JSQpREN2VJ5aeu4wdXm/BT92
SyrAYQXv3w9laeHFMOQ5WmMqPtXcoVyoq4ZlCn7tdkcSaWB0BfXvkRVFg9DsQsoxJD4dlFL8fAo2
5lRl2HYfn1C5r3JM0Yz1Te3PdAYwszJUmJhUAHv0ZxuUCRE7U+9OBOdNGSF4OQ06hnQvK+SBbuP1
qMx9EJjKDNAqPLQ9uvo/wn9uz759eAYCC8tAPHKjuUvt1obEAZlEqAd1Yiz8jVyt+37SFl0m5Yln
MD2nVMotCBMb9fQ2hH5SMCZKKqpqy6lAi34ecvt0Yc82q9HKuh/eFui4ie7RikY4+AoM/B1E7uog
s55vm0TtMb7I1B+SN1Hh9k9eOJDlZ0hM3no+5S4HCfso2Rgup3Ex8CtqQq+f4gImHljcKLXlskLW
W77ZhMcqF6ePViE3LWNBhiCsVrE3DsLtC6MfZlYk1WJsireSRcpgnauBsnN1I+FZRFdTYNCwh5S6
APH7TU0woWnN2dYMcl/0er0XiSfl4XveQzHdA7X59h36u7Kgr9xH/ZkuCfkaEbjHLRpp6OePqPh8
1lbdHAYu3AKobG+goZBE4FQtiJUSar+5rA61SH+yFUJCjZXybJ+jhYZ/8rX73N7Bai2X17d/zzc8
33iuUYN5J29doERQkZXR8Q1T5fJTX3aHey/g4EDTCxaqgg3tFkxJq9wQ6QsxvM9wSPit1ipmoWzS
Hhz11jbhInKFIwsuTMNLTpONVQGiSB8iWxPhE3DuXD+n+etw6BZF8BowouASmgkPALexnIO3hbJx
Zc81hyD+d659wKRHKygseoA4O0QnGtM7GB7Di6gdiEOVeDyo5Z7pIsVZYTwOZ5hR0sl60+W5Qwt3
vEOIkFnObUuL5jlkQcrI95Qw0Y2+8O3yI6NuJsJwUvKxQ/dx8p2iBokFJfocOtftOaHNy7pSsBQR
yFHDLpS1x1in5OGWeDXGf85siJ56aQRt1dL/q0hy7wuXV8ZqjPNdJBrEBllJ+Z60wOb8HfCCGZbw
KKbby+Tkx0HcAZn/fHKHACJFTAKGt7J8fC1QViAZ8unh4QUxgIAmFG4djZDkgSXlmfF2oc0LfUZG
4TGWASM/uWnJ08zloQ7C51fI0q9HwRnqMaY+R4wes1udx070eVpgJhTfwbdbVAneQ1Zat6CKCoMG
8HScLv3fGq3RNGqPveNqACAPaZpgAPgK9ZxVmD13ucJ4KLwJof/M74xjphV2mhZ2V1HJ/XfhAAqi
pITVneMat8vTZMCzZ+FGvkil2Nx4v6pUmtCOy2Ycd6G6AGWPbtYa5G8/41qhvs56vPTau1nldWBu
W+5hfrSZRvEKSrmK8Odkc4tDV3qBAJrbs4zeKtDFfkY7Lqw5oTzKWNLnH8xdosnjgACClLjmMpVE
1eQ9cNp0CtI2arTBAGRlZAYaLiw8680gLBCfN2DpVzfyNXCu/jQKtMWm/FBZp6EB5Cf4fb3dxVJC
JrUqQo1LvkvHhicqWFHZe6Ij5ylHj+WRC79FfctnfUvF1S+DWt9we/Rjni31woRnMdI7hO1t1YpA
s3e2wy3UArdiyID6pUMnoFaTddghxy02sQlPjTOyhkOXMqw6gpXfVgK5DZOWV/vr/RgeFRxD3t1k
gdkWAtIHPfdUvyoCjh9hQ3F8sXOQSSxw8ULV1MU3ZAKz4wgU7wBdDhVxdggLvfZKLYl6ptAcY011
+5+sClWnbGMFFwfzq//ZpxHXekWHXikQ1bbaDiEjyLlQYZbupnnBfa5e9Y0D1danAEWVQqBknY8m
3DHks6vUdz5IWOIafefNQXv3hL9Lx0M/BAqaGfSB+NYldcwm2saRVEa8SIdFMAh8L6codVlJnXII
0YMuXuw8VfCVEx6Ege8oAWtzXxRnJxNjTwn1Amyjl5eq58TcVKVPvtzB25uE4WEXbD+5zk5mqVVW
hV46L0+U2cv5a87w+LD4GtQINK9tryWPQy28pT1KK/9336OCV/Xdi77a+mijwm7KnJP5W0pANv2H
/cGPqaOF7cs8BFatZ0DMpoXZE9/Dzw8AecQJzTjQyZqH1/4UpDH27SfoIdwzht1bsU8LKmg4owpy
zK5d2s+/019ETTWdUMI4z7PMsrjx/o6CXgARPNxT5AnBt4ztZKTuTjV52T0CSxFbMmUVvj9OiuFo
y29Q309UP7bStQcFA8lmOfimsJJlff27FPYv4e17IW8BsLAb/LZ/pTbri8UDm3mgK3FHrEyufY/y
tG2J6SIWgJIdYBodwSjAtleYoiNl9NrmLYQqkNCZHXXB6UwkrZt2p9Y2m8eRDtaHMIMEhJjwigjv
3mr1U9HTsc3KKvzMjwQGIe0wePrvKvAEoMwIiEuBGU7bkNq8rrnp8VIO/b4yaFlYq9xTpFj9S9Xb
OLvpTd49QXEEX2t1RfLYEmcEOiTG/C3MzpMTLupGtccmkG0e+gLiJEFM9BChYtxQ2IfAcJda1Ns3
TdNL5fV5kQwxjRMXpkkOVjlSQET/wjkbTXgs9zNTd8rONHNRAmEh2EdiY7VG8VZHtGiQ9gQDldyK
npQY11QgvDxgQa7uyL1Iz5hDw5Klq66EWeQD0ORg7TEdh1n8qqUwM2k3OEF7XAQXEgESY7DrY82H
OM9Zk1g6mav0l3m1wR9oK/WNfJqOqBOr/UP57ooVveBHMsYuCCJK9Btzd5Sr7bBtx2USd0jP+MXp
UmXIY3EqIUAaa2aFpdZWuGqhEneSKo6UJQ6EWnUjkkZlu13LU9rrlDOTaQD2/WjlALe88gD1XdZ4
mqQ7nBulraK8a8Uzxsi692b4AENj4t2ptGXSGul0KZKadFc7enuJLy6Dbpv2Jx/fc3naxGYriJf0
vh/tez8bnW2LurnGcduVeQgDHNMUN5Z/Y5GYpeBIDKGo0JTb3CNXRR177IdzfOJhqS5n5T4wg0qG
u1vOOH7piLf1/H7DDrSumLUwFP+rOOd86tAw96usrfgbRrIyqezoSVK8TLeewhNVKv/J592a2d8n
EYfqdTygi7L0nVV8IczHiHr2vdS3TSiWQvdwHoezRDFZffoNMONyw77dAHoTDMzVeVxNzPJxfm7o
ytpxMkZJFQ0PRR8xFmK44fG43ROxPqTwKhxLTrajCoxHR1b88c8Ne0Nn9o2a5sff8vb0BtcYYrt9
UtXnvYacrtk9GlHawdcUZJzZn/EEGxx6M2gCdSUzwASiO2eC3JFaRkNLeLjPBoE1Q9fLW0kPnf/q
+y/178zLqpcf3rinKE3aYKFsKvu3tJVFCnglNhqNsQ3lLoCARvHxyVpN4YTkay/qyE38KqwP/AeA
AXNQ94BYyicZ6v3r0lIPHUs0HVnBz0AmdOqZKYXn9fhh6FnoQtjdWh+sV86ERMIM4Cb6wVrFtTqG
3uEtg67HYQyuRsj7MQfck4ecY6tqdGN2IhFfRDCgpxPeZAsoyJYPgHdoVA8KHvtfhE1YYULbduAF
9PpaZCeGK9eQuxJAZx5GspLfOCMShz7TV6IFkIgrgH4zhhGJOhLcFuRjqsH5MUVuTXZNdvPPfz52
eGfElMIkhoI1b/ahPAXd0qbD80epzU3404LrQZEzO96Do7AQDFBnT2xk7eoJia6pUUNL8AQtQBKW
9dEdtXR82z78L5H9YV/lmH6BjbdxzuesTmTJfxghUhA0K32dwPYMyOgYJb4flzaT+PCfHApH4Yx5
5uBmlFvxloxp49gUWOnK7OKyrr8aMDtpUDjpwnlSXb46IfhryrUB/buE3WFW/om7zGtlLdTlJcPS
+Sl8+ILJLfpUP6oOI7OxZN6fp66GcCaXHiSygrfLelCFLab0JhImvgmoRMkH9NBJDmgQYzfgBH2P
IB6pKJS1eoZfbJkjsFqKk+or2WtfHzcGOv409n2DP1xPBHt7BtE5/LVXU/s+plR5UEEwP7FHPLXl
ehcDEoYe6SKE6KTla3IhRPp3ijOpoctdF0CJntHJ+RydtRuj5XPU5v6NNgCVTwsQS/rkWf8uWHA/
5DTYYb98i+5730EJEiI+dU7ieAOWTlP/ldAaeJM32eFeJkqYqeEk8pAQ05Zn0w7MKrJ62iawpTFq
QM5qcgPtLcv35oYyJ46WAZczSzJMakXW94FRj4DygpsbIpV9nSmo6YsxBZf4Iwq2JPkIXx97OwVl
Wb4T9HXHVAJSQdrjM5YHsuv+DTlaYAuoczx4X1H573syEGuLME7mn1MfaNEyxU1nMco4kuBMXQ+N
uF7SgVCRvwHDG0vfu4CeTa2/UH2wULlzg/QVpRhwxKvXZqhlyI9egDITpzFgjqvu4YctNes3oszI
Kz4McFsfL5iPUZr5FUEp4j8bbWTTM36yjXn+KEasUaBmaW/2U/q4XwudT4wIZrFVGj7qDyxdGADH
HFE3QY2BbScAiIWngFR6WXqcQgf6AFEToM3vDlGZmUvTO1jQZ12Io3SUV9z9TGHyWw0+2NZPQagi
+V0RdJcdoux0jPFfk3XQ6dzPVF4VxGMT80OO7Q6uzbUIpeWPZWxTsI7DFnES+9TreJGo2POon8l/
sE8EXY9JkwbnCGrQqFke58B9MTAnsmvc5pMaEnYeXsQNxR4oPtVe9+6qLFZnSjZtEqEETH5YCcqn
KOQ7+C4l9WVfIy6Ofbkd1eh8D8g9kaKep3UVmduRMYRwSjNWVSGP1HqPNJfAN8BLszK8LJP2XKtC
UuJ0f8GH7KXsveWmmvavcpkCRb7xR8tee6bZKM6Muf8dNOqNhGq45MKUfRpz2wgVd95bCMhntOMR
imummL+1GpfuBWQUU8XA37WVrS++MQfqKr3aex6V2VgGIs7o13b9K1UL7QxxcllQUFTOVgpDqL6Z
bNvIVYPqXxlfUPqhDuACGCmSsHJsSOZSp21LOZLCtedxMJsUIgfxa3Wk/4YtaSIt2+ws/LZkATBh
OAP4ky6RNVryLDnmnzVNoBcP8EAH/i66Fl01dO/IwEAAse9iyzwdtcCIjNex8+tEsi9khzvguifl
VtRFOpR5LV223GSikMRqF5mx8VWJepShAASIHbly6/qSEGI7MzqU1sud5gmfls0mkGjL8xHZqH7v
2+aEG5CtTpOKHZg6YuMbbw2Lo7Wjpsd1+zymQEZohLnz3Wo1AMmNdpQgaWnFfyG4gGr76DeqooY1
/H3Om7WSk4pkvrD8WBclj45TNmT8kim8Z/CSwFmDupoj+bPFJEaZGMMBOCdyeGJghQ2QyjV6qVAt
zKNkk79lzR4h7FbX9VoPUQEWBII4apnyDubUOoHEj5hoz5jDqL3GPYrOTxn6vUXIgpNVe9lhASZe
/Uo4N83GCkROAeWgglzed77rGCHC0LHH0PUtO3VTCvuLUTPiq93ZB8FZWN6urYjangZUjHs9/fk/
O+bc0tFH6ZA5VI++OIf8hNX0qdUSeAU/mTzjIXf3aeRUhurUUsI6DLtAh06tHvZHjZ/G+KuKrKEP
wbtbfuQcrwZxWU7SCz+9WQF42PeuBR+SP2bbCnby9lJue9u4IT86rd4aLSbnuTpkei+Z+r8KMUeI
JoR4uC6SOwwZoTudg8ogttEA3ToqQGlU0Mxe38yRVR+XaU3Syf+qUEIraZNKqc+Hyoh7fmrpRze6
iXJEbq+6TS/BRrN8fDEJ2pYYgRib3cA4Iqrzs70wq/x2BhqyDoly1bZmCINBasDXEPZhmCpOT4ml
/B7Htuo51i/3YkwW66lgF2CvDhKnH76jKzR411Oz1YH5IH9xVya5kKHQmKImSKDXg3HSCrSfONfh
Mso7mGB7nBZIOD1DZ7dXIbgehgxSuTQeWlCog9XL0emgIB2IW14wwOVZtOC+7X4gJBt7OtraACHq
z/FTq6YShu4zBskCg4uXKnNDQ9s/qw+K/FgVl8jF5QfQ0tVzbcMPFiSFlE2voFt7nrB1m3ShjNX2
CfXA3SGf9LsVnF6Iq+dDunnQLxFSVy+Ii/RXwO2b3NwRKAbPGYGOPKY9sgf1tvHumizEvn+czuHb
R9JFKk0cQBxyWxLXHQtfZyRE9j7C77iWac+uoojza7o9N1lWZxWVnWTO4hpH+GKXT4xsF2XAGYCL
dmy7RmHfnl3yGtzsO0j7BGGrwxybuwYGnANOjz9Q4jFukA2P9jMlZQoRHgkxTz+q9EKT9X2PB5sM
9zTyy+DBNkElaIRIClG1LhbnPaVWV6ldBvyJEH3dYyQ/3eb/+x504eVMAExwiMbbKV66vwPZlX0l
0jQEAOwxlP5bBBv/MXjp912PpP+v+GyQuizZLgmoxQslpkDOAV+VcvW4sUutt3aJ5l+wgeIGW332
/clOIfeKujiCTTSmmZgdaMzeU6xPVfR30LKjsVO0PTn4Z5bt7cofbnJ1N3Tr1qHS9S7NMsNYmQoJ
7hzvC3H8Wq9COoBGMM6kV05OCge9GjRKJ0/lrf0AwPcdQ2n/+XGHjSvg+DoZN4JrXnHUgzs5ww3/
VTwmeql1xArh3GPT8HNT0qZ9XpGPU163DbwFLfa4XGDUDuP0tZVIVVkBPTHQfQGeIUfALWAtZGwX
0cvR0JmkAyS2V0x4hESx0iYdi3c34+1l+eSoGSZGN4EW4FxPq/BLsB9LSPZ1F4H7/C6EMJOcG71G
rRk9nt0VfIXbQyzjyNS6FKvp/7HPJGZJDmdCzAl95rC5gvuJvtX3anbjbfymq4s2LrR9bJED49n4
YnAEd4ju5Nw9RDu2tuPwnwvxlV8icqkfip3wc/b3cAzeQ0FS18GM0mfzkE02pGKkl24l/9baDsZQ
BfGxtSRKkosWUhKl6ZpSrUUBez1WpquB2f07uFE5RjSC8+hgAniys+Lpv5Nc4hQ0SJSpmNYC9ML9
x9JhzLIHzQpKxQWcyURScEadnD50hZmLTuwJd88LOY7EaQSxrrhOl/8zzDChm7udRIdJ9C4PCZ1w
7fV/C61IPjvZH7kF4oR0dHRKyio33IxLkh4HLxXNDvuiBVfnAN7R5E12FMPAe7BNb4htkElenkO4
6QU1ShkpPN33bbBrui/M6xkIKjDdzX5XO47daS1v+pYzx0uLPY4yK5lLi6O0B3FJdWZqhhF+Du8r
oODNv5fWvBhqW6Bv//J9s8ukzR2HRJ76Nsu22FPQEsJfG7JjEAtbtPnanaSmlwob6dKwcWHnTUWM
aYw61xYxoCEZ+AYwrnK+fZLHiWWgIygO8UbeBjBCMlzS4XSvKPFlVNILHJ87kiYPE3STBfcrgQZL
r/jVOIODwVa15Jf3OysYSnqdrEEn+bHwFq0ePof9bb1F8CbJQj0TPlXfm/hnRJ0ucnTjjkRZyCU2
aN9BaWcrfk3s7YUFo3VUJzcxtlUZAFSK8dgQINqoaKljAOYnlt0cTlrzg1DUnyKVuvtyCanD5jr3
+Duy86T15he+2q09eJVYYOqxmn0kddwiUem+bNi1862IR21CPaxvvrPGxYYHyHaWkefiFIzoDn7I
DqD3l66IyXGt+lU0F0hyVpd/nEuAn2u646ZUXNUOFOY0ZLJKBaCSjK0M3+gbbrhqeCdJvjwXIQ0n
X+mbgkQQ7KMZ4oIN31cl9DhJe2xOPakkTAT1WvnMqX5PmB3e2TE3EXdnJb/Ye/YMQUaaMUUCrNY/
O16Hi2VUAh1Ozl83vwAJPa+V4PQCq7kdSFQAda6EnmVHSDsvlZsfLlnAhlty7udrWa6+jLF8rKPU
lJP1WJB+mHpduvT5sM4Bx/vO51V9OouaUlS5OKs0xCgwrtEuvm9VoJLn1i6yQnLO+wdbbtz7D1HT
p65uNaMwATv77rMpIhFQgKddhhqgyJ0xjQiMuOozquoFOi+DlGglwrsPPqW+F8qZIzW2umQ0jDZy
d/7rGdEttGJfPTy+AefHHupuWRe69xSBA65p/WVn+UDoPeXA0w7MIpIZ2KqCovZWYD5WLyrPd2eV
tPE8KJaDHcGfJq1P0Rin61mKlOg6tLdRyL7tRnqKAaAyNzHUJVDVQ1QhDZ4Gj8c3IZEvzQ5XF8k9
xGJPNOlLvfkKqI4eb1LqNpPgZY5rnfChc9i4RIhB0buHjEeCLKOhgNDC0k7kpBjG43zmLXeInRst
vwOrnKfPucaB6sigf2ANBgoZpCgGE24nEUOQdrCWNQzpfd+w74qbt3ZmkjTrKR+urvuHcthxM/hX
Tq3HR0FAT2EiYbdYZGgk4c+Mk7oUAzgW6ti6m/WLsAzD5Gryvhi+YpBJON8Lxl/tkMkzcTZQdN1f
o5ekPJ2yFhwiHaMidE17pH06PWsnhi6qk44tdWY+aljVMc4SCBoWAXmS4+ZTDQCBqGrvMY6dHtWa
e+/DDox6Km2MAIc1ogfvZtIdli3jIIlKAYMpmeTCInn5fCsQZy7nlquXOG6Rc7HKTuuzkZpxoHYK
mlsUktiZ9LtfhB8FKpWPVl4GFpeR+6T2PMqWorNpl7eH49Me5scY2X1XkVAK6kDcm1kc90IzhvBK
rNQ8tlQErbIuYA9ddyC4RvyFDMDklo2IBnX3wUUiKFWEPnPtlA2j026o8SDkRT/yzNoMClVQWE5F
PSIF6Pptd1//9rBveQ4hR0bJa4WPYtXqNBA+433Du0aZRDXxWorpIdMQwuMNGBp4eB1TFPppbhqG
2oGGPpS+IeE7utPUyZEL6gBP5//l0MmjD1rLl8DLgSS+xV5TCirsZKHLYKhSIIGEhTCL984/DruN
xb56NLXQabPTwpf6S4fgBhePD79jXJ6r+yiFRN7uzpS7KxgvundPBbFiSCztlLKmSPQypjTFf3mN
6+Q5THplgMLIKIEKmUO4Jg2x2nlDWe+YjBRAnCbYj1OZcD89lDjOSRBsuz1R5vbuz6Rlw5tBV/dh
cJA4QH8lKiXBYuFmcB7PwdZx4H6sKeRZfyu39do6MRemjlSR/jbRDFe1WIGRXQNK0NUNKuvqLsAX
p6TVd2fMlJ9Ckoqh02Su117Xj+haV3SSjZJgSVbg5VXB3+4JzeIOJaJ5B4w89CaXgvnpDYDamoCC
0q37WEuEvhlop/mUGBcfvpmbgu2QgbndbqyCo5UXtfKtbVHOfBO5tIA5b84BgDtgkUl5h8Dn1CW+
sKWj6sjQPwHfgzeQjYXQ5J6znzmW+BUJabvJdszYob5x0jRd/+UCElgEeJv6UiHZqRq8Gj35uVFU
PbBAfdGFZNDcfmfpLWGPEcbydHZfMQHIULcOe2R/cTUb5sQmI+fGAFXN6Za1aWQhJfTjvyrrrAsu
qzHGk10i6lZrq5F2sVUKZ1N7/DMyItnOlbcF9PFl+uDX1iy+PouZ4oPzSD/9b18c7JpcUvsx2xQV
9vR/Ia9fYG+YLHzHJ6lMofzzgQ1KDePUDgSBFtWMccR9+H28gx5P/xiY4Zh3YH0EVH5K+IImlwy4
wdgMQqM80TX/XgbJ0+3IlZvLK3TzrnR9WFv4jmIYAoKTUorZHg21Xg5A2iLwIAvL7qR0/cr6PwX8
bBM9ON6zFcTA18wFF6BTIIemUFcpaHuG2wzjRl/YhUNVWaE0mlX+fE5q4oP0BVJQyP/bNua90PlN
+YqvGCGMr9wcFkrlm0tKjBPzyQYIf6yxynVpy9poDNGmKSF9SqB6W5VvCTEvZk1sW+Bk73B3DfcZ
cFzNcXdqEqbO+cdOsBzuPjKzsYiPEDxr45eRYMJMrnzC6zXfbSJ0hgJgLxu1hanx55vJReCqio6K
68TIlBdPzzwWgi29VMv+RK954ryGItQjujrar1NKrj8KlyV5jcbieDujCxzqMKQasXvCAyI86sVM
BubklSrjmcaJUK5OtNnf9QIwm88j6wLFHWEB5dGp84GTrTlN+jQ0FHdqRTPPZt8JcU6GIEaZcS1B
b0ALNX+U7gbYCy1VBvtB1gvdSE3R/zh7NCu9HuIzh+9/E51J9gaBeMCx+SIhBJsPUmLIeEjjqvsg
bWhBqUNYPxXUJuRkriuv0dp/P2ikc+MyjbzzgzC8iPRBa0orJy06+5rZefqx1NF1EbQ3Kl3xd5aB
A7JiwuCDMgTsN0U5DflEMIMnV/97lzHbXaowHeH0gu3WbzImR2gL+hWGkwMSrYQUlyJgyM2PVLsm
HkiZvQ+dECvYO0def+cE6BsWm4yxSBEQiuzdcQoMUtf8dKoaeL+2ToKjWxmr4qG4jsTuGcJuRYeG
lB4ohiA3TMn61QsniupUe4wmYTAixFc+YL1tg5AbouEnmWc1etwl0SZGh9/Y3XQikY2HTp0c/YuE
Vcsq4tfyJfSpvXbR8Gxx5/Uq/OzzAaFtzVTxCCsLG6y6kjp6xHGiaIOghdtHDP6ui9odlB6AQCw2
95brZp/8nLvHrXO7BeHVVftNlbwOqQmGEcVK1xmSekKwUvQPbtHuJO2cJWxc+gA+LvD6cxy7YbK6
eUugZG16KMVdDF3SQ/u+G8pYTskR9nYfO6LUA/VZDxvQIx0e7Nd+Np0DfQdFeuoPBh1fWHYXsz+8
9hFGOygYxrHc5kDZodSRV716N1+oQROfiW8QkbqDjYZ2vWX8VXEc6dL+Wzcy43QmGyR00lr7XKM4
LmNZV5Z8hZTx8TYzPSHVEKUl0BBhPHbGjE//0vUjN/T8bEEVD/tKbVkPtau+JwADJjG5g+iBMiaU
Opt0MXVNcGEXO/gdEiBluycK2b87pLWJ8QIcKexTtuotR12EvabgSctwZ+Joy6qeAbk9jLEqKV6i
O2CvT64SerF5sZ8LCgtjOGDi/xg73dYCCEfhua1IfjUYW1ctPVoT1YNyXyvtqnHCuGxWz+Baoh9Z
KBda3W2/vJgK9MKOXmgCFutl++JhV95KtHKB+yj7fH3NUljtJkav93YaIUBrmdqDLZZ5X5ELdL1C
FxKX19RZMKVh62+yVZQRfqiKhrXfLfDgnaY+ZseddvOZO+iUczciA/n9p/0QoLQDqxiCmU5L63S6
qnmvaB+Zrx67+Ds5qYuj6S93yzZ2LngoIjvHH1SUApE8QWS8RpLkN8tY8wlZKwvK828BpOGlzf1O
5de5W5sUXMm0uaf5nUcZpY416w25rkdI3PvU/7GOYkDq7EQnlfsJ8G7NBphmVZtJjWsTsl0CVlzv
r03Egv3cPzvrfEHD8NXzzoyX3TG6Qkm737Du67wuekd+PncF/bycanTh4Q1Ht9N/jJe1ccR3OstI
D1hRDBV63BDGpmdIFOz/6cXrOpCwVSzImpTS6/gnqSXoax7QnGjRTqOHlUyT9C1wtDF1cdoAC6Su
29icnZRJMHyow5ag9DUBfEeFwneXhx7HN0bhVSRuXL87m6RAOcbAa4ZXJrr9o5PwLrR/UAobred4
tG3opTtEHAGv7ucJl7ObK9O+HAknosDqyQySSEkzhCLfEw+mebKzr2EPjKRMCYEYs/+iZ5mURkTq
K8FIfUZ6BAqyMC6Hz1XTPrFkWRYZn1MgjDkKIge+ShS6lIyM8R0uVFPYV0I0USTJtiO0L3WrPGk+
5IfUkoqdJeA/agoaiGE7rl7zm29TDzZw98HupWf+ywvnakOK25YlbI/AGj0pcY+Ux8HULTvcLJun
bwcOW/9kcjgN1Ph7nnswGcuUGJY84kssxeOqCEcNgIkSZbXk2dq+mHIh22tqomB4qRIg3vJdS/x1
INwmoxBis/6JxtYBjujNzoWuvy9lWf2cO6muuLz7mqnPNeppHur3NVqqTWQU8RhbKdQS4PPDOaET
tkY3MOdjXk6kZl1r1KQTKlynFYuAtDm7HZWjBNWjcKh8+ppuWHYcvVr7KFwGzweAoLfDN0x6vkVK
LNCDyAC1W777oFK0V/YcCdFItjUZlKp9/hxz9AmdW+8o+tHVVaPZzbq2+t7C7+S1ovcdG9KjxRl0
HdCPFPipuHrv2coYD97wCu2I7X3X7XQ9Bf4DBNFhcyExCrGVEwuUJfhqPrUZNjP7AC2pevZLIJct
XVOlnEq8pCLOGX9NMT9NKvonJZisDYe7o0YP+30gNUCauKaQIgM0BxvVmZeSNIXhhiZ31q8eYCqm
ijEI0EDhvnddPTNHCJXS7GfTHFgJeJn1zP5jD8p08EAlEnfV0RngAI/QP+6QtGJXHwpQzXNmMzff
hrZZpXPgLPOlJfPS47fF0ZPhmM+1DAmNTTyF7mbgcuMNWbjomOH8vfflzRvrHy+Z0F6i7a8l2Z9w
qFMDTPn5eQ8G/VGXqt9vZrjmLiYC3mZbZ7g5sirJqpYcheJZTKPPd4Wi1aDgJE+r6ojS+UwBqSIZ
mkzzlPAWDJ5IyWGws++utZSfLmeDkEbn4ek3zHsd/jHe76MZm8KndnpBGlyY3NJe4bzHmrVWzOlx
mHlZEnvjz0x+6nu6Gk6mdsjEmkmVD3iazTXonoox0LvIh5DEHZEaX1d2N+poDfLwC0BSjti4pKJM
VqxyRsPZ/yAgnlAqxgf65mFwF+LixsbSIRLEN0CEm8KjvWvUXANOMbZj0yHybKHYI8ZCs0o0BEHZ
OWdbcPq8DOT9wy3rhl2PcHdiH/q5FbaqmzktoL9yygOTTg+MagFYhNhuBqEwsAbPZZslRX3BDfyM
S6SF1qNJ6tczjeLxhP89Hz4LGtLm7Uo+ZN++uXPuiUWCTO1JhjwevhFZmODVs/V5N4xDjc02kywd
pH9mdLIY8m2DWHcWwJvOFOEaU+dKjzm67Bb7A+/2Gxa1ZZGC4uj/+bAMCgcAnAcq7P9AJR6DbSsO
SqZsyiBwHahmSHCdY2QduFA/z6TQqNlsGviTmWktVmMjXIjMLU4uBJNXyYCiy/FdEYxNgVqa+A28
dCqEuAS5dPdzVA2bjeO5pCYCX+JjwF1a0in3xWnlYHIfYNG7J03xny1BYEqVwNQaArimnxAYFt1H
ti65BXQTg5pJhphbrFP6lzYnbiTqXz46AwqLH/w8ynokRfIBNvDXmiBlST56laX9+L0vIVtCv804
SOCTGAT7NRkTZfoRDy+7JeAIzh54GrdTlcKzrTt3cL4tSaa+ngcQyLvQNd+sZO8UE0bK5AylTVjY
poWqJiLFOWJrruQImHu4MzjAdBxHjozMVVGlTha3MsknW4uFxOFWT/QftLn/aPmmsbfBGul+dCHH
xSQKoIej0fVXN+cRwbeAMlRWgaT057/r8Sm8BbSLOkqdTofOiaFlOiknKkvmc+JDYCGZJLTXbOQ4
q+sMUhagofLw9MBeyYMTTpAt9ah+MTJy3Z+Lg+r/vNYir/nvtjUKTFg6QrBjXxw6n0BttS9b57kJ
4LWaO6K6DYRTzDjDA70dM1pAqnfRKuplva1Ip2Ma7LOTjiKE28AH8PM6tvdLIDa7pE5chGXFeioz
9vSuNe4uRdeyoWFpHarEhfZIqxrNqysgWG2XZaUDY3zef0LOkukePHje3kE3t+NdhKUAA8f8VdbT
Xf7sGZEVrYBy/xDWVPj/v9FZng0XvB3xLIuNYAe6FTVcTPzxyttmLcQEmBWaeDLQfpV0RkMKO/1u
nKtuHIWP2564dQBx6kDDC1YwHoM0di++uXMqBV7FUMea13Pe9thja8PzAt9Le20aNZmykrUpvjG8
bsvJYWe0OF8cuW/mzk/a5UVcnM/6+yy7lHrUfQ6uvYC4XSkyoGp0Iw/RuKVO18GfZgIIYmK08tao
1NU3wcXXMBvHopaFDFUzvWr8MDPBYLk5iFJcYdu0/ao7lJSoncWYBupWiU0WZibzSbYMAwkPdDOc
dofG2D3kKUbB7aaNvzDo4Q6BAFOS9IJiEaKPlgmebqcVIdzXCGsnpycvM5mxEhJFx2bsMdSM8Sv8
d52MDgiG21PYzBDt6zMrMdtDXEF7q0fxFiqiAmByRDjX13sa6xg3ZWX+BKCHAOsRGFSZ94uPU0eD
Ao6wLWmk8OSqLtKWraJPgLWVUoFMmJoMDuKCmHDGpHvrvaeLmbrbYMBECll1lfSn/SGQTf9xQEg4
rFhWUym/bBbwTl9nynlclAUt8v+LGHtrQ4I1KBGzyb6Gc8Ft21DU0bOh5+4qA+A1vHv41ZSAnsyV
2GG3zecjaFTxcUg6UGHsVa9AYBa24Hw+Qk2WJTrxZ2kclPFm5/t6jHByPSyeB/GoY18YfX8NUFWO
E94hGd+eY+SB+1LtZ9Cg/ZLBjtYSOKrl7TBKjGyzyK8myjlCsgqeM3BnrIdw0g/x7ITbipJqy7/u
xure8ugzvUrIsuo5doT6zWpyJnn1mTj9Tw0ptXgKsBN+oDTCSL8FmdWlmm/Kb3JZAoEXAvF+KKZc
W859Vyd3Ao0YxO9f36+yJnsbwxzD/DFBW/K/Jk7Yg3MrMMvzavseWpsMCjDOlf5cg/jNkWUiK1Wd
mnbzAc0jNR+Z/u44ii6w2R6Lwl6BsXJQWCkXcspKVYhJfgic1Jm2C+pXGGsssfhBFGAOSKwx0t1F
idaQC4e9J0CqgHKLo5O8U07HosLy/lW1Mwn/j6vHgvSniCbjvYNgDm+4miOIG1hLIqkwrXnLsz3y
PDpp2FfpgB8wixj2alpZ8Xcz+dviT0eU3zzk3ehZ+CZ6QvI/PgLER4bgeXT+eFz+WK1pbCuk06NR
IPQo2RBG4WottsHV2PiXCQbUn0b3XdB4U1fNPuMEx/sVWqCCRnaexVY9Lcu1obIY2cJVpdUaoMSB
OZQc1WrS+33wv6mQMhMSxufe2uFEOSCbRdFEwq9XY9cLMQf23f75CZFvyDbFff8HyrK2c5uQAAFf
5z3JuOtY0w1z/X25SdZ9fRgK33mrBoLBYddQnDYhZTrDPHjqPmVJfHLE++y8cNbMUit1TSCUwrIb
EbnRRTTias8SKjnDdijUAXyMyx/2WFrelV5X8iWxhqlk03w7kDAvjW7T0DK90ciBbO455xXDtN3i
7zxwFahdE+G1Qog0iIYqiSzgghnk6SJp9oSctlWlUselzueZHBK+CPxFs1kK9yPQBZX6cm7xKbD2
mduijto5vVkanyOH2PS09acVRvNB3vdN2G3jJJYCCyoSNpAhoFzFqEaqIQaGmy+IuGZNZgEzpgM2
R3mw5QDZQ1FBfMoNrBm1+TPRJYm2dZMFx0Qc/5I274tbpBYwStN4O7IIoQjjCnrpKikxABc3gs7E
1R5EbVEoRPnKcO7Ly/aUXr/EVV3mpL6Tb2RSlpdCSPYvGl4dRDLuTf9Ch3L358G2LiDxQOqBMU63
nnpJP2dcanzaopDcQYT/g+ivcagU/S5l7kuixZxoVhCHa+dw47R/tmR90gcR72sP7HDNqLheFyp4
vLQax8/1fzMiXRXeeMzyQFZzCyyrdJTnHsq3yK3OYYFe/NDvgfS9k620n/Umbmd9aYRRdU4xKi4e
koTQsrxRANYLer9gGALj7kZkKUOkGt8yq7n0NqCnX4jWtpo73vbxZr8jtF1aG43u9UJ830KOGjHf
pGW/Kral0L8tovAmSaHcaQ82sQnNMSIdjV9nDR9gMwWGJD0A7V0Amzzc69UQGlFpSrZ8tfn6cExs
HtfqC81X1I5E7YelOrI1k82JaiM4uDJNZ/LarlZupkYWZTQjhLjIQw0d3aNO7mzDKF99ZK5tKSpr
9+5/RMoPbuX/gCdg8VfV70AElXn7mn7RvJk8z9vxyHDH0704UzXy0PjWO4jSU+us0rF7OepMe927
b/yg9uWB6d4C13tWLzG9zoBzBwvNXbuvbW14CswkJOM2LMIfPX6CSRnGExlnSslW+dguUUGjX9yA
hFG8v+T19s3mVoIMWaNwCsYKYB/FZeTo4ZX++gJYNsOo5sYVBY8i8/fEyYrxMzrnS+4JBZz3vD47
ulcAEVu5rCV4yozNW2ge2fhOYvMHthEIW4lpX9miX0Um1OGKkrm5QOkp5nC0kC5MvN64ceYOfUC+
GevZxw4A+JXd4nbOep9UijnU05tyULY/XErUzYIZfeY5Hot4S4RILQ3pDnsdr7K6H9pdODfzEOJE
JWWhfjLAx6GxnW5SjZ/FeOJQmvsr0+8kW0ZdQq0ZQxCIzvTz1lWF1+assD+b4DtgYh9NpOfyaCtq
vYO02coGsOOzWdM2r5nY0KbzfnXkqdSioq1CSABuN2kmQqhX8EmV0MA7APcnphfVRzPMx63lu1C2
Kh19Kp8IZxZa9y2dSgRxYxsoK550K/G/dAj5IwzGvequ1yLnjXHQ+N5kP5AoTr3GsVyE1zEO7irS
DZ4Va1qdpeUszEZlm/O++1wNlGMtPLIuhfD7GBIFTr3+jPPs5KPRCfQQZNpy+WrGU94+8LF86Zey
htmZkEnOfGt7sU/WiFoAOchfZevc1CjTcJReHDppO6w4hWSyHhmUrXNhLSiQMfPKIMUEMmmVEHfG
84EQC/asKRXtbrmYZCrHRLz/ZxcS/TBzicyE28+6fER8dKCaMSHiG40V/C/av+Cj3e98OBmp/eOT
uHWv7icLN3yca9q213XLZ35CyNMSBAQ2rvQVfzVf0olZcgEpMrppVVmHIex8CdRh59MdvaQTSU0p
+XV5Ntfg8DYlM2quoQB7KQih5ckGlsWHRCCdGNihqZU3pIaQ1F3LZ2HwEtsWG2IJPnDlRP/vtL5q
lqH0NSTmtpc22dKOPMpgJ6T8ObXcxYU7zeMitd1daFj9MM12mN+cZrxMJU9uxyDU+pUmXQ0igEd8
hREKWO/t1SYboZC0yHkrGNIuuhU6uIEcN+YFu42uMY3yE4U/j7YO3SmCL/7RelqXWp9fyFl440+l
RvdAWtrlIp22MezRYALbEB8/HigFYVpoIEcPxfALoVQzACyWSsyadiCa0FQVrXcZ/hRu3Wu0c2Zf
JRsX5ZvnGCg81B5y/x9y1BgGs8bAj1bH9XSPfRIOFXLv4BsgayrauTpuOu2HG0HFGnBDa9QWUeHa
lXszr785Oge7P0dFfZPZ8TgtOEholJ/y9OUQI3gaqNYj0ncdYJja6n0l8WVvTqMLQzlvqfXPMVpH
EcnMyRZ2i3VH/Zb7Hv3MM+/BJMcbB5x8W11AzlWm5ifTqYPhQEhr3JaSag0Zzzd4UM0/FpznuBAy
4FGYsYW3SbU2j5pf0O8vZAHuR71TvOF27nYZK0vGE2PakK/sW7j7bVuSE7HAfUBLyAkpneTCA41w
+iUR146q7r0mt+wDaSnX8+BK7Jc6SMJd7rWmd9UZ+OXq0inEuKwbs1dPquGiQymRKNb8f0yZugiG
WFy2kQk91ABC0GRoeL6RfA9Xg/aV/8i9JXsZKpB2TK4hOqh95O5imbOPxAISxMDjMphN+w10CRWN
mfAu66ZIU7U9nagS6YGJrFKm7UFMjr9vKGXLvL5O1wfzYVmEkv6j67V7jhPlHca/KV9K/aC/rJSS
8eFwgjKCaLmyJzv7FC6hZvzFVeDRQ0uQFa1p+9fbUG6o52wO0YbH6JMhgcQGuc91fiDd9ad2KdxS
dpkern/vv6L2AguB7odMhppUw1Hn/Hv1ScjexMMLm8Px3J4NW68lfL4F6kFoVe6cYxkimJ7e9N8p
KKDx2AD0sLZiKi71XQhysy5XlytJOhSNh4mvu5WaXcJ1PTOsqLhtlHPKbE/sY+w/Xr7QNX/fewX4
+76MwfPnmmpIKCKbVhwasoIDqYiXXHOUoXpH4T9XCh/PaAmPFiIa6JfI0BE7R02QvE5Olm+cHux+
lmK/RMYMjlZP0B6zO6vvZQTBi2lyHw8VPw+jIh1n3TlHm0/3yFONLSVJG1qluyVh6U+9Q3zge30y
+HjUTfps8t6mO2dfoK+tFYLscSYTe9A7mBF0/D8Qh+AmMPCaJSs28+DKubi0lReTb5zGT9RHXI77
oyQvvLVxkKlnCQn7wm5v6YszWW029q8c4PDeOVS6B757VeSiTjxHqhrw3OTIS0xKBgp7WGkZ/Egn
CyMysAqrOchdygG6LaC+nlOPm/1guTHyNRUjgZfeyBeUA33U4GQmDb1KRkqj5G77Nganogd/g0MR
VImTnOV3Be8yAPLPZ2FKq/t75CmeTEPO3MySr19lYlTN146HIxPF3lITAS3qDU3g1+QGPmcZPc31
7mbrIH3gzT4+h+p/3e8+Bmf7lSL2bI8A1jA0oUf7tU7/VOxh7XjPM0WU/BbcA3+fSV33UyLheoow
OYsR5vZXO3mRaBjYw5MhLnd1+AvCJKfPnXopk04hcwNiSdNjsfgrPpPs9QPsm/u3xvPIYIoD2gYl
6HZX7qAN37mZtJyWEz0PE8ZA+XXIqJFeKNuA6pzoiqwYNxCPYXiT26I/7bfhevP1kqjZUFzdE5lE
3xLiJX8qUtbLG+cmQ0VVzndsfJHjMIsXQyxgp+PI2dM4UY7yAFJH9KYtio32WX6dN892tGpZ5JBj
bsVYpvdN4Uw/JWfm1GTecGDFDBVKmos94TC66xSYqfS9QT/vk08FOuq+YEl4jkeh6VMl2tzhOKWp
C5zD6PkZX6Y+GVn/AWUGY11gTggnt61TWXtTR9k9nkuWOTKc8REjffPmYlPmjgyiL3c1xay47sac
/eF+/gdJn32BtpTYzvjgXBxNsWgZ1j8l+8Pm0li9AT+ov11b8tUULuEo5G18mF+9Mun6WqCrMevg
oL6JdvKGdpf1G5XSh1TaeJpicVVGTzXg1pPDGzbZoLYPJY1jWi3TtHtL7Orkv6Yj/EoJOq5u1qrM
ttNnnZyQYk1mnfL/MVOy82EFlmjyhdr4ziN2EF+x7tqlKlIQwk17T4BlBcoT7USXrtjp2iooFWnA
gFAiG5C6qZdXH42NQhEIYZLfl0iI5cLPjvRoU9MQ7f6Z4gSI6qy7JEJ6VRUcmrS5p6UxQlm2pzor
Dx1p4x0UqMSRHYv2kufUCYjnnmUTv8ffCcthlsZ5MnFuTlDQveJJWGFWJRhEUZWaePPehSuGryRE
wFu1MUlxpnovXtGHrtanPc2ct3Nq0uhWAqvYzZAp1RDm8FkQOtkhzuYjcwgiWKVPiNPnwRxo2CJK
aM4kGd2x/hN01HiTN9Iv9pumV/ntgrruCBGaUrRHTHJdRuwMtGcnWmRBBuoR3TNtv6ewc/xoFbmJ
Td13qzC8EKblpbYbKiPi8zfqJLuHNSqxkBagqu/9i90UnxtsZlg8BQqherAX2I1k/rMUIeb0JuBa
hxp8Rkbjw4SLcwoMcurqknTXzoSxFn5WuhMzGa8akK4UEJL7WOBNoYGJgCBXhvDpgCgoqYeCtpIC
TFURZzob2qLUr8URDLhT7ZPmWi4TUkdNKNFCNIrREEwP0n7BX+vOnAVYiOf1cFOHNzB+9STXXfYD
U7n3xj8ZETwZELipjhVs/cXQysOJW91hGd3P95w1XAl5jNzg7ybWurnCiz8zP2JAOutJHz2qCWHx
hZRmdb83l0RPrKXncMJUk2C5TLfGqmakNzRXSuRne9ZnAo3WiERocdM3gblg5Tf/rW8u6pG9OMQ7
R5iUuJL8ea/HXoNozSttnC8CG7bb53TTiqTjAPhCeoIj5DFby3YmNCgltttzeAiO38ffHIUXdYuH
8njQRBNYjopQwJmxK1W/ifu+4vgO1b0ntu+/RJyMfsJIp7dQqtqJczRSN//CX9yNuJKwc1hKPHZZ
wsHuKi6BYX/oFBrxFVIF60ayalfe/Uk2wfUJP0V5S3hL/Favwbh4Uzpec6P/1UCJh3c2hz8EPk1G
7Ts2P1DTLWNoTG2FqXE/Mcy8UVnwIir1nvMj9IVqeMd5hrKRqSDIRLVEKHbsa1qQYJbgmCLWcf4e
3ctrX/gqc2bB4+88CjJBTRWnBXX5NbOfBpwmTCsSQVWpRYufsM8x5g7phPl8mt2PVk62od+QiZ2n
c9ErwedZ+OG31hvz2FHQ44OjQThJIyP3fr/nW9OyddXDN0VWGNYNsR4yO7GRkydxtEKQhWcT4xjy
i/MSW6Tl/16SjFBYfiAVUIiGcdmBNCTk6/o9m5hsZIEyMrHWL0lo3bX45d4xjkWhK3viqwJdC3bO
TZ6gy37ff2AR1Aoqbdb9XSUxbePYegFGrtINORHEw1EsK5j9T07RDHYsttm7qPGctxLbMDVWm4bZ
0L850NIFZvRFE9KOH5fosjaFWAStzVSg9IQ9cFaXy8gcKMx1vI+gyQGLy+izqxfWSEe0KbpLEf3R
QoGgf1MLcgvaCcUjH7ftMv3PeHcFHF2nPE1WiGhkMgtqLMeGEcGTHSEoD1ZRxtsom2eJahfLYmAb
gjjpMHz1R7zLBFPRwWdOQeLIF0WA5kp1N5YoKmXJZFynrLsx/o4bY6OAnCFKGParqcrxJY781HfV
XVE70xM4NMDdJd+j1Ab/hiVqE7Vkhor7vEpHPk2w1yItjzv5wQ5p2swWPKiAqyW7mhiuYYct+L8G
RKuDyDzwO/xj4GIpBFXU7Vk3rgIqKTqqezGG1fnAR9mMDwnQHDbCop4frryhCRE5upcp+Y8YtazH
1fUwvyN3PNZRnpwmvw1td034fklEjgnSD8ZSzGd70efF5i6Os+AdEFh7BxXAFUH98LuSyd5nA+zt
PYAM8slK8r100+BAwEDTlss1fJ2PCma+i/EDZ5rE6WTrsmlL4Ty6Qf2QIsM5GBI/sKTZ/WnL/vWV
xF4AG8N5noJM0baNGMo6ADYN7Kba+W6IC9GhaitL4wzsQmUUSaLBw+qrRcXxbXORnNssQUDNAduG
NrMfHVIOCj0arhlm0LzqRY1Ov+eLjMD0xlut+WOYAlvKfn2k2yonLLZtaNZRKBIwcdWL149lRQuX
IZl26Z0e5uMx5cx+UTOykflch5y4rFftspPaCnMk/cAJ05Erw8WSoKrqpQXwHA5I3d9CbBDHN997
XyyV1DpKsPytajatiprThw0KLkXaPMhJ1UrnIEugI7S4tePJbySaHhpB0EA4veuP7v3CNVLCeB2J
qayXFDT+5ldqJK0fNsgAhr7JaWtUFzM6Rb/nPgCNgeJrzI43G2Ifzjtvf2PND71MLV0sU9WO0gew
pOGbkKt23fL6OnziyXieRhCgFi87WUceRuNCbHkiy0xFJxRH5b+xZQYdnigs0kSUacxHNj01BoOV
CPT/8uoTig+S+F+/S8ozFEMpdVgpSrcro0hGw5OPRT57XkzQbQf4w7OFefiPxKzV7xNTGXIdt5Ld
7u5+vXuAJNl5bixoSBWTvwmmp12UG2XHvLBtCqee3meLKPc8dzRcQKvxs4DgZRASDjbRXk0+55tB
AUb71YDG49FveP4Fr5G8hwDQiecG1+dBvoscQgPXVTwwuR3nbFBckC1LqujH5hNay1SIs0vDW5h0
6If+eGbThAA2vdeRMEKAB2crR8z/T5K0aS9d2+AZ6jyqbyBBb7VRewEeUEb12TF5+xcbqEY7qJ0d
g+nNflbtd6rtC2JaN9wnmHU6tRymA6KTkjw72eZBP1lEYGoKT08CgFXLcsqTIkTXDZG/3IkvMfyW
sog1lf3lieVnch3CiutzFk4BkRwxzpvGlqwMXMNBrTuyxycdciHC1qW6e5YGP3t10skdHCu2DWNl
ZDFdWhl+d3Rsjl2ArtRhoU46l2BLbbppiASr2mkvM0MlIXRX1ERYEezMr38a7roNpab4K3jiAcWb
bnQVQ5M7G8y5jCx9CpeRNt3z8oM05ogAmxLLIEnNiNujI3JKVNDurGtHcEXMyL2oOSYqQSqy11mq
7kCkUHo4bD4hGVjOLWYYg3dFFEzIWBID7EkqooS4Yirv96xLSUltJGoS2wd0rs9iqvXSw0Msuyjc
YMWUG7aiaH2hSFQOlFFDB+Trwh1PL54zHwDDUrs1AGsqtDVECK9imeM3iR+E9JLGeQ5y8qyyfFgT
yC8HRdmCIENB649IFFWmFUkdA4EGmQwjW/WOolHaegNZqIX5P7TrEc49IizJPjw8KZGlXm6MtVuM
+pO+HW53nFTiiMXt4dml13Ucn7EqW+AidzhvLeiD/ddCXBG+0rlGrHbjTFwcC2j/wx/2Ix2nHLiB
qlj1CTE2mxHqB+G2gX3Jnx8GgsdvjYP9+gxglu/Jdq7ZXi1aIAapE025Bu2JkAp37IjsEnRgyWkD
0NHXBVtpXQcS7wcJ2dgOuQIFaeH4eOwYKDyhFgPms+6TcuB+sqLbBmnbmuIldv9mQd5s7WsI7oBe
TB6qmedlMWYG67owRBACYraZ9msW/atbmagm6L9TeHwUZAwTt2PneYoSkAUFeSNGAPAuo4PHp874
cwmmG4ZPudWHixjDbQU6mkbPvqSQXRdDdivWsABbbAlPhGUfjfDshwqnYSZf6wph3DVrQ508vbNZ
DpcX7+ixHUEevxrfBMtxWY8j8nM/++5E5XPg4zT/et4bUuMFZbsAOMqN/3hUWt3DjvJGCphqYMtm
OoEss6yBzUokVK9IdsbN53ju+VL8wErYKN2ANDwyhHU1pPji0zdCSCq/k3GXlE26JfTCvC2Old6f
iGkGetrsjbm40rGw2bjvR1dFvRC5144rgX1NYA5QQ2L9cuJc0jPj1w2c0w18rYdbpbBSKCdqf6Kh
unfmt6pC1imFRj5y5Hl98AH4hUhFq4INUfAC8Nis3Mj7/Rh5ZtORERD1mh139vXv1yvEZeH0Bxhx
WSwJg0FQoWxpkLPq/SvXtnlNliF3gEe1jeW2jbbPl9GEm2JSadGmv6kBFSHYmh939WG0TWOulLCF
GCWSYmsOzBSdZ8NBMQkc1Swp+s3ylG+egEvEdUuxHSHEU+0ERpddwM7eE7Eefyuf57i+jlw0Buol
kg3XsRu1OfQTSc5A92Fu4bEAi/cGXuBKjVjrmLnhwTS9l7ry9UKg77q1V4UL7OS5VpWNG7ywBbEh
5nFV+r5/24//a8HzCFPVoQ8I1CnvPpVU352VF+ZPnfyQAm5DmMAhqR1fq3oTwImOStJudpCMmrAD
zP6D+ttwnRrffSeOV4ii1QvOVtueAkG9PflWBv9x+9UsYYmsdjxv1loEdWrNrn5RBhWsCdEeeMex
40D15AexGez2BI90BkI2AvXBW7EI4ViAvamflAH2JZftPXRRMk7JAkb30AGC2A7K4qZCb9Q73esK
8kvZyTE3ovBh0QsrZTdAZt6MLA9oqwas8jd9lvAU/dp0lfnmGI/41dnF0NbVcSXzQ8OHzimjjxTU
ZzZePh2PVNFM1XmBeSQ2Jt8f7M25rVq6vafVooXDyTKVUm9dbL/58xO6HtDahNKpR3aQE8EkOjDC
Ak1g/dxVL4XcyzcAw/miN+1jSlDLae/lZRUQLsavnhJ9/MbQxoTA4D4JoFhIp0V0Ifj0h7wATN3u
D0T9ipVqiB7oTJB4nwalj9YfYqocGyrgfZPe/TAeOUkavXt/swk50DZz3qkQb0x7StHNDN8FQDHi
Ybas22yh/zFGJfc3ggcAoRdTrrosHJmPxGokSIHjlJ4EOrWyqXec7mzTNwra42MNg0cAf2Gm6Fjv
2Rt3IlE2sSwZ8nYzA/EDOVeQca6sly+Oaobz4SIPBizprIDYEfS/7q/yFgFTAMO0dQ5rH/6ux5Uz
3WyAED69hWiY0zQlMs7mOhdpVNC1X1XgeSgG/CxIhB3NyvBIhlpIDSHc0GjfTJxWR3nGB8B+5BP6
O9DPZ4ofBU2gAAymdqG9N4Hbxl6RuezrYbDCxTe/8MEz0e9IbEVDJOsla+eSumuVkneqAQJ0MnO/
Y73A13G7geW65F4a+oPetkmnXS2WPjSkJsfJ65bBB5F7MTkmSXeGMQQwix6D2W9BBA126rjksx1M
2aIy7wgAtPY9lXJ30h+zk98iYzmKNVdmcJ25i+8KoF3NmrpPH0Wa8g9yepaVVUZwE5r8sNGSrfDy
HTrltZyX/RhcSWwAIeXbwnaPCFBAsvOzVcZ169zAEv1AzKeV3frxMmbhiEa2Ik6UY5sfsNFAYdMI
zPT+hlcIgYAPB2EbC5K4kQQojNMVAPXyoqNu73Cfc4INFnL3Z/86wplInE21olz21KGnydiAaqVf
RnHPLSLnUhmqfaeC89yZWWO0JzyHVBPRfRA/Et9g24J/xwsT0qROr9/oFeV0Olq+bINsjybCRffW
ImV1bLZZpyvOLAvjzT7VxW+RvXrUREMa7aeL7XgPiHzOAX2L5hTW7+OrQ5vbzN4/2vq0GkAJ70zJ
+8G4OVwkwuKtkUGxeOogbT8FjZvv8gT9SPHC4AYg2E2EDaVE598VJNdE9mAD8ITPudoHlmneoVPL
ALUDx8my9p3WxmW6UKmwjMxgPX4AMK4s7qgxO2IxioceHhccNfASciGj03yQZZFS77k9enlv0gvO
8zHv7YwM2UrjirgPqYbwcjm4FUDCTE1qR9ZYrobITkfFBOyAPplcBGca7P1kUxVv+yX4gA2pmF96
5VwhmWIo7LNzziloMz8BiAXPrp80cx/BwHm63egIdzOHHwgkiS++QKxIfEO0lufw83bkmeuZYsVy
KENk1IvbpDp9hdN2qbCBCAkPkh15vUZeVCfJ1lbroLxiQTTFHxMV3AwFMKTsFTEHpEFDV3IzvDNL
JWNiS246jkYhIqasoMB8f3+JvtEVCTgGfMcpae8hWDWq0FcPYL71hZe3mQn6DXKYxmuVsMGMa1EQ
2+KlziBTSDhMA1efy/KgOtk/dEzr8ksmZaxSHWq0OGYdniV0W4b/Lr08kq4RItOzbEIBKbCW6ITh
R1LmQfBbl6rTsj9Rzeomh1F79574gR8rhuuz2Fy9GAoH3lYTJjT1j7GTt/Vy3dK+bZw40EX/RaXm
vaSbf57uEz4Jn8mwLDUBVkp1lrz91JaASpHMDPSMpu2/vU5Ek+jQK+bkwZVPnRkU1UKCLqDlx67a
qv0uAxSJW+ZRIuVbZcb4OT3w3QD302+fnFUqm/7s50oteIbZLnDAoYyJ/JU7yQ5yJziC5tmWqVRk
7sfAYz7s5Q83tl6ZJygngk7TXcqZFvqw+6ZYqQ/SkfnDidp28vdRe2yJruJX0QVwpxX21WPmR5mR
taqF6YQOdgY1gNUty3PqZaScwlS2cLrVl66CA41f5YtjVCKWRFEP65P+91BZd2Uubu7X+pVkIL1I
CENe7veWLMyjdpDWEpRyN4HQkNkfXyjY7P0BEk9J7Vswu84grckuf+KrVUuS1cHx2cyqyKOkQjiH
VjZGwUw5jYh77cvzG3x37k3crtW9AN3OKa9xYmqSMhGVKaftqH4fBu9XL5z7R/PzI8uhkrcrUK69
WEu81rzTH3fkrP5P3TfQtnZCTGg2pImJIFcdOeC8GTHJDi+nT/Wn/D3pKBPEQ3c90LrcraLZAnCZ
VWJQCcU7r106Xc6hkRhDvT8ZjGpkbbGSbd9yosfzExdU3zz415YntXv/6H0xOgL5IXNU32kYO4vm
/BCkgbq4opQjht5Z71k/hycvpGx6GXGpiTKBqoDEM6UqxkC4mw+tB9c47gjehgwe5DdH1MwIx3sG
MlBmlhXUFU2MWdxhKHWYF0sieUcTajMrSMTsLbNKJSJejOdgof5XKYUETOH81NjX3a7W2iH1wjfm
GNXMtqafTOfve+Jse/xxDyVEsdFBon7ZILneOTM6izp7QF9a9tu+jbb/Vw5oAvSCd91cKa65sHcI
WiJK48o3M4WlQsMsE6+IVH9i1NznqIylzkbnf/C9/4D+divTUvnemts8Jin1Vxc+tdYFZ4MR1UlD
0lfzR/0WW52BQTqFz6kgxHGO3hv2rSfxR8JTVmxjNFwVU9AaIChv6q5HB7mfY7N89BGdDp5znwf7
rcdZlNLpkPU6WmawDqc2b94qntvr8bXtUoHMPfDz7hh+L5/X6wn6t0Cv3ZX/0zb+XjEJUQJwR4iD
CewexIZ8XXMsFNhXPzJJ4Mn8xxxEeJInWkVv20q3W/eimJkyypny/4x9U3ITV959pkQID+uOuU4l
83MGCOwaLl+Jq12zbAfCIuQYAGW1S0CDPe4mLCi00gXFNo0MgtadJEhENJffgzcYDgVJksSR2/Ty
0eehuadq31/P8P5Csh3yJcg2HzSgknFLqrtjnhd+qd03MFHRZDhBTKpN9aeTZ2oex0Y4l5zITGPC
AxmwrvCBmb3W22YpRuBwFWlW5MkOuVDryvWXeJg8sz/uFzwdcbF9Fn0rvjUH89pCw5j8LGGRaXzT
aTmZRUirDHEdtE/oLX1Dv2vskcikS11rg7sLMlticU3b5Xx4+TMkozsLwdgElyUU1ti1VqUu1l4M
yESr0BBZQnw1W2bWQ1HeA3xXe8vjJ854JdqPXFMZlws5rbMVBiKTtge/aupLaKLyPbDHQnpxxl1a
8E+eGFD1iLrXllW1AdpTZvylhIsSM0W9uopPMd1szNRgTsirIXMyWzFPV4pjuOQrQmkhqVpWJmJl
YCZ338PKums7xxbmi1SJpi3H/HuRQBW50vAyYkYEAB5FCty/T61x49HQovloXMcbdWbuya6L9Ecd
zlvDaRN/f4irUu4eP2ONe6z/uBFn0W9TGVNfZFSMgz+sCk88xVXO9C4zT+8Ehp8RqRP9zq3Gf1Wh
F4dqgIt2XBKpryBruOYYn6qCkUOGR9k6VJjwqx+R0uRNjOJTCWPBIouBseBrnL56fShSGNT5LaFo
37UR6YzZlAatuOpBZiQ8VPYGLiXS3zVQiQTuROMXTBTkD3Q/w83l/z979y7H0nH22oRtFyCawfQV
LeKqq/oZdEHZ51KWgi6WWptPrnl1RjRyQAW4mo9BWgm/2yESuy6KRrb0zJ9LN+ZXnnYAE4xwAy8x
U5tI66mV4pkYDje6h5qqZXLa5XIXyGM0esB0YgrCpzhsWwk3f8QVYXYmuSd0z9hBrM1V0nn15d4o
7QOsb1OoCCDwcXkyD7Z4rDx21xtaWGDEE4egP2nw6W8kw5FhCgMHGpSQ9VVIoErGAmGfLsfO551z
FjWl85yNLGcJL1WuKpG2Dh6UZIPyDuJhqd2Xd13Cagfbtb6Oo69Csi0cvP6H/7UZlc5Dzt1z8Voi
IdTo288ZU95YGv8S4wcV/rtTkDP12Ign2pJkblea0UY0IVY07ytjEDNXrx9tEcypGqMS3NdznhzQ
SoV73c335/9PWJymJk8FLLqplGhw8DAKbIP0/mNHbHNePzv4kVi7UH3wgZ4Kh6iJx3wwDEIKUuX9
99quL6YhtRLCZ/JGWKEfLFFEpd0CiC7nJZ+B7awMmXsnRtbs+7S4DmE8bWsTJy48KqB8rpUbhLhl
Zl4PHkM8CMgpD1FpxSlAxdaCqegKf6lmyJEL5NlkAO9PBCbU234VNIu1rzFHllzn2YsrxwoPCW79
/gPm9RXqp5kBmLaGGpndzB3D3KRY39g0OZG6VZZ7rtMmO7HgLXOjGR1bPuI/AIpR/hAHkRuU/9TN
IiBRPRyIdpoNDzwOXbjliPUBoBqXZAzJl3TNIEZytY45kntWUST5FxDRPeXbbXSOiyj1/NI6S1aF
39Si9oL1Gv9IePgmCZwRLar3hcTi7z5UIa0GFydinNO9dWLDt2SyPKs7xKMQ6nbGShbGjtEfxqVp
JtAc2am/cVR7BYmNlH9LAoyJhkLIsogYXxvBhiPNcCgxE0rdiYmznUj+Zxz+8D1SbmkSgWkWaImn
v53pqSjDaJYH9hadAZ6uJoc4IfJzQ1lVQxKkrlbey9pFt+D7cwbdD1hBgcVtPQa4sU1YlNIiM1H2
bbhnBlyYFFsTc+H+dETDMnHwJIrXvpbabs8NMTp4yjh5Fg6QOzmMfi9JYdoZ04pomjFjM1A4DpvZ
7YfKPUQpK9eiJGfO8aoBTDn/R21UDkESipQkCCW2mhn8E1crptFRbY8H6yfwTTBGU1ZU3oCecsRt
K/fsUbaUh4kaXjUgngOsY3dWR2pWwqvNTw0PqXqCfJpj90d+If1OZeVDJLRaeHa3UjDxO+geLILN
8L0ZzWo8GEUx/srxIguVU+cHYbg4iDp0T7hzbDXTMX7NK04IkPkveKDILfK+1INAShjdHvBFQEqn
AahqW0nYTNLtXNJYmlHxdAYZViEf/PJC1WNMSAgifPFautlcdMTryl58Vc5VNynHGgpgDFugbIFC
RLh3Ked4X5PsLzbmYC0zV2U00/Lpzyn353tl0PpAIv0TwuGjfljs7FHDkUO/J0PZBSHvcaaHMs1y
oS7zb1o38VKOkzgeROoCaTDMab660vhAP0rj0bF4AKX71BJYrcVa+sKt+BhbK+e+0aurTgDk5z2C
RZ7KlPBiX9RaDk/9woVjFZ0mu9NidQEaqIp+Dj9yOfhPvKJgf2IU4gtG4L9DKuyKwDmNvrNdOzQn
ZvddQaPZHgWywWtzVzN8zJ0V29VgralH73g2rJg7u3snLepwkyyJzQL+0FwsqONfr+KoV6atyZH0
jsDfonuISEqbRGgeX2cmOSLNqjmdqK/Do6MsTHdXNMxLrfqfS9h96yp3eiFURKwChfxsITMp6QCH
Yh7MGzIQ7uSPMzL4/PYF2kEmNZePmogGVfJm2rys0u4c0hgO89ROzjx1fsG2zaApgxtFgBxjngSn
XRH27OxBDgOfMeoJrJ9KmD6DsdNSljC/5LOkWHwP1meFS6qIRtCmyt0jSmcPiXGt6ZZxbMC7+acN
uHxyQjnnaPe75qAm4B0J7RMpY1ozcTky3PKkemyy2ht9B3gnWnmytK/8Qnvif4rkzZV4C90icZwH
AlxgMj++pQ3E1+CaG/ZWSvKJTBDG66GUTwyX+5K6cR8JXqFwgvI6jqdMPnAuDifFeCj4+MsRW7Gd
e2Hhrumatup+kXB6VkTm/ccKwyyUIyavg72oI3wgtzVyh4SJn3oU/02+AWk7miHcnOOI6Y/kLHal
yTyvJRtE08VD9IsUHYlOoFjXmocF85lAjarL6oe7xhGF5CnipedA/KXiPegdu5n48HptgCz7LJlF
0wTKmYN4yqjdiRxRaCZEQBKiE5vAe2caVLUHH9wX0RQTpbWFx8b9ReBhkWfvChTmBs3AbOT7MWnM
siJw1VjwXLKRuCT6guK5ZP3qzmF0BaQJsNWZk+iJ0LGVF2wp+DT/2VNsg0A473pkiYaTo/dv3IDk
8dvJLrqrcnbA3Np7cdGwpr41ZvxDBk7gm1yg1VIWC+7AHuURN6a8/fNHcnYc4rRaMC5EqLvKX4PX
SnSocaJSuPKXFGCkoPSUwl6IjYmok9absUCIFyujiwzctUyByhcM7fXJhXu9ttOhYlo0rEkZFQwx
Z3Wo7grviSEp5r+i0SvNLrn0jyepcQhjMYa1tMSCmureKO59e466nmn4Wo1YDqdI6Ns4D9tX9HZ6
w0+q93ycWZYMU/vpz4zWwVVn6FTyaVlH2aDbyaoZsoAQtv+SWXuhCFzUakmOTY3fAHr9him/4Iak
exaOCaeLAwUCTfKzeIR87nnvx3FBaRctUqrjYe5pCe6Bl5yufrT/HtdyQM09lfgFmZrMmRqcbus1
xYpVFvqmkea1GXPWfGbGxub8V4793RYiRWs4akQA2vY1ay6mhDTbNKHGqqRc4/teqhSa8qVF8D/J
X6+oB9KDf4TnRsdmqnXP6jJ97SeOi8FbzHbOWhh+kNCOh54WDebkaTpJGekAkutTIjQ2/o8wbJtq
Y4TdelE+as6r5g5uQFxpmUwsQ/WhxceVS31hZFNHIzY+cP5k9LAhWES4aHXIv5glS4UqThLmNkdY
UwACwVFnBuyTAS0E4BAE4V8Xptmdw46XmmcZ+oOLdIoiMLAXNHzZTJoXoe7T/bm3VnX8VGdqBvSk
pCUCNrzbyCQz1HMQb7yScDdP6/WLRqVmWlkLZdJHG+3piE63p1AP2wV8EQ0rjdepkdvhlGOUM6Ik
+YZPhT5a/+NMRh54EfCbver+MhFSPdzouyWOU3NtVG8af+FVVFrclGDrBIt14FhX2Qunulkit8ZG
aTqEoRX8tDo7AuUNQIm3Itbko/ctaqWK8mApVphkkWqTe6fv2CxmVXmOr1Sq26Guq+ngphhzvP2l
oG1Otl/5RUQ/FNVzGhyw0hqnU5bduQ6Ix8gDIifUswbTMq+ogyNH5OhPhLm08Z71TnYGjYGrBLrU
mpfen8emC8VnWdP03rapoysNOQhDd/T90Mh41wwN3BQzlGq4XpHB1xf6PRR4ZonpXNIzPg9gZsIg
yVMMWaopWzmT+2uajH8j/kAkgGF6EEHcSh+AYI5ah9Lp5WJ5Y6I5+ip1UAxl2Zjz5OPgp0aZVGF7
U/+g8fVeQcL68txTsRnjvnNUf/Yz8KFqCRzkZeFXQrN+puWFE7iL4Ck7V5fAu7sZqwliwW+sBlc1
u+uczNxDRM4+ejQg6nw38wF0WGGm8rVKlt8P0pbKgdOokuOv/ft9sX4ndYVXrhQWczQbZ3S0tnLf
oF2nNVQoOCD8r1V0MYWfcBQkw5GlZiSTIqaFuG67VMKwq+012C1KWgX2BhuKycN25yimZ47cQuDs
wwWBT5eQksQcSg+Ns9KJ3RdvG2R50UBPTubd9Jhz3ZNLEL52TFnfgrk0ruZWZ3iggRXA2IwkYlAe
Qwm2uGUSXRXNvxYTA4Pz3b9GDQX8Zf9TWYhOHtkT+k6GKxl/jLT0wza/9ca4PBkBV1gqnIKUtJtF
3plehsq6s0hS3jx6rv3Ha68wlcbapYAc5OwMl/tdef8y7BmOYBX/PLKPzSOo0WSwfAASqplivcgd
bLscPbzbNy9bGtEnUMOXFLv0Spswz7r9sXOhIQo+Sts826ykKjfQ0glwm4kyDt0nuiO1af0GRtc0
FYV9xDqnsyXWYYUQw0A9DXgTpkE5+xC6nCM4hL+GUyIcXq7IFk/KLoeIsy2AFnfhGSN6KDyy9FWb
Q/zdE6H+RvMExC1+sw9IqKLtqTB9IlTYHzDtwr1fWea/4ugCCY+eNEIoKiTmWLtAzz/8WWWWcWZ8
3WLibG6qeraaS6IAVuSOzuFuXmO8BP4Vc6sc2zeppVI1sIfO/cOwFBKG8bgKk/nnp6vlE1LXR0Gl
df1FavTMe3LHIKd6xdv//t8gu7KyU97nYSzOZQ/lFqIm+NyGLm7LRc15BiLDrdWYx+GaBnbPmRV/
Tt2JF0SGZBa4m9CHNyTNRCEulH6XxYmbsRHYiaFXZMJerArmInpWh0dxV9qomI8bINn4DmITYx/6
35hC5LU9GjPKpyAsURv4VWGFQZCq+J0j8W3uAktOMeuxXJmPxSO7LbcRclnzXRueCZ+tRt3Weyvj
XGOxcX9xySJX6UA4yBwdpV2IV1J1vwrX5yiOETmb00j9YKCUyDfrnKMutzrSSTlGB00HeiLdl9s1
OfFqdlJoK28qwNSXOQmtaWZ7JUIGFy4a0TOuE2c+Jmf/dxgMcWLv4Wjgz9L9dXP+102hBIKHqKWY
qUVPqO6DyuDtNku9EOI4Mx2S9LVCWhY40xj421N3lGdNWT8TB33wUbe5dh80EwKeykeni8q1000i
/t2TJwLLJ5mrT8pWaoKPF+tDUi8tJJufjvQmuy4tovW2slwrLZhiO3ux4LmLBYJmlqEyjiLXiH7V
GHK9Ec3CIu9pOXyPEGcOwGeFRz3DUR6q4REjWKjfTjMLnimoyJY7NZl20D17h7Eqok3ox9N2usq6
Rv84HOSYIvUpFb35+vF2MMXs+4Ds0pvnT6NK4FGS5He4rMfRIo38ocPRk1gBs2v3IW8MZXHqZKQ0
xN2gR7yY+lX5jciWwKXxe/XOeVaBuGJWGZFHvNtKO1sjW9gYmxLNaR3ur1DB3xgUVRFXMtw7OeTf
ly+47D7Zb2K4xPua+0qL3tnhRNpCMOttHGkO6ZL/oDrA2l6rq//SQXmKQjFMMg8upCyYVgQuG/dw
hEkuQ7Ivr+nwQm+1upqZd2hTtfjl7ooiZKupSpJLmEX+qohEk7krB/N0wfDOMI+iOgKcZ4M8Nu/l
ns4sXdD33byCoJQpG8ZxuV7WoxT/4fm5z3b87x6fxdP8iVCoZNsQmqhUEUvNa3XO8clOSDzYIdIU
HXhv3K4LwMmKIwifimeJNdCWGgzins88FDCJclIjyoD2iPg+SST/f+PEk8ZkLtnbg3RrUmQmdy8J
Ee/dbIJANnMqOx4dfw0aruv6q3Jl3LNASmtxe5RjyVPZefZBqHkfyvzvGIbmryLEp0VsrPMQdiA0
lH4hVraiMzn2bgwF3IwpEyw/xAYw2dlqgVkd8ZLWuuEpcDziQIacwtCLJZT+nPFwWogNRcWNbazT
swo5bGAK24HCT878VPJoexvYez0h/8V/6L4bOw6LCqcLIt2W77e4KveA4uIhQiHZFpAxYX3xdJxu
js0mlFEi5/CYHTQIIM60JQk72Vf/mhAqih/0Q3zyK/M3WjNh5kG3etoW9MkZ6NK2w3U20naYj/P0
w0OaMsOAZ9THYZ2lGo8zOgDp/WjJx4fbvwiwhhnUeo88LDRAxtsfWjXDIbt+qW7dyvGJyZ0StF78
5/uy6NBk89cnVeMlB7z1NLvnFJa4VcVBgy3ujLbmv/RyeC5jr/2r4h1A2+Mfhh0cZrYTGoABKaHC
LdzAvC5FjvHuxmBLFGsULbGRhYXy2w+sntFDMcX4UGqN7mPtBwyDlgXhtT6nxK6HZ3BrRJ3aD8se
efgO51S12Kj3WzKsCFw/6L9c4B+QE+taJFklLjGYij3YeTV030+2Pseua96finFkstNxsWlCG8s1
NSuKAR/ujSEUmK++4t4a3Ip7s1UrzJbDFI5HHGiKLldyZxl8Yn387PGrZN+ZWuTevDc6hFRTwa1x
UusIsTqVFycLuwIMyuA7riGCIrSMhjt7PbUVvRe68O1HNORgZCZEdbio3d2p6Tjn7SWkrUS2Azw9
0IxPHI58RwhONE8GibVrwdTBBfmrkdyObXSPkZjJXTh8lF9tPcDMzo0cFcxGr/QPJd1kn3qWb0ZG
Xvc6qmmbX0BVCP6jQRQTjOoj8AVelB3dvt+2MiNcDE78+ZwQDAerj1OnZvb4Y5qxutJb1Ikxgvs1
1K1vWfAv5PdBmOBCVsFBn7+3h+W0kheMztJCJFMmrax7jW4YQyVbWWDjtOosTvNoSE5dn9mUJnLL
2vJCPM5oPRTT5Ei3jGvWn6/78MB/e0HDV5naZSq4hhYstc4kq3Ayd3WllRHRyMJqzCPX6UL4LCAQ
Ib9y5dBPLgMWNZ9RNCYTgk3KOa6onwj7tCdcA3ASNGoN/4AsoQe5Zb/6f4pLvCPGh5HgaD+7qnR3
POgmpNC8QKvFuRn57sv7SIkDdjlZxPbSpiy42MnkqhVjIMkzit0mf9IRa383J5C2CwXyiH3p2Lmz
SmqoYXRd1DCtke6xsaciohQXQdJ6mSf2gLgajiiQuU1z4s0OpMOBCgBPfmj6Aryf1uBQS4XW+Z0X
WYhekUCdBYuUY6XZrXi23qK55+4UmKlyhe6+pN05jS98OP4mfO5wqpT6H3zNVz8+evFYxFHMSEjc
1dzPSYvXEVTtbgsynxO3yvWR+QrJ61GI7Snqw21aeB/KgNgMhl7Zu0nnofxWIbXMce7v1yRSYQ6o
+lO8PTT9C8ajgEhvzlZ84B+s3YPvbA/D3wwroEWWWBzPGyoEA2tEX2CD3smbWtjxlMqN9OmCOpx9
3986bXTUjFeynJm5Bg8wUIEhnQHf2kiDQzvllGQk6zxk3YOJI4Jzg2ac84uKWyDdKPRocOoogRAO
+Yz6N2mWynTQLt0NiGPxvMsAdXj9Ql5ccEDhMdMkSEaU3wf8jHeuFRLDjZLi0Rnl05xPnJUXPAFC
VbiYTx4et/agvn4KjSNYIHWR1QzcUraQm9YVJ95zKuUyAhBIJMkZlcVIvi6S9B/iLFAe4fTWg5wV
Hr0fwqeM+26ZWUvqfWugCj3wHRdgkLGYfQ7TORjBD5TABB+xi6E2wkFTPb1DyHnrobgVQxCB9Hgr
exyx4XsgfJ2qZiiMLUyBRfQQCaH5/aBS0zyNoIpK0e7XmltUOzg72DfN4It3PJ1b32kRWBxMfG9v
sNb9JKgFNAVvSCRgK0uxLCtE0hFWyu6OpuQBo/kOnc7QjEr5lPP3lBBzbP9nxRQ6m8Cgsytwgfsd
sl1ygdESRK+fo9F9RWVObL93bB2WaojJG/Al290oduGKJ2bSX/RrreyrUrJVvr1SmaLYbyzf+Yyt
dr3UJ1Kmkl9fz6prOq7SR+oIXCTd9Q+JS2u8JRw8ezI/3haTvIOyQvROnqg0DG9Eh28U0T4VSEuZ
lXs5v3At36yNrXZG+q6TczLmv9X/RbHHcFsIPzG8VdbtKpa0yvlEJupa+UDoZ/Kn8S+voiGsqvUK
+aH4p5q8pQ/APzUlIyminuw1yJR4Lqdi+umJWgWnz7VCGNktApj50ugfXIzhLOfVdzpsYmuMY6fb
Oow1bStwES8SLEob/26qGcPdpF8HIn//8Cw6c7jNXS3ATxNGOjFJvS6jI6qXHjOaYuR2caIJAtar
BwVgOfABptCSto4UMuM34Ko9VTUhI6aE/Gu9cWA5EK6ktpPx4kfARvmEvJFgIbc+gEiU+YQHkqzJ
3o7EZ10wjNp4SI1qHEC7WD9/6BNSsFKn/Z9E8D74fLnJTae9eVMItzeG+az1x5JyaBJU/a+VmE0H
6Q+akG22Z8VNdZ9GNs0tFrqOQwFpLlOxKw+jn88kUTH5hRV143wK4VtDGUADfuRDKhr9qki+iVjB
Vgrz3d4coYrbgS80urIQyRdlLVKanAbcIwh117dOVWPlyHCw8vBacs+PDugp7uAVd7MuTZRi5OrS
AYdN5109TrTCpCCas83/fKEpNSYuSKxACkRnPzrKtGcZHi8bk0MdhY747VBePkW6Hozyh2rOtHIi
LzRMY8JFkHo0t4WdUTe2+ApBZ3Ga11fZrGZOWewevVp08OMfVrSqRfBpkNIU3errNkRX03CV/IBp
2/+6eaD1VtgEnWGsMYQd1UpT5EzqYyIdGeNMIfyXRwEpAGSpYBL5BM9cdnEzfd40ZrRfraDBr7b8
9Ol/ZV8PNSwv58cENxwRGZgI6DHr64WibuYClCJEKnFyjP+kevKUT3iwsr6l3KnwGypWH4FKXzNG
AsPN1tD4v9dTQPgInzHCUjAPwvjupInJ3xG7irbNbEZgLjiaeBEkXuvQllbkHHQdU3SGKNe4wCx9
X9SnVYMzcs9+LMAZm24PjxQqcmVeWMIYhaj0Z04FzdagMN82Fc68+sdoUpCkaeUC0re3Gf5osLcC
CsCdUS4gQ5xYiTzWFCnoPVoMwKBcG3fA/VEwDUPOJ6lz4R0SSCLsyiEbVmUcJdfGqEmo1pIGs/p+
FuJ1Ir1Y7qdfafTrnPHc3KsuDer6RuHvefG/dugiynfAvoH1DiIVdCM3jV48VlJvB8NYA8wV/llM
4CyrnXTlgIgyPgTS+fGb553AKkjhP5512Lo1tPUvUevl8tszebHcV4sHJVVx2TEsm9spXcP8MaGa
vBZFAUJuZkO7i9I0k3FpZBN3DyBc13qkQR8PloPiI6k5A1d97aiMjjZSxNGywLZV2jtWbL1+DEvk
cFKpDfJCIb2lCDnrGW4AdSYraSTIcD1w8dacHYRGY7GmpzG1EvbhYyAYghSEFvc2lKsBvRQakJOC
CtfD1KYyVLh+L9ZgmjnkBre5Vv00TxHYZMzKInKCYFFttbMfnIhtObrpjECPPxV2y70t++t9b/EC
TF6C0GVOi2uibs/FrwT4i/p2EeLYlnFcBirHb1iM0bsF848zIfNZIETK9YwnAmzfHvDGSvgsfr5D
KhcR/PQYGDFDvMXlfwCo2VWF5iiNE6jARCGi4PziNBDsFTEH7fairR1aaYnjpTDM8c4pFQxDJnNX
V9AZHmlFlzXZ7xj24oMteQg8NFWm3/I9p2Y/VIHhBr+2Xuua5hb8vhH/jNmOMogiWA4gtaYJMnnr
XDUY4dXYgHyYhgCc5SSxMKZvFTpyx+ATq24rAriY/3iN7Ue/FLrIJAcA1cKMkqk1Yg6eXx6/khgz
66WGdWhkWirmTRNtXtb3eaV/aPSM2fVLiLkk8/8vimS1ooekgBoe2gS4zsG/MM3v7cWbQsz8mdfe
98tcVc1X8JKVDP4jIc0ue7iVYUGHS0ILnXDAZBkW5mCpyZHOJuVcShmmRcVjNa4ZbxviRL9Bah4/
PnNazV4NdE3SmrclbOym5dGKfxBvA0njsnDGP9TPjq4Biiv+OwpfAMg17OLTS567TParzaYbGmDr
uoku9Tmf4C50tFuuItLKmfpet/hn+APAXNNAJwbnE6S9MoUIK5QDFwbObznbfRuGUAga+Tj100Vd
MTGHrw/NUfLhpQO31hU8uPUkKunC1yrrn9eX7BJrR69CHkWNMQvtaCJ2VXztMnemxjW3kxQf0oXA
lW3Xx9Ew8NmqWUDSkC2fddDIdsMD3Mu1td61r9i5m5w8eBff+BG4Fl1wrEtUmVwhWiln5AJXvrn/
+YwtXp7a8sPZrebpKt7Kndr5meLT9x/+utgyHpQCYkM08rQT4neItdu5Iokpg4qytHqhopfRpPEc
pqSMYK4M6266D6/286/1/CWfLjcYH0Y8KxCtz24DaDWj5g2XOKIM6ym9zUXkquUlhqzqJR3HLzSL
uiT1Ttp+rikF3LwzCkGLe8n9eqhdbli+DdShEBnT3TyxX64Zezf7dZGqabZvXqy7RabA6TWOA8kY
LehsgYysAbmHul+hzucKWiM5tTXcuWQRbH/p4aeqnPlcGocULLuqHTjqxfGPpoacsSFydKIvNfC6
VczUkNsleY6AUs2Eg024XTLp0o7u6ZtF99LuXhqw+iuhHmW4zfXUd0dSUwCTmEtPK9hv+Od7TPee
BWmzxGcVgg9yTJYMuMDo+Ejub6rj42pENSQskYyMtHGhzVMdrv87E3HehhFCXCctFXqGuNLwqmJi
IeVcsKEI2DZxVLaLmXUTJPLzOKv/DI8+ptTgQ65PkDCU5q1w4whKnAtiOL25Wmrzcy21Tv0l8Sq7
S9i4xYkizJ8oPYjCQEWSi5S3F/k0MACy6/CaTzjZdqXi9E9p1ylo2Cyadtf4/6t+MaygsDe69VrG
4nY5YinrrXk8+chYPAAWf9JcUukn8FO89R0sMkUcQ92MOi6RiG8JarPXSPh/Z85Rx418R4PH152B
nwB97M9NGDBuFiPKoYT8TKQbUIVf16TC7yFWszvNKEqIwpyhvk56NfxktQEdoAmpvjAOIqr91pP3
RYNbjE5m11//AuXx8YazIFAMv4n01vASxEq+CfuQg89qHkPTfpJREPYsENsVruQ0Qln8sBP1CuAS
tAsQKWMrwW4sih8OtDVBio7hnhfugF7WVedfpGhtOSaFs9GIoGA2DI8cEQfH9CeHJTsdX/qLb0Uh
60BO8vehT+pxvMv0KJULQ8JyLNHTQB5MlQh5P0mVy6LKfV3tJZ3q4Juh5D1wBUgX1Om6nnk4MmsF
YHAV+5fb+Qpao8/6R4u6cUiSfjgMHyotVd+qvEzSCih38sFM5kN2CYIPjZP5CxEWYWY7lDqDwJF0
Wr31lk2R5DqJsql1H18/B+5wbAUQnjxXGXdjiGs3F9QKyYvYDgi7KVjhJGWiwyTqEGJXxPuNSXMp
SH4PlIDO5WMVjhVN00/qR7GhBpZoMfogAUEaRyuqz6//gzautUQhgDZme2MqlQYpR4dgfCxqg7c6
/EcQNpVY8cvGTRS0TXYqs3693K1y2LlarpC02QbCeTdowWWWz0X9WOZQ9GL4nPGEsQ+5+X0NeYKT
GVQAvbrqc1KsdSuX2ecXjgjKHL/pnnALkEcvPzQE8H2iKkBzTaBU/AfliGMWak7iMkpJo809yGKc
WL67w3K2FYvtabnjqp+QANaqYPk/d57iwMsCZmPwgfSG3is3OuKLpN36UkumV1FBbZwJisfXulMy
NShx6Rfa2m9gplX82M2sW1p8O0j1ovTxT5rzAMRNmR5YvafRmzc1kztGofWj4reCkBqwT1TxtAOr
/TDfzgHb6YbVQpFKI6rXAdVo6eIoimYiVFCeVoubGqvMgwlb78GN1+57l4OUeGYmr4bnYjzYaPrB
eqZcea+q5PER07nTw3u8PbbCT3JmezwbqJle1taLxEe366maDUpyQ2ExtQiBWrYgg2NHe8OE6mur
UYLjGlO1NkZpUZ/GS80/n8601Pjq8Fdi5TPOb/sUcYpVrDOk0YnD6y4Y3gbXwXH0Oiz6V50s4hX2
m3jDhi5oiTCfxBtxclCafpYXY6EkwHRlFg7xnOjQf3WTZN3QuZoA4YcTcKupA+u5SJp2XCyHjHG8
lVVP86CrjQlCwwL3UM4ibPZXRTclKIb0rhUsvqnEmCNo0PokbSmR0uZVTYpzHMNEkfx23ePPfaMf
/ERP+UAJaTOxarrUdzRtA9AQGi3Ki2YdXL5YR27nH5z/jllJG10OMyYVWIYEKmPgSx7qXfV4LfOH
HDrlrA7QkVqaZbps6muMhAuuQkDFOtipVoraVO+DT39slWI8lDlwkxndHJsFfXoOtYVk1nr5+xIb
UhAxarh/QPX5oN575ltvlD8bTFOe0zC+VI5My5mztR95N6MDkmmJFenFK3Q5Nx2JGiNxT3ZEP2Ev
EJ/6MFFJ0/Xz2wajSLxpAQ1ed+vLo3IsGj1y1CUnuzl9kIWxsGuxqHiSXfdON+Q8708HZk+cW9CZ
nDOHZv25FqwrPdzBlcQUr13eAmBNdfxp6vyVmDjn2TI/c4s2fVkLCy1E8C4er1uKGH0rJPVzSVG7
0oUsYrPjJ0Zr/tZMR5Emz0RDRRtuO6epGP5h1QTkj7DxWc80nj2Ek60EoRcJAwAFyXUk8bWe/f2A
epYASigSIsgYPr+NFItShesHiW/aCWgCTWQnyuCqPTv73MOXmpxkAAfpRTdhOeUIEMSZ2OFI2ZF0
pnul2K+H760MPSlsOYzEqOm3w1eTRENEAHws1G6z9LA+RyjnUOisO+plI6goMdBY8vEt+nlBPa1U
bR2ztmWwIeILjnb2rFAINrVLMCxl/D3po4bwK2yUAFvXnvRVlwQQREiGNi+MLHqrT9+9eQseoyxV
SAr4Adf/4F8Ei2AJcHdMa1f80H3Fkh50PL/d93Bx2kZNi6DqqKWh3nTOc4dnjlQo9Z9Kva2lg5sR
iWXnQLZdC5Y7JTg5573ZcoRi6E+LjfMIbfPACCxtCKyty+AMTgRo7kaf1ERkhzx4ZamFKSMSvIVd
GU6CPiZv5dV/TuNJXJRAMIlTF4fBudMBunkaHjv3r//DiyDgh/Wf0c/B4HtoqPfJaxB9cUIaFV/R
edrGFi7VRbc8YOikgCXZqF4H4J58yI4LitKVvrkhfvRqCCh1a8zc5ZGdc6qV3ZA6BcSFCeiXFCMA
AePjWTpfNyBS1aIDpyTCtkvQaud2x3EEU7GSzwH5cgb0FRceTcu5H4HrpO9pMV0dV667ZeTwgSzl
QPtqw81XnHC02R8S9i8lSGm1kAMgUNHi8E9fngJtMn6WSupBh5T1YMV8coIHshnViiHzyRSKtghZ
iEsMIc59jQJrshRWk91/v3x+y+1AIvzkAZa30Mve26/a39cyIzlcQTyYccLIoKH8KuDSLqe/+mxp
CxMAwNMx7qCxuPE/AKW0o3Osr6vlBTFIMID6NfqGtMTTRfIAxuqyCvuqOPZVq6c7dcgUYSqMLCAH
2vEZZ6ekXhHjzVuXKUxrhMHWrNn54rzoaWWxBwZa8S0tZw8tYd4h/2MvgBpqnRiNtYWxc1glWRfX
Bme+cRdUkz2daX4Gc/Ate5k7tDAIRMd+gPARPjRcCndTpMEhJoU63BA5Zvvgt2YIRxKALJDjaAjH
D5S4EFD9NrPlxcvB8Izl6jHS62bN09cpHd7rVbpdoWaxmiXw/8ztmMI8HkFoGtaVKZeXvki6jC9m
zeMstZCHQ5tcuq/fKPCNUXsx2GDzhGwhsjQ2oPoqkEC4mz0vx8WwbUnkE/qCCp6sjY1o90DdqmbJ
KJr9O1eRy+IK3umaD9oup5sKQ4hsW0iFSyF4GFmF9DuTnwOTT0N/jK2GM8nknlY9/Huu8Ci7JACo
vcRNekXfBeifPmCTk4ywtT4JcHgB3cc5nQmuaMWYuD/Q9hC4k6hrndg+PINNmRdENOYqbsGBP6/o
DLe6dUaRVB+SjoI7DrjqJTgMg67FAYcqTvmLBZj5zNhR8SwMieqO0FEnd6d1Zy3NQgEJJx/jAGUg
k+5NUyMg+KIKeivEwzp7x7TDYHCxyXDAvaC5GdNBu5596hjKtUxnylJOiljYyipiKQCmRrzVcI4y
fVM788naOrSn830ECdwocpkheSJuEgm1ir0tYkuI7xV1nRk9he6Geceb8kD+7u2zmiHZwseH94lS
z+S2rhBOjGjPuL9aXZtJw9lXdJAppjFY4LXsN6Joup8C1CQYH6WSOHyFwP4Ft3kZ1MlCW4z0r4wN
xu2GFAeQ7EEZ4uf4VIvM6ctvEfRW4Twf2bZnvlrqUUZXACfrM6G4AglMFKMq5PJ+d5DZSw+H/sx2
at+6HbWOF4N4+WVhQ00PN5TsVohbUWUO6sUJ/rZ02ln+ev3yMp74hjS8xxQkW6F2H8NCD6t+BoFn
dQLJDJ7r6IDS8q3XiXnxQqw8BZ9jBdtpDlFtBAWtFeA/VfkZm/yXwmNF1QzQpI8N6WvShCQUgKJm
qMk8ZyxZyQhgTWBhdo+9Z886JkqJRyqg6xi5OcDrWW+tF9ISVN+lZyhQZO90OI6nNDds+xcCsB43
pLjtvLFRkxq+3G6RyjLF8uQaVl2JbN+R/goZPJf/vIIwEiH5rZlAskuGk4Lu6SPMmjS24fsTXMV3
D7iA/PSL3Su4E324XoIWOvJeXrsWIJn3jST0rPSXOOrSRDM4H4IFgco2W/lycuZcLDr6vI6DuBrI
CbWlK2htdGaQFJ3o6j1bn2qVHmXP9diuLuU5OooRa6oAxIs3eHTVTyXGlnis5RkT0kdsWDqK6++U
3x9JhftWwca5n95U7nMts6zy+JVMdyrqnvTEi3O6USisuy1CtgJxyCyf2X1aLTR/RtF0nSypOdnm
2vQxx4VAPqn+eBfbz6YXIOAobasKidNAtXsazCdT9C1KhsoOeDk04BkLEJxlkHmGZIF18HWhmF8u
F1uVRtNr10tjsJh24JRGkitt1oVdeflMM0+wsqeO0xsAxHTTX1X7jj3RVVygbBWGzHLN9+3Ti3Y8
j0e7D+mwW4kp+cpS4IBUgKgGRepcPEcjCS1/kcc14L5tEl3ZJMlHbZJG2OvZS8SJ/9ewHaVvCi9U
R5+7X+9ml14IpxifXQE7X/f4hQS21RsXOXEYauoGzhvx3HsvM2ycBIQV6F0YhjUM0hUamNOD4mXP
7Hf9IRBiPzGXdTxOMfslk2t3X1/kfCS9W9qrXbHdWc95ut+BuH9CSr506dvK63PWbGTwmvb3RVpg
WJFSVRjGFXSm0diFD+YBUE2hwmt7sjbJHVUaMQsuomSwfFk/p1lyP2Z3dc0lqG0ESxc6nqKF7Xk+
purkowhNSMmWtM8FdMXBn2Ks/taQ/r0nYlSUTX5VNZBtvUhFegSYJw31tQ414qYTaI1Ips9hYWI+
Lg/7bUuAY0dwmlic7SOmpKQyRPYxXm3Y7XI4YmfSJ+ap3njbztOS0NkQ8szXGYbjFHvLJ1YKrT0P
ILT93rDla07rtHpLrVgiP+/Irar645CzCAflda77xt+qLgNu1eZUWP3/6XDZ5bqh2c8vMjYxRCW5
+YR2tvzLYWl0qh2tmw77t/UMU/JX5PmiNhyObAMP4luRqeR4RVdxYfH1voYCvjASEr3GevT6IZTp
TTKqwcsGo63/dQLnH+rEyKVfTRBu0zuchLeFbGyDFcHDLFMlOWQs0n4PzxpunJ5zGSUFrgFIrgzB
ZJTHgayEbXshCbK2yfykGA4dFqqRdvfrGj/0OTvGF/GeNMPAgEUL1Kow8H1HgJ+fmYkMrE1I1AhC
kZXD1ffPXDgyQwmsAXskh+7u+fkk1B/cHDosU1lHf8mRaEVC/Emqaw4XWc05VjYrWvn0QVjaMIYh
tVaD5IS7Bv126x8szJy1qzPK+oeFO5B2RYSqcqGc23+J/SC8cOy5gGlCbGMnllaCj29d6htrMTMa
yugTBfJLflYs9srWsj2UssnkMJLDIzMYhSzvlXFTfABeNHJwmOtiUS3rH7DgVX3+2xbrZzUiRdBD
0HzC1opIy12smA86sHHkr9kmsRosTF3qDtWfKUZLeZT7uNk2cUnr2E8VnMU9BKnqLjSP2M6ei4Z2
mjyru/pUbyhFDPbF5hpL15q8/htF6Qh1fr6AuX4esJjCwBbk/Or1w9dk0LlEv2bPXw0tylAUbfgg
1M8dD3b4VvwjxpPl9ZQMpTwFhMm+1v8AsNsQVzJxlaYgJW5tpuJ7wbBHHBO8/IeOAlAuF9TSATEd
7R7kDYeSHIrMBRkcE4uLY8BecGKCDd7LgP7chWQcInaORvxwxlu3Z0wtkHWqMIZ3gSTQiGkbR0/w
cz3nwc4H5nDJsPY93sPCeuoRx+bSmLUoO1RK98tWRmDxKx9D4mgcYYSSB9MV/A7WnuCjwg9e9TOV
cYNeBJm+BdtkwArgogrVo98OTsLf9PfKYRvnOG4XLN9EhygwufdX/Co9hxquoCJ4Kq5xrWJ5miUl
y24NzNwUlswQXq25gpU30nKjwF2Dd2uUxaYm++wZWskLPrLCg6tcT4XzhOc3K5e/wc3XFODfNvHD
yEafDpZJn2f88RF2rngdFZV3vqskZd8kEadEczrARgB8jUjY1b4KtaIRa1NnF4eq99dIDhoa67/x
z3AxOTpHvHBsnphSfJEHNjlSd3CXiD4p904eBVS9zOO3uXI4yieILGaOglC6dXdpgnJqVDLNojNQ
y5tTVHeP7MI9kyYNP2I/LyAkeWpkjn4/ZGRVMYVL907JFFFEBrt4KsasIKsek/f6jVqIafuYKlzc
f+dnVycwA9DA+G4RMpwdqpajLtpl1KKTztlAi6EQQ7zwuE1qI+6Y5aQRbBmKFQX4N1DSrWI9L0Tq
yXr0pDlvp00JBaR3zm1kzN8eY0DoxieljU67IbUpsZIExc1Y1IFzi1gGWXjbr4JULdyoB8hd7lR7
NCqlKtaRmliEXfO5ksH/xnkSyFJ2qoaWZwG8kkwXbehTtW2AN2PwV19KKfyBFaYMv5R5KIF3MVUr
rGK3cqdiHZJqWCHg0u1Wd8GJzP0FQR/kr9LKg5B5kdkPaz2veNw8MzZsrtFETKkn40o7I4uxqmsc
bBPbXJHqRIIKthLreWVLr/lvyIBb3iYCKrFTSfKPSM4QB6JxWOOtcyu+Mn4/Tlvem3+YXnRPGzwQ
qvChqFlZGlnYihZlju+VJdKymy8AC0DtEzjBzkeLDaitcT6udEk3haHXWm3TttWZaer7jn9FIqvn
Me6yRA0CImXi3QlI9QpY0lZlCX6SqjZnTZzXeT4qaRl5we3XhYql8UlEehjNgYQE4u9t/mpfbEDT
rzSdB85d5ATRuFVyL2uDw9EZxs1xSNPpc318KqTiK1gQ4Xi6qZ2GAzka9JbyBH3epJGJR9t8s8SG
IUupRBir+nWzjw6t5lVeHnya58Pmw5+Va/eQwEWD7J21w4n2rnG2dsQv1iQpdrEFt622v/9t63wA
9HVthGgTX7LYKe/kIg803YOg1LDjhuXwQd8dwlllF4BMs79gEBDcUhnTrmn4sh7yAGpd6AgZihkI
MN4OMgGYcLKWINY1rx5343kQ1kBKO6I60SGdfKhS8iy/UCpoAdggae52o/3x0e+XHZYVm6Io1sPF
MKY1hB5RzBzWJEtX36J1OqYvCCtlWg6LO/XkaK/Af6DmtPYmirIMI/b/E1/3JI3/P6v+aRKN44Js
nsgffVs8sSdPB6ZRxRTaK2AVH7GTu+n9IIJOQFLYgld7Cmt5NKa4iPGDzqrUKh1EpR3aprI53ArZ
guVCjwKXpeoHnpQLKxjyW0TPpMYLx2v5fFaIDKJ/YqGQgdODkz48kiPjkbEGl7evBvZoVeY10mJK
/gbRUnBmIwRm5ssMbACMCB0YFOW1YG8IicLxkZgBvFEPmBOttRKJvrM4Dcl1keUWpIUgfz+csxsC
HxeAQjhT1NIsE8cOGRaFsNnl3VkCWel+lXvFWkIiJfyrIKWxNSHGiXAwHmnsQKdwxY8qjuTQHy1j
2Xrgswg4QAel7rlF8N2IV7aIyJ1qPoHAdJp109MvAws++2NZc5q8/aUYM8bITMLVDsZNEXU7OoBx
D/L5X6dgOkg+VubpMigVDXifPJJnYS/QUV3ZOnIHs8WqKDPARSvSZ/JsTf4Vw9nGXkCdUHXSLf8a
rQwHO+CxO+SBwiI2mZ8X4wZ8FludI8ucRRece4m7ANMt0M3ZLF/2IgUcQxn501dFjbf1JzNMFWhv
VZHFtI7ZFyfVerXqtDgqJOTG2eh7dolIGBmAvYP5GwU9g+cmXldGtmX/L0NSf0rnRR6h/vwuZK0z
Lj4P0xg4VKvCc7ipVqUoxMOjBICWYLbuLEFgGp3BUZCAUcitJ25m61HmHYUTAf5kBUVYuKps7JKF
Hd9wrodO4HPAi8fmOqeTWob/7sqZYXCY8l6ZJFitKOoM3k9w/AmO1F1hFpEFRW65kMSx+sHpcReB
/4WPogZhtPvvOeKp+2+aiCW4MdE2dCwP6BGMx5Ck48b1JWBYEokt4JXVU8MJWYCtnayj5aeilsXq
76vNWGM8w9ci9copwIqWhCTcdzdZW2ed1ISiTnGz+ruFiZ3hmWiWRepcAT9RgEyJSN++Ht5dDHHy
7PLbuz7g7X7nHyPq8HoWAe56JQsrMMi1yZvFXb8JRfJxb2HN8llnoseLGCW38sDeqBq6cZ2eizPo
F3LT8xYGrStbXjUHLvlSVgUrTRsN7MKVPUZ9Rg8ICbTtFwDsAbKsOzhlsK4VqTKd1qyAg/xCrWs/
IynInz9OYob4/N+G0cg6NIuBGhTVegyRnVe6Gfkf4k6chXLrkW2YQOSPwEsppqYdZO/33mqtJ/fy
j6Y0Ecxikrtml7O5IQy1SUMDtn55h277l7YMv5VYezdBKUoHr/5FyQVVBEeEeaJ/3cmcMZxsWD69
xVwbzLJMJyzF2EZ+1iztvNgdQhmjIclJonCgfv5Jmakkf8KMucDGO/mvb63mrSh7ksC9PA3lpmOe
9tHnhQ/QYVHHpn9GAqQp/hH1ERNm58eKnciCVzkrek87avjxueNL3jX2SqwxBs3T9QrveFEbWLl+
pkAkWQOt4Baw3hP0kC6BSVUXMtTIeeDuPI4ZzO+FmamNR+OC17CPbi+G8BTjLie+fuLMqNtf2H5I
f7ZKmzRadoFN8Ey3hhjVHDGkdmv9DOLRw5nV0wLBMTYHi67XUpPGMG6Iru7NHgrTBS9U/vKYSU25
MmCy9BdxI37oTHNgJE/j1oObmUWwlZ/5MNSLqJNgoTCsSy3y+UBKpA/eTx0NIu79KRUOWtlQlPtt
7Xpvc9QGwhi7YfCAtJGMiruEk/BuARRH0R3lNH21mxIFCPExJG+XFogPq7+TEGKhqKvC40u8PC/E
XySqKaeQd5oVHW+7LGPDbIsyKDSvEpM1Wt2SEJigazX8fetEK3aTElO7OgKBop3uun6t/q80waLA
N4BLaL8hJxGf3qIsqO5UprM9LL0XnXuf8Xy2qCD27TTN1t7rvDZqXDC/FzIZd9jwcm5RGAiKu63b
sn2varYSckopBX38j43/INZXwdcSx48c4TxuyyYjVBXcZBOWaCJo62qzNXE/0D+ViSuqOWjnEXIW
0bFrqdlq/cmZ4qXIO5ftyw5YlHfQdB6EY1YZdkchvzsUYyV7hTGljrtb5vtgXcX6kq1ZN4/8MJj7
i+XN+JaLlWblEQiZIKLmV5MkgpAYvi6NkPSTP4L1IWyOnePbc/ogxtw00tecr0GrXKg+6V4kVy5H
2ejkraU8LH5d3SFF46zrYVE16AWh4uBJOaQviTmjZUTk8o7oJdbmarRzxptQ5sJiD6BHcCj7F4yb
a05urY76d4SfOGKg92fWsn86S2DWSGph5Lit2CbxEaomyHXpmb8fwEtZHc0qCkZCLtqnS3QqwwLN
KI3CXNKp2bzxyRh0bYfOh44nT7R1vJ7yydeZPs0lYkPzT02v10Fl+y5TKBvGuwUs1pj2+w0odh8h
r4z/vmvLipF250n3hhS+EquB4NZbmnUJ1dDKLzJuD+Pk4B3wdUVbQVIoxRhX4GFzlUveURV0RORZ
Jas4N4EClQnKfN8HM8ar/EDbu/4stRzhhvtsJCIVasDuNvqcVumno0UunZY628BVO2DcUIO7Wnd7
GtBdVtIz52ReK6kE+ATKyT+YtVHA54lR8+4TVuyo16XsH2DJ7XeXM7zFOlRVyfeGhXQb2L6M52Eg
KXe+VEeXyohq56oxMjExdjsXY24Pj2qbJ86xCJYW9CaPkZCAn5eeu0dqvkKCWk1RJ4UaVaUxBh54
zRyrNXgsFsr5Z5fvacB0BTnMVfubwExireWTMf1t+M8f0EvEVaxyKd+uVgswq6+dapv9XoprrF1S
BFtq6h5WFDjYC6YM7BrSvnkanDvStXTabJIP0NbS3S717tTojSZV6KxoXeiFPU5AFUpkcdLYAZ9d
zng3OkK1lMFU+WNdv25SLQVstyFDuA8P0ivN9sekg23pRTQjmeiTUEEO13WBDwjOqp2WksXhsku4
tKeYRkvnBUvmN6mEmprgeBiuowr2MgZA38S48egkeG5ckwa7jPgcNR/vgvXS00JlHfas5m4lN918
NIcsroQZPendPxjL0l/XvulW/2pVWMK/SDWn5YATyO0sR72280tf/Nd1+uxJVpZccKV5xaxHfPsl
PA2zwCWmyELlBDrW+e7SV58fADaKTPLbww+rSwzTfUeX6zILIzFsGGZDtw6iBR9zMTFhgqu3I2el
CiTR2pmphB3EAVu/l/NfvHqzEmSjl6STYFDoBIZEhwwBkzLGlJ5Xvv26kDflgIGctXSvc7Q0QaVE
Ie5n91vCutHl2OaFmJZ+5CJs8h1RObnL9D6rReog6zd1ziyp/GN17dfn6qKL+myTGCvPw/vQrZL9
LicgOyRDJyyKCLwYkJ+pIh9JQ61f8SUz+ewuSGTr40pjwVVMY74wO+TFZ1qEPzrkQ+qBwbKFY2Os
oDsXJEvPHIN1Luvr5/jXXl745bwGkYIfaZHwY8HB8/Ry0AxGvDp+gOgxdePDlFHZpIX1d7hhleLU
E4g6E4BAQcNPGPlXISkn3+LIe81t7mBWyDkQPpPerrVjnIZoe56NdBDPnaZhzdzpy24JkLjPaNuq
Iugauawz2Y2JSJBUCMxDaURheygSCUsaTcrOVEq89ULrTFIXRfWhUIHKdX2uDOGDr/tFXdQkknv6
MqvDUOWwsd4xKYZkbaHt0erFwlOJpQie9nEbwoGHxrtv59ftfOhd31+XMT+jFf3HQSVDZFXHHr4I
/nteaP6TV0z7PJFoKddJdkuzsktIPsYbgTGhjQwc/nAHLjE5lhL6EhP/e2sWAXX7qqFkLTPjzdnc
NdwXWvf7DGM7DFivgSKZhnlmKq5rLqbHNQCLlDM0OxPJJAiIM4E+DyOACXv3+KV1v1B1Rrti4+pJ
4EUWYdk9fbLcuR0LsgTZQjd3oDbN8uCyPccoFLlRt+Cm6GMpQGZMk0f6ucTKdhl8At2zom74yVBv
Sx4vdGAAbmk1a20nyl9yUKZDz3eq8oFbOSlNvcFvXmZSDdmBQdSR1zrvlS3d89YlEg4Uo++kdGi2
BPHrT3u6XDnXEGkImXiRO/n5cPg1nngxkro1/GOMwY/1qnFQtWBq1Brmj21vKflGFmkYnaFKUefN
+RXMIZ5+1g+Bo2/6wfi+qjYTf6uXkscViqmq+38fpGBW2sCAMeNBnGrPwQv9YZ6Qymh9i8hOMQna
STpOGdO+R/3ktSGSRHaWK1VS3Q4mIooZu8J30ToUOLVkKHED745Cb7p8wyg8H1x26mDMpEWy7Xrz
IYSyqu+//ClxdYsT++BsIsvAIWc6vp0JrLDgvrXd7HGogELUMiAIJHv4kFFIKNQz2x0UQ+t+Ei6w
agu0Oy0TUX4G1ardLgxAsq/C6Md+0RzMuojKpVwHkS08dp04FIa5VX+7fFZX+bcA+9gEOpLd+IxD
TqffU5F9xyxZ5cA0/fZNhp9kuTExxuyzaN2z+pPKC+g4QaWh2JAnadKLDp1ue64fmyUzYavSjo4U
9PMvx25wxLbBTP1rUFp2xkg9SlUUDKa7W1hKbf+3jFtzTUf7wxTtGh9/xrZxl5xz5xxn1cIb4TAh
R0o+Ur2IJ6e6t4scwlthLvsUFsUCltBGn3m3yN+agqox7VWddEsMb9gTHmRexsYCwNO4fceMW1XX
RFpFMczviw9VXkAK+t9A+D3HqVPKfJ9S+F5kyYzuui+qswQzIV+xybrY3FzwYAzPKp8wSvhuzOG3
s7iPrDl373VprbHyUAVsCDbyWOjZYzxgzyKeMMMgir1PPzecPbVFLVdZhu+Q4ft3i/UXEpAkiR/I
cHnxXNLGpPhmkGYQ+ieGAGHHdEk+s/BxAT9Tz4K42Yfg8j8p8i0nh4PVfgCSc7U6dbSbkVy72lhS
pCoetLIQw5nHuflbjyHdisShlu8dJR7mrfPj11wcHXRNqFzcLYmJi/PrlAd5RhDMjxLdwIeY8LZh
MCLNzO4BZSqgoipgT4zdDSJDKvLYN0UtR3chfOvktXL7Mm4eWN1peLub1BrOOoBsoUEI2Mqr0xzG
vGO3HeiHshAUrgwoP9qpcmmG2lbJIFPXqRifkztIBEh3bxpcLgFLV/158aidoPoeairUyTNboMFR
sxBt8Q3tzy1ZN6RusUkQljR3fsXa0DCCA1j6A7m9tLPsdJRDr8N8E70e8pOFBMiQv50tbPhfMmbc
QVYqjWMzW/runb3GAtA95SRmCfGRoC1Wa1clCIxg84KwWBV4gGsal774yv7lHql80ANcY9TZoGk8
4Ff2XGuCpY2UTwXGmCkdOf+eZNueaZHybVL7cLcpmFNTah3YTfdnl58CWBLIJaaIBAVIVRNq2+fg
oTZISQtq4zsvmT6wwW4IT0/iuilnosSuCcD+ky4b4wV/6fr1qPdNPAkc7gFh8plJmoG+4dSxYaoG
qULhEMskorG2SD9sFJuP27Y/C91NfxvvPshdSoHjlde++pvceEDuPEuhT/XrNOzQRzDfHxSpiBnh
A4SHpoLEMhqiqF7nplpCxHXZBdgyCW5KJ5TCiArNabtD1LbQNWlRc+reP9MhQ5RscWeZZa5/OJ0C
4AoY6j/H6Wkr8pEbGU/7AmAcXcxfwgXAuc1SvUx5nQwYf+72hG44eUZvD5Cc13Uk5krQ4LzrwFGP
TBqa8318sOp2OHsoWfaL6yzkQ5kOFqLQjduLtw9Bau76SN5/X0hPh7hnTkPyWfDIfIC0gf0wOhpG
6LGZVSHNKI0McFA9Pv5S2EbD4v61fhTjpa0UM6Q0J1px0FDHwdL8qjkDufJQabt8MqXJcb8z8S6A
O2RG7Bg++ik7mIlY+UJp42XwTCV9s+z8JsbtUvb52Wwyl701/F9YojD2B5VuKdMQMwUCKXhCqjiu
5+xpNxp7tlHCktST3O/WC/BJZEoztRj771aJtD1eqmxz2N3VwbPuA5okDC+ftQNEszPigMoK5/gv
5so/gKedgdwgCgaO7UUv4LnufO1n9ScDskboaC03bSwLNyQvEKUA0S+Q+JKfbucyUwBftTTzsYSt
Y1/HlCzaTG0+DRmOWxt797LM/mwI7C4B2qeSEy0V9pPz3DPwaJnD9HHTNEZ6bsoqbVYjvrbYXjjp
t+3eXIOUqNlpIKzxDOojEaLC9+1loVNqAkNZkaBu0jvUiwkLoWdQCAtL8+I72/qcTnONV7ZyqVQL
YVs2s3almx/6parnOkdMrm2WxIFARZuuttVFwxPQ6FNREt4o6QoJ+DQAzPMLPoR7gBt/HUNfi73n
YOH3TWqS5PkNfOV+zFDTlncB+ftZYFC5JiPIA61BUd3ecp6B3p60Uk34QV1r/sYVGaP9XoZx9Y5B
t2lWlV+rnOn37rTk6j/2Cmls5PIAzkU3b54EdJAwCYbeFKWjnMx4lpWY3KVr31G87lL0Qnj6wbMp
iMRYvCDSYUSf4s5bOY7+6125H0BSjxIIJKsMjrYhU0r2ZyiZYcT8/dKVHZ6sr6EZ666WyztJ+gOL
3qF/ep08SsNpjU0HBXUB56bsF0dIiFOm5cpJGQmWrJ02SScJS+TwwroGJZ9RO9/z9vo8ryYdIQAi
R5HcZNRJ/uIBbFLXT43sIo61qtjTaI6oF+ztU6vw/M9ZKNVFXb4MlAaRF1q01tMD8e0rrv76pwXO
WvgKfFVBLD+fYbkAwYcNtx4XHeROI4TC8+d3RkQAYmZZqdUivmMPCnhbtBptj5dljx5+mXLWJnI0
bNZWA+LnzgqrW+L/KbdI08yUooHtP4ez8P5OAQ5qxyRy3OVhuEe02KnTvcqQOMSAF4uMY0tayVR3
2Et+h0PajDTwSnoTiQN/FB14PwvTOe/5+q5AbNHjVUjkqZSo35mJNnH41aE/zJWlLgmhFgojzcZf
DJsbxns0cTZe53xgs1LLaoVm0QsQVXS0jKJFEpxy9GOA03trajNsNJERfhxq1+PkZRWLIAKyykqo
/LlbvdhkDmVwKBLl/r2oDgrS5VEVR/7N/0Oaq8biNVDRMNlyIZLLH112MLrDzKVCNqS+1Nr5aa6J
YY6Fa1pdn7kvQeFFl82DC3jeUBd0hydgq1D1PYBdeu3VmVf3pLT5ZQ7YXfuWQjDsBTWfhUNcVUem
aRfup0jQpTS/xPY8gld0uX4Hkb2oBHyClsBvEKoYdO79LqXsLic5gX3LkM52fFLvDPno0CvTZMhL
ZCBbQilHS22aFHIlalQRYTF9CYiwbBnZ3uh2CBvZd7wo46X+ehvmglYo4U3o8w26N9Zp/nbXnRjE
Oi5mTf3B4kb0akAvyskyKeAZRhtkhUQ0cwwH9roV9lr3pyKz2WvwncMJLBJqCCQ+zhk4uwbwLrfD
vDnOMgY9h6AfcUiPAauV3+/x/IUOySfDlSPZ/ne4+dqvKuVwX7FAX6kini6B10+YuqSS0fM5eg4x
c4ga6gfiJvnSSq3qWnaC+/qq2NRoZK1UcOsB9EP757kLqL2npS54zKQO6lbzYAYf/LeplaTdlYSO
Jf4ayRffReS4hN3cslHI+jm5DfgJD8klpVGmysVQkVQeErjL2Lcrq+Ti+QU05EioJxqrSBmaL9ik
UawBhcXQICnTm4ZZPvQaeiljFyK9bitxsh0RzPTkoO33iMGwZHnsTZT8JzaLCCUK4SCMBNG1LqE7
SckETEHol2bTtZNOQOkMQ4q9thWVIDv1mdIciho21fL517dl23z2cRKSd20zuGYupxLYxWdR9FA/
hGUY3zB6YTUAs6hyln1vwjUvqDMAFGto/Q+pKOLRcFCyzCUltrF3dp3Dr9N7D+WFJEzS/1DAYFVt
mSb3V77P1nGzkD4ozcZdatLbkt/+ZY89yYK17giDuN+d4Py/PnQeE1AXyBHj4PtMznqqslhSBjEg
2+telVvz7JBgRO1JIxmE3gW9UYf5TSDd3d7Ov1AhVM0WO/F5IfEyRzLPxlXu6qyP12+Fh9MyUJXF
xJXis7n4dQKWp70pXpcnqolFxV3v1OX3J4mlIq3MyNL7ETM54sV6dsiJYPg9xdQxcOFoqNopHP4j
bQlOqnE/3RMab+CtcUGynKXL9UseT76D8uHOZ1cCwgzS2Gbox4m9dlf1piUS7IZ+FjfAICqamuG6
CVY8dnZhQc2KkzwMI8Zf25eWCqZC1U9TsXIgacOYupRbL7s0InRrrdVDhPWw9Nl5tl59otLz/HJo
GGIIrybdH9dDpXxJk6mqTuefALZlGt6r327V3rbm2fUy05vsfQVhvzcmfPAVPJPi5Ey3LSkEkwCu
yQsumEz8RrOkr65H7Y4tU68RoWeVTtBx/gnC5lXxcjjRKl0uODvIDixKaQFMyaPmgtj+kfkTGBje
viaCM+rZOqYBzBT2C9btp+z2uBVXcuKdtkTvCR2f0N5rBUlpLr7IuUfMU8wzC7ucneiFUZbeO7GN
V+pIZLn652W0r1ANC76JeaF9G5hCv7xNSNUcioKBxII5eDQzMp8ZUI+dMzBdfgfMykFLqiOiV7mF
nVd98UVJacaqSsw5g+S5XlJDwWoqYPMl7CtYZXlS08EoB6NgRPHY35j0Cd2pbL4xD5oOESK5+xgk
K82KbAle1IAPak6oz7uLWx2zbDuhwq3BoyFXY/BrdpI/OZIt+C/cO17sQfaGyML8R5zDnv5YFMTk
JDuJmWSYO1MTY/X26X5iF11tb7hMqd9LwSTqpHEVLFccvbKesmxP5bd96dEdShl/Lv55TirNrDpL
Ci8RTt1nPCmZVzwnrUGZ8/hprsptd1KhIYcPHGwQHB6QkrUdCeMTfOzNsUugWWw571nfWln3jBta
ivowrYclKpdOoyST5ZrwLh2NcOvdb8lbULMF7gkld0D8C+fG+aRTMeVu61hnHFJ+3aBUivwiTRZz
bvq0f/DL8iV0GFIOoatuZaOO1+EjbMN468a/xqAd4QvLM1V6Yy9sldXQ3UZh+wKoI9RtBSaWpj9m
9RnHu5L3P6GgIwU2wtzIo1fkaavezceLpL/L996c7p50IM+3BQODAxispG5skZgyOazAPu2yW8kh
6oPBj4wJXaripcqPA0ODmXtn9gjx2kNLGJjRzA15epqBCvwT7tFjX62i2WEyXhM21bli9pBh8Wg1
vYmHt3YJG4WIspaJaUYbI5mkhinY2TAA4zyq4Uz3dhMr0qYE9V6+iOenG6E5BvFdbaFcD0TSVCJ9
I53i+ycCnuPn1ZQj7dsBlF5HmPg8pmJ6piqqFTOoNBFHFWGrORsBJNapYwWqDXsfvEuc8ONYJGiB
GV9G3fl9HxSf8nkb+xfyY6pa85xQCYoSNITa4YmAJElrr87h/TLMAPHQ9XH51FGdpcOjjQoVLy/r
LAs8pAdcMmpavkJdoGEaMe71EWeQB4oYh485/avHXQMu5G8bDzCgvJX2pZnyfyQLT9Z1emtf09GO
PYh/G6KP9usQ4CIYONX7uSvVwjsHAnSF/vADk6KUEr9lKKwxBskGA2RIMElVodY1731T1vHD1MG+
YJGl2GMLpbhBsEQswQkMindRLIAZvVh7buDMS0ULD/1MeylQJTpmIoiptq1x0BoieoLppAbDEBZj
eyq0wJHCZ2Ieg+mpUNwZOjr6AS4CTy1UVGE06I/5A/rsXxy1Z1bmVzRZMSUlBdofMBt7TfbIcw0u
QB+0cEr7xpuyucBthQjDpyhoy7HyyNY1y+HEgqMQeOhcPqh5trwTQecyToruUvVVDIQGNpewxfHw
h0k6Rv+9cZMhLDS/VSEQsb6mDqLpXixQp29ix1wr9/luPhcJMxDZiCue+5q4PQeVAV5XrZafIh2o
b3tmhN/o/n+8Ysh727/9uOq0REFvoK+YWI5Kt2OEB+sX367WVuU7U388OA/iqrIWRu7k0we4Amx5
v/2L66yoORzXHwEMHATMI8BRW/4rGqDpuSpPzACezk3Ch8EeNc3kQAIPsx2mS57yYMRYg2cxLTC9
kW48cDChkTdJDLiTWVRX0y0PXJy81DFLXVkP+5sIVV16aevmKKQuLmX9DgJFzs9G/dbeEBRHhnII
CgVnQcPpLSBqLC1ZwTIaL6gzXYta1WaSts1VizzzQ0RFT4eSmQQm6XEsXdw8tslh/1ZCpAiegUAv
ZGdjQEt2UL9pHwLtWFOJiv+n254VOf6uleLAmwtIcmdDrKTYKNf62s+TRlpxQ9Bw9bOd45zOCD2K
pNlPi83oLt3sLcip8d1ZtYk72LvKow0D1EQAspVBG6hF1kQ2D7lHpkZfejJmycSMq6dtlfMHx0vr
y/TlTPvjrl/I+ly8Q7h3KrQDdL6IGgUi6TchnFK3q3U5Fzzbf//E43SAj8xHQbRLhnlMSItBFDl/
ult/gJIo34+3dHxoEqczzw3rA3+o3O0KhtM4vz2mV8NAmwOB+Eatd5pQ9NepRKqykmw6Cb0hAtjC
fAJxCuWin1Ffhd6cltY+rWdDkiL6Crj5t+4trorf2p93Hb4gZZ5mWgU3TzUzXK/XjBXrONW5hXkm
ZnEd1ar+sV4NKDN7aGnJwAIDwJhI0JjNBt0AMpLRrssoPtBHHzOkhZVn+RbmZo5+fcynTQ/R2Id6
KzSJe8f9EdP6QLAHy39xGzVwqwdnUZhmPzeeRtH8Xn16Gj4acKv+4IHxt+2E8cbXoTlzWoAtI4tx
9/zASBlbBKSvKhbSwZWPBvWSQ/ZIshtkkm32pUlzBSrVuFDnGmGtHxjA2P28El3TEjsgRqLK0Ix6
Y8Z77FEWMkeaQdiRgRwPxurOT3VOjnYlNYAt+N5cNhfttstwxdXF3nnLgXBiNhla/YTmIriTii4I
pCF4xf/5pF5VQeVGwB30Nm48hVw/+uUsz8WkcEvNIMyCcsNQlgqGRrN+cK/cuhVyIU8u43qw5YaQ
S7t4U20Cj3A2s38NtaM4PHsvbMNNWTCrPtbG3Pcv4hKZwGxHPpWd3WpQ80nfgDDMELcF7gzOYW0h
d1esyqLP61H5IY+bZgfRYiYZrsw5aBUcFrGy01DMTS/qy5iDiJE0/y/2wkECUBdP7yINxjnriyPb
7LY9eMs=
`protect end_protected
