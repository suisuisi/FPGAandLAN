`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R/8klGaE4rNh9MmCYuX/Iy4tnSar9y/DvgV0TXyRlBt9IRZHelFA67K+DNrfMVt0hQWYPzDPDK/8
hhTYXcgdog==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZvVrjbQ7D8uRXx/5e1R0+OcxXV88iVdf0pqBD9Knitx91Tg//TSUXrypu3RlMAA5cHZRKupVzRG2
gLrg+FPEH/sgL2GFocpUgOVPO8fyhrOEbwc7uoI155NkBeTp5PWJozWpLh+Yr1Sgp2aJhVtSgpYj
YFDXa/dt9kjTALZaIf4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HMvoHCd6MwP8Zy2lgNIVJjb4pXIOo2sqTbNp4dDZKqJPCqlFYKs3n08l6Q+4mkHxf5U2LfKI+mRB
4Z07LcZ3n9SV8/0qRhR44llTnmXJEvdwDcaQAOKGaF2xLL3rG2Y4TG674zgBbyeA83xopNDaLNrC
w38QNySdL/pxlzAVYgaw1NJSAxE+mQDzcQX8IG3bM91yWjc3OkViU98nzlYDiPwWcDOhpYq5y30P
dywTnWePsX1WYsppCwDfIAAiJJfbJu/j4S20rWiudH5evf4IDn5iWnEQHB8pbLPwHZYkk8a8tz5F
WsGgL6AJXdxxuP6fUJorkAAOzB8zCi7Jv6njbA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D/iXIWDsgbYOLrw9tTn7AqkXSZS1S6X7c0WPnuuSvZZZszI4k2zv/uqXadj0ziTR0fRUMcBrTgW3
/0cqsCjfy2broeHqze9cef2iPy/xfTuuFeL4/1hyCegKvwG/ilIGXcFXcONfCIpNJTiiLemAHx+U
/zx7fhP1N584mSnXGsY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u/IvMvG2nCOkwNyaSTeTlfkSkdhWkrKtOOsnX/cnnmCpNqVaq+x5AgWSYo98Cl05zmiglhAsHKsh
FGaPM38pSULjSSkj8teY2eZJ6lIi7Ouc6Z6Nz8ERJHTGsXnW11HQOK1467Z1tlji7EM4INEJqMkv
x4BJc1l3L0KHl4DXDdOiMpPrUQGeEnetvsz7ahn1JZorG1yaVayzjyMUl21P8/wvrQLVUq2M/+Lm
x4+c7ChAlzlPBvXBei1gmwIj7L0Brc8O/MHp2LdIOvnhfbSAdr+j1PsWawlTi6124oEA/4rbmUqM
laQ6qzxFVDBWAdjND0PX4GfgU3VfLuMptGifDg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vkm2u6bKaw5cE1gJILxPQNDT/0Ayar9EVnKG4+nwarO2pVND1GaI7yYgOpErI2H7L2PxiF+T/lzA
m1ckuj7lnTN9/B0TJMG0hhSc609tITg+nRIhl1vC9o1Zp1/ikQcx/TqmHfAkdiGjmUAuvPi7H71q
1IYLAzE8L6PvTKIFvUwxzlD3whVgpk8QMqiFY5X5HNpQAkwX1Heip2jpHwctRixCED9YpguUg1UH
giBUYyTQ6BTCGM7DVPXx/2mRtHF9ZJ7+T27SDomiQRDeLNxaLGn+ij+vwDwzzNd8d5TBWMc52qvp
6c5HTxW6mh8KQEiDUxBXBarfDoLcLMAaP8IjGQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6768)
`protect data_block
ng+hTw5QCzw6rCTGKSyFSDjt0bCrqHuFe3qE9SqXT7bC2FWggejeeEU00FzFlQS6MEnCB2aR2HNx
9J1JLQnD8INwzdIYyXNny2Flxh4cycHCsF7/quEZP3sGm8IeO4GScWM2A0Nc9B1UGAHKQbY28jzG
YPDNVFe3qx8ZvHbCtVaILtleG/l1+Fx4Mk7ROFuScKfUuor6ZeQ48ynPruGXF009zhS8a3+9iMVM
YqYCZfLTYfJuiFPUrq2OVXOqPWM2j4yPFoZfYVEBOhToonQXW1uBYSTCF1kM94DdcIFptRNY9KLh
AL9EuUDBXR9JM2lY/V/hPZGE5igUIoI9686cyqb/1JMIKQNIHQitYJSxvXjeADN0tKwrgpaKpwpT
r0tsKjLjrOQVY4f9vuOkoSbeeFfyRperopUIfAUrB+KyBMnLeM4k6RHlZoqcwvvX6PiuqVL6IYla
CUcXMuWuMpL/dNmkCO0cbm6BwODqT4LwCsSEmgqZY5R9pCc2asVuiHbddyiZwUVg4WCmPVPsAW4r
KUZyshIazmN7dZ2z64U325wP0XfrwwHdgJktxpWqkWn1h31mG18JCWduMFxJsAB/bBKSXSJX0vTN
SaQvw1gAEuO/X4p5QjCysSA1X0k5PxN+XuQ31w78D+Zdgxjghb/CQChTqpQYWfxEDT3RXPITg+nO
C4sDktFgtjMEbH492d9tEg1sx2BAtpCPQAzA68EOOdA3E5w4ya7qQ4504hF7roblTekmfFpDvwjd
YH9mIMbvD0hKxoCxwnAy3OZuEuLnDpKYcGv3gVfpehP6tigNRB5Em8W+7DCP0qjeqhB42Ug4EQQD
zSnwG9ik7hS4DnjlQk9MvaqJrfcGJxqOp9nW4XFcBNXaqz1157GmjoT+XjSGiBb4TwdPMdRowtWk
wwj2aw+EvGeCZDV9rRkk3D+AnhT2SZicAWtOI6fbvBGvW+KLP11GX4EUAdGfC5fYdQ+iutjxYq+Z
dAGP+Jp98IDJpZ+WD5YMRb/gcWVFIJapaKQs2cPPRqH9OA7VMfCpT7NrLEPFAhnhvj/1LA/tn+3M
/dQ1nW7swryH9jIIvzAdQqXtyinxz02OJPKIHC2zcuVxPyqbDCGcBPKlOx7UT1RGnfyiRKqTmMeS
N5LvCA2cScOHDjwbxu0JXiz1HAVn41dE7F2Y87/Wlwq9pvbydnu0+NMHQIekUQRfvMZ4A4cMXbB4
VbbNK5T8vJClfuuXB3P+st5V3d9uzAm1yZDIqSFj34u2flKS5fd/G01K/BjcQTF12Aq/chjZgVjU
rNXqPJsJH8Jda1G1wN431I3/UdycVt3VEYsh4LJHJmO2PLkF4ISt9prd3x/co7nfw4EVu4Y91Oja
DvsyKp7/qZMZ14ok3wurMYXrSw+mxw/Fz1XUSlU9VSB7r6h7hWgfVVRqgflt9VJkHaUThyS+GQjG
pfJQHRb2BpoHQ2UWT/CLpcByNpk6YJKnbGTqKOJk+haZ+tG7/RimiOgA983y82ujhckYbK90luLk
jiRPDCGvKGYp6q1ZrYUiQKhSriC0zf91C0CNGV2VMEtgejMaRQt8vF4dHLZGKta6Dxks7XFoJcKd
uSgH+7+wjQ3sJEvEdbyX0W3x57vGeuXOB26vpjjYz9imXLhcMfnlGJe6ZSKG5WEiJesGKrSCazU4
WHKGY2OsJi0pAeX/Uk4X4UjmJKAdW4Hn35xVqawODpnXwTsPjV3qcZsCQ47GMA+DEO9sfYuMpTPd
7KXSjZdb0uBNCb42hW/CihdyedfG5D5ago4tUTxbTappklY22ayUTevBrFeA7HMmbT/oqqsIfVx5
nUE3fD60RPF5Frwyy08v7wRjrk/iqOQegZ+c/gOtz00R5nWT/8LGYdZ6LdB2SOJHmZXfDlZLkZEd
rJhJoNqs9BqxGtu/G7dThONk2cguzRIwYzDkxeKmdsJOe6jWb9z59EyPQlrynXqGobqn5bkb0aLY
eN/qdk3/hBkJhVY3PJbwsGfY6t8B8BPJ8Hmu4KQMg+vhgTqHeUY1IyELCDYeUtjMS57nXYPYGyK3
Kg1JeQ/qR63MjIusD/hyWH/9IRXkFUkTWPNgL256qpqRbcx+SpSDKkTe81rCR5e00zHm1KQNOMqK
XsN3T0X0x9l6W2unyhnqrKbxipI4Sg3f3Sn5QK11smQkCCqao07l+B0f36PMZDZ30UKD7qHwabsW
E0rAv/LMwlApW+a4LJLIz1EHTEjbxOhx6PV2905a9UMN7nW0hqljk+Jd4nqkJogUvXlKLRKTScOW
ry56kkwPA4KBHTZpA8dWQhGPzWPFZ/FEDfc/2kZ3gD6zQ1IUjoA+l1b7wVATfE9FpopBEbt8wjak
p+hsuVtbkiyEbTMaC/SA6PblOm8/w2AW06QqzfwplWOlY5O/e5+fnEzYPOLuvRVeodWyJB4q+txb
zrM4lSpj0un/CvggnhtVMsIqbdA0Ux8V20LFmsPya8W3JLdSLzF/7S0t7ViqyG5m1Hh/9Kl4QUAp
I6/uV0T80qr85cWTeAZWBFJpNZWwcJZklz/y8IV+xlGb2/j/sVgkN3wLBfFh+D+KTmRUkBnhHYsy
QE96zNHPlh7ury5abffuywlcZFPUd2j2YjclhULdhJgg9YdDuUe0u1tbz1Ma1Io1Oh/8oRwSIYmN
gAKyKza2js9oLUlNdqciIBXMubkD+wEQrzj+cyxD20m6xvq/gg9/Qv+i6JO87dPYGrqWaDDJk41B
Xf4sYY0gdkXfImiE+IEFOIXEP//igAvTPO4VLHua/CQeL78uTcJf0+k1pJQl4z1oyQXzbREEsmil
DhI3PUY5wob/H4DwthWFygxq7+9GjD12Ec2g/bsyQRS6lz2Hd7s1ZKkvrI9tTv2sBK6xx+yZxFha
LQP9ECGrsARTX1ntcsyQce+f4BkQkiSt4xKPgnKi0xNcLYnK9+cmJGC5GUDseGBKjEeP3sGVLnoO
KP1FVjjhhTrQZN2n16Yp7fVWpVAxzm9PniMT1BJx3BIK/tfTFCojPmRQeUKzhg7LbDTxb2VOHyrH
3Wdqd9M5Nt+1hTPgQ+PcD/MMprqVhDgZ8Y2xz1Pksj8xQ3SsSibL+fIZwEF3N4wXNbF9fTN7FWgo
jdImtX30oOEwf91bDm2L8e7BXrUiVg+MOirE9EjFgIdZPzbyow1g2ZyM2MKBo/Hz5AHUfhnqkhNB
ErtPHGuQJal3W0WakqU0oUDDBlb5+9fvilzEWIscSyvgX5t2UG7VAUqdFqc2ZSiBueIH26cK3Cg8
Y8V5P9FFF8w7gVsseD9jyR9NAmQRVoypTLIt+J3ldNGut1a/D1anvk9d77CU0G/BRoh6CN/wXMss
8CbLRdHw7FC23v2H13NNmmMV1/zlOdF7HWTUP0kf6P4hs342guhFJEHyIhk0AgsOZAyJixkvS8gc
Xe6LJ5+iupNe3otDuYzBTLwJ/e/jVPopeG5RBJpVNN3CN5c3j7ui9ihjji4QHpynxdfGqMC7ri3h
7k2D6O+5nPcA78MHLuEZ41iL4IiR/7CkUMjbznAKfrbOHh0tLaLZzSqmG+Onb35f7aH1CCuQYDQy
TbwaW0WdHBzoFYl3uOHAmaDvx+BEgc6FMRw86PsjrRjeqTM/ScwR7FM6UUgy0o7Sj7ELtqMPfOHE
L2USOBWUbQ7Ho1QzkR1Oeo43yq4q0WjaX6gnyYbnsI0MP8Rrf2ajQj7vHLdEdtzBsNXQzg2mB9ah
9+e+gitigdeHs3NpJ58n0U18rVKI64V/Fb3y76IfxamF5nQ0XdO1ad643HlbrwFJGZhK4jB6lkXM
eeScPzyu9lEhNOIe9hQP1XHWegLNjdyzdOLHXM8MpGpbvOeg7EHH5FilbLLqqNn3DLdkJIK0mGMn
KdMdKxfJLPGTctG4VpBnTKeiCdCANCmDkORt5XQSnlvvxlVfFyiwAwlbsnFJ9Kwll8SDg8y5CVg1
eYfibhaaUjKA3WLwNcPeyOaPZ6iIlDDdcZjuCRs2YmJFuK8BRaY00fFfMU5jtWgcKaACgqa1H9hE
cgYcXCnU4gYIMzRfq4hWn2B6ILf9QH/IxrP3YBkDK+QM5886CTXSr0IZ5vkUQnWxBTiuNQqhiHU7
bnPXzTgXWhlOKMlwK5R43a+UoIQQpzlGKRMorSi2gRH6MaOXFa95QpTDRVmBxD3HI4Xrqm6B97ZQ
zO5HCxDkkD54DzVMN4Oa0+N3b2vdCWjijowNLq2LJ/B6F3QVRz66seaHSeUy/Qy34TMM3dMGSPJV
lU76iMKcjwhQ+YPFr/+EcoGtjsxqtqs+r55VHxCu7LrSDlijhpfd9r5cNi7E9u7peGEmPtKWaF2X
x6C3XBBvWLAQdje45+s6i7Z9idc81PJfSRimLhtIEGQOMb36bHFeXGCd3iBmOX43M3Z5phPJekb6
tvlvq9nXmKQ6AyPie7HOg8FsFmTiVcnzy9JjC1bUpFZVAE5ilEyi9htA/GFeowBc5LSsCcsAzAfi
088rgSUa7XxbZYTIAD/15A8LElYwMlBKdr5UAwemHO7E127zMKmiSz+nX2l7ShhVqrEfzyGVpnO0
YQzFyO1/J5+/gBR3L6MVIOblcPbtE7A3G4GznwRT4wumiGFxu5lvuUYDpGwhAy+/UsZBF7xDONmA
0SoOIN4eWFyT4wV/S8/WPwqt7HTykP8JGmy5mZHPZfq38FU/qQn9B85XfgF/CdyeMixoSsCnSAtg
wkdv4wbeysu5+6hiKYI6kjrVJQiWyBwmJWtfFa3iViuJz1nBXeGs/ZAudUcpOUBP6bUIduJ7Tgs4
457/eaBs0DS0B+eUr+O8WOAMiSmqSEFwgLT+LB4dHhF8xKiNj5BsfYj7kmkcZgH+BQdToSg2FTtK
B7MVSksSJ1yx4HhKghR0eAsGNv3qgLIwx4/7eaoGjbhQ06nZXJ2OmXdULvgFu4b9XtQ2jFq4dHO0
sKbVlK0p0TUpkjqhYhrzFDF3/K6sTzVcCFSu9rqCrwZHJ7wtY5Ge/LsST14w+TjxfYl/BUt7zKd6
OVVn55/zozmFPgkiUKKy6GLEM8mqIxWsHPKAomfOElvLqtf0+C/FLtmwsYFT3hwZa9jbv6W2Unhp
2xdgcT7LH/VLperUCwwMI7HSiW8BE+wZ+1By/2mPyq6KuD9aqd9hyncQSodB5TT+ZKmqR06s5S+G
SAspTobYk7kl0SrOoGxy5xKmMnFc3BRXCYaYLCeEu6PYWWmSekUb15tZ365JIelTkdYNDWFzDHlY
5e5hUfrte0P2lYk8xva/pijM+6N6fWX6sBZNXgF6r4C7QIfU74dfTk6j0ELAwJQcfK9EUEf6z5in
ddsOSqr0JLRvw4QRUA3095aWX8LpTj/PYV5UHppe2VXqu0yzB8+Ym6GDKyErlFfuznWktSHsP+jQ
aJWeEyFcELQHcVm7Ya3txlgE9oZcx47BIADajzgxCyEgL6/1p9bCnAOauc7pIeGcZt/faQRkuYEQ
FboACpCIwMUP8Efp2YFc88YgvAC7EfaKxY8GffC1YAZKbPfTyD4d1qFkuPsB/wXVY1sUdMjfmnUL
e2wX9eJ0WWxIf1wMwiCT/qg/nkP66RIiPPniAJw4bFm5JqJKSDGMk4WptQpVVFdeuo48LTPGd5qS
4+9N3/3qJsE9F0dzQtCYrIhTkTphz1MzorysVZVUQmxyRGYGhAqkBZ/N+oHkhxYeheRSV03mt7yC
mRiNpLmCx8MgqYSmMNyX4sCHOWtU6kAuyZY7AJxIrPh7HSCxVJPOLTv2BAfLLTLwW11U3LRa1d+/
hgS+E+0AG8bw2uITs5D5iF4KrWHIipqkUHRem8dUYh7MEWfZjWTxFe+7JcBo31PtKyRUUKGvDwzx
SdPXmS851ri+TqOP7Cvx9xAsB4GzcJExhHjifOOKxZA6bphJUkdBOXuFvh2JNDEJq8WL9erm79sq
C0QlgOEqPdeWegJLP1u+yYFts2KsTLhFbPVuwZ7NTGei/KWRRbLbaySTIDA5cFLbdcQK0YURNDh4
esg8FAqD9SDMnt6LfOG8pwzE0CMroxlxRAgr1bxJfZfvLvn6e3ROqgKRwTQCVBEb/TL1fI9jqb0Z
4UugMzPDwDgLMijXUGq4iT+NVoL11drNbCM2Ucp6pWJ8NYQ7HWRtyLtbF81iPsA5v3Q1JUvm/HGc
kQagGfAU6A3aJIwG2l8tw0wTM/syhfEm4J7plPd8Ldqwm1aFTR/GgKT0UGaIVcg6I3qkfP527h9i
o0hh/yewj2o9/pl3i/tgMtoPQOijD5xydvD7W+GWpbcqMsYiS8lmgzyfkOjOby1Yj5WXbf6Ui+zE
HXk5nsfOBdtzxYI52bzwlTygC8cuoEAIM0SuGt8/o201PcJJ3WAfoOVxLmC/xQegr+Dnq9LCkZ+0
krb7QlvLPzDxSXQsI5hCzLCO7z17VEraqRodH/AcZHdz5bE37iqQKvTvt9o+AzP7iQZt6kem/18R
ulzBjyUtdWnbIyBzEIIoAxueskMxD4Xu+of9qmsOAQmbonCrS8Afd/ZMA1TN7SlkHRTNrltcz6zp
v3ymHuh7jjOTuNYQVV6Bcx3cLKRNhCUUYg4SDSVG5AwIJ/UjySKlA3kRjshVqMmVpq9fDd0yeR3p
cpsdNqkIgamOmOxaQrSnjcC+VFSBejjTDDYZdCb77OYwLSw60Ta8yMzEDmnTjY5nJDScqiALGjU8
hQX6VsgkDmOPQqvgmbmfaVsKFZjvV+WF3h2/Q5G/iOnW6I3PxlwKphmf615mZcAF0DBuYfdnUhuv
ux7EkY4QQ0G0jBCO/7JVfLLSdztlmFu6T5u5f85RXm5mySSMcMdOCZwdJS4359hFuKo7LbiIplEp
bD313LN/aJYxS1Gy7QsH8yD0Gs4KephiysBrBOgUNUqYxIi9hVF6nfzaxkKHJSyQCt5lmOU5zVhA
/3UQ04mDo8oxmEGztqRAeFeAc6imh+bQBToWywwjGw+bIZCX9Wl7h3nSoV7Hjo3xsgwOxOL1ERiG
UCvc5KRq0rgLyUsqiVWqtn58MRRT57Gfhs3Rfjv8+AqjyKNWaiFV5BH8XcOxMeMY5QqHeW2KHGVD
vtYHchruFMOPoW9ak6gaoDCnAltCEvKXD+UEAIP6WbkvTq0ZCA9RkUzSvT+oBGVE532+PPiyWiNe
+PfeWpdMcbtv+dmUv9XA10pRI4JF/U2PZVc6vTMHdk73YAUwl91WWbo4gVmS+LP3Fw+/HIVToad6
BTqt2ZJHj904QcvTxrbo2cGGzv/NLlKnQIs5kGyaUxN8Dd3mplJrLqW7gs7zAVXtyQ/oiD0CCb/k
YEor0NiZrE1TILDgNt7Y660EeaUf3Gu9z+TdVeR//C/LWasZRmf1R+KJctWLGIkrWTt1Zna79PWR
W2FsGJpYLjC9t9JYRCXvGde1KiY3OgOtiC1UhX/GB+ZJLgnska8Z1GO2IUDTrvocTzzyVMk3K0sn
EM8hAz5Cw/8BzgJqUUGIyLtT3QRPpXzRJw9VHk0KjojRKNbTt50ztSXxmZOVIdg2QnlZVruUdM/a
O+OLNXeZOUiXRvk6R+XUAHyJEoBFtn4FLss7cVFL0DiL3+zFNy22UqXvTascomvPEF1yANkjvFJK
Z6nb0HhX3ulNv16/TKN6VyE8RN59B2kNQIo3GUt0sW51P6DkVKMv0HUxKazvmijdq2TMuQdo19mN
KHMYlzZduIZUAWQxDU8IwgADJkhfQkLOHm7n9ZZVafVuGsZU9P1lhio8cRlK5culg+2UNCEN8g70
6uWos2H1uTcboisgPTF6+DVj/BGKs9aiKHA3SayM5O3noZSX96iv28uC9zZ8OT8TZB8r2Lknwbbb
1JOoLXt3XnoK/OceHtbZQowtHXkF2qACtRosmVK0AvHfMBNnZeGrW38P2torgqEOBreMYhxpida5
++IHvGjjFOIqHVuLsat4aT5uDAB75nkjcILVggxg4x31hGqvyJzLJ72iwNaC3L6UIDHmeDrij7Km
Yyk0YMUbctuOxVBwqO4+iHxot5gxKAkOMqikX/2ilLFbLHbmMvtAiBJitXsaYEW2SXg/7VW8oRpS
q/uRTqZBZm6f354riGEFy641M5j+cOVfX/5awKAMt7KqGLOngjfTs1A4WciadGxU6a1H4udt4RMj
lZ5uqqWP7cK+DMfSsvalSLDllOgpYSeqMAISEYrVpEmwjzKgUrCYFJb4raOsEoeJDyOKy5iubagg
8TfQaTelF9yxnjuH6WI4CWQRenE5Gf8ZeW8cQOtnfiZhuAWDT8OG7gEzOvosYTZKNW3QMWF9nZrY
pFIgnbjxNpjgMfFsndbVG+MTF7CUpFSr1enm5QCH7hKtd4jpLfYKEO86mE66IwmhsCKPoQU0Dlyq
aHA0ZwEq8r7n5dyXmaQmHBvTHxBCa3F4x1FHNzVjrRKkYa1TFwmQQaH3AOsLuyA1W809l0sWgfoS
5Lv3jeEjfaBz7Xlsyas0W9OndAUE5cGzqxCWCwHeVBH8z7j4Kp5Lo13WpNBYrhp9+FDw1Hc3KhLd
YsjjdF4oWIW86EIz3fiaTkRrgNgBjD3XNK1IY8yMg77/FwS61jhAAkxLqjV904Tix2JbWO9f5yjF
gpSMK/HtxFY3LOsp1PMljV9sOnznDiKPJ8vhGK/2vEajlWrdaohTk336f1AzxOPBvDWTSkjMbTj3
3OUUrVj7uzZLxwRMjGP1eD1/leYzsEyXHDd+kGXBCbRNokCdqszBh2bH3aeCqdhT6fFP4WlmXklL
60aw5XUdiNvdK9J757C3CgxcUUOFF+w+Srjul+RnfQy2nOP6os+EkRb3QM/ZQqvaCbaOnn+wKwCw
krfUq9yTTiLS3rF8DFTTsMn5tfs7cOJirh0RjFMUNwoUy6VhphPRel4JUAPEI7m0wabMUPomS5XV
tzdJKGBHOJOtChjZs2Sqad1jT97B9JZX+qCfsgdxTSRBN2J6anbYDGpO9Rk29GNXy9kvyrQNc8at
dLF0E51T7IT7zprkBeCIPidJu1+HKRRCa19zQ0gv0WnB5hMPSfqZUW8C
`protect end_protected
