`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lOovj60F/36/SmS6HGL2YoZqU+R6HMaRWxyFEmNfnbUwXUI63tMlaQSgHxSzSPBQJDg9qS6YEHxY
xHTVdrG0Dw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VRGCd3WQIM/QlAXLFeqeLkJonwLPKfgzsiA+iTNkSyhmnaoeFXllv2y5XznGwnukYc6aq2TmSHpo
sCmaBLCnTkuk6FBvkcKngPCPDvI65AbR8Sp+iSUsBodg7Za/P8WblbA4Sp17AkkdU0US2JwaxCkO
l6aCv6PUhnFHVdonSPE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a5W17eDlPJRf3DEqIhWY4sCFWmuQ8vFQ2TYiMnZdvyW5ti8fsz0fz4Cx+wFf0qqBfp3t4NJLXnTN
/mVV9NqBoCK3X1uMAZTSzpZKJEEURoBzMNOauReFuZlFN8pK3pqCx9noU6ugNyjAqB+Sjo2KQRQV
F8mlKKHAO64izY58gl2ZoeqENV0h9Ak+la5W+rM7V3HWbZjnS40i8OiuPRsFZsLKAw5f7sxbNEKE
mkC+mr16HgsBjCGS3hGodhUlNLAMFC6bbo3rPWk+Sp62LE6Fnkij7hoBJ3cYoebFFuVrmdvRaad0
AWxJusk1cH/brTz+rW/Wx0NAvdrgmGLOswiQzg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/Kf5sf9tZ4xHVzMm9AtacMEqNH/0YNjKEh0GQUyxICblVa3UkBoDtSK8EV9pzxphPSten2yV+Lb
gsOS6km2fKlQ/s/sG2tAjnhJXvU9CNBe7jRykZzpFmqdInRzkEgLQV8wbdL9sKvYEo6Mz/58q4iq
7Fha7KJV0GS0gj/Aekk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qld2FMhlHX+jtBJiVJ8G1TlzDdkfnrRXO/gx0+KIAl2YaV7t/8CzEqAC8ah+OGu+hgXORGYExRAs
NMcIfeX86MCrW/EW883fIdupJAsW1iyUlXBtezbeE9+UzTmM/r/7rAOUIVau08GDoeumvt7Y9X3X
uR6CTceHr5/G83hLgUXKCT0Oi6lSp8027/k2WO628f8Veu3twv6MksloNo2XaIIGKdxYOCr8gCd8
AH84A2lWPMMiUrAse31apCd6vPk72GYY0JjsD+gDCtaHOP68iHCZJ5EwtcfnphfQ45rgK2X3yPlr
iuAlGtmeyBhX7LO5t+pGk+1x6WYxkwcxANCOYA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dXCMxoBFa4HuiNpnO4iJDiL8354Nga0YEylkDCw9SfhrYiiaWYdYIPDUboAq0inT/vEM+bt3/tBt
ept8+U+DPFCJAkX05h2u++Dtao/lE9PB2S/9phDTIqrqc1wFkmRiVir+h1trMVLi4GgU3svUAzo/
O7O7PiW+VNB1oGyQLyDtdnpkAWKs22i0E2HWTjU2jioNImqXCjv9iudNOrSDIE3k0EsgWDO9+Nkv
fq7GAK08JIu3nx17lWLAtHg3JrAtYyyLbcUTeAEcSikaBcQXc6ExpSpaH5f8gshMtb6H+4/LEYwO
GDQNl6AaOOKGwORorQZ8BVGNqtle0GIYQkeXHw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6128)
`protect data_block
SRnPres9zl3dEAaeg53tBC8zkUa6h7OATb0wUDgtOlGgjdVHBgfPzP3e5uryd0lPf3AdtTsgoiQS
chpfiiKBih7dIbLGVCHUuxjFVwr3t0kozcWZMEkNrEzzYMpPWmKNxppLjyeqbeRXC5VZUV0/YavK
mYFO0hYk3DNVq3PFjGyS7C0eDHpJUpI1MOG/5XxmZVo3J3IWKdfHGxqZ6PqXWX3BUEP8e42W/12q
8MqkiLnh7WDioOgQJmuA0XtuJ4btn0XNe6GEtK2+uMZNt28shbbVjAIKjG5qU92Kmqt8pNXdxi6g
kVggnZF71noTRVYMZcQW6kjLr+QDlSGYHoxKGrBx7OnZw5zPnltCuBZcXFbbxyCzWeSfFKeBaLYH
YCWYN78+NnI0/VsurTevz5NgkJ/7s37tJv2qRn26KnhqSinXpkbwuSRNwbaQfQhNwfQFY6LcVHjG
cou/MJzFl4YjC4n4F0EPUHWlGNyU4DSa9TH2fYNmTZcCKGeqikgapoT9PYQoD33tlVRtpy37OP0Z
M7i9Zmpm50msG8KXMJh6YT/8cmNf+wuIKfARzKARqs9+7nQarjB+NC8RYN1G3p32CCucltDdMlQf
oGtssbzeWMQjwjKak0Rugv4iI+/nChugUA7lM0E5nMFcyCmyQoGwy+iPYg1J8sHVteqYlD9qrDCN
dKTtpuYTxs32KU8fSVjvqdlCfH6pkH0YLT/kKt/YaP+2fS+fpjuedT3/amQ7QpVKenWe+7dBu2f7
yIpzvciIyPlQI8oYNAehZ4pJCdEIAR1ltfMuys1jSPA4G44nqnsRrv/XphOZE+UoEL8mWCPY+hbA
+REKkFIncYNUQf9UIpMivCpTHU3n+a4WEfYcAo5SoibsGEwWNoTCRAMxd1ngagNyVaTJ22tdW3Ag
SgNqH5Ci9uvJ8eDLnbfdW9/g0m22eXRQ4m5cYUeoos+FOpIVtNQ5oenULUbHWwof6GGDIgkzerDu
pZS+tMLhL7Zgq4EhujWss36BreWoXukqp/VH/fDc7rBNwBQP6ELotcWBQBtIw4q/rPea4FHr+yr/
JRaVPFzQqLio7k5RwyPkeVGY4SnPSnjObXohFpsVWgwM7MGUO7srFyvCea+jWlN5Vv4xd4fgm+yB
D8/UGupVY8DajsoXiW8cwt83+Vuu4DQsjuwdmzvxTMNjLhTnF2dwjFyfvKYR3AF0hik8JS9TdF4M
swoVr8+0gVOwHfCalhD3RndNzhOvtm5HU/APFZvCEMf1MRIGaAb9TAcmmBBd7fQ+UamuXAeU6JDe
pKSFMzOtPaHVoRoP7jrt6EK4AgmrAomeSRE7PTQMagq9Bsoyrwe/1rWrhDbaKr8GlN/hWIsAYj99
ewFb32MY94fZdYV5UYIXnKdGsNAHI1QtHk2xcnLeVlTY7fVZbpzkIzZmCmNNcsr+CTD9wzKcY7M4
o7UaB+ofqTAuW8uIViPEbhA9StxQnnQVqKHenwq/g2Y4CjIyGTvcM1l4gXHeypkPY1eXJIMO/zoP
g6mgiw89Q3KrmvMhzDGGYllTpHr1LrOvyq9t+wcqxK0Ibr8+lF+/d4NB95HRvgINyNo4lIGwG+U2
AInVjL0A4EwnMHHehjVaLcBbTGOW/b58yU/zfnhXl4ss21z0vM9E6y/aqM+NZTP03dOUrVavtoPe
Jaoy0BrTQ2WXQvyRxZC4WAfe/QWYs/YV+YGPsLIIJ65hUiza5KtNictwkeUkzo9Mqq6hoAr8dbQ/
lnTg4N6x7fH3whtmyaIFldGrcqkLjLry7sPohEug5hVacyMF/jfP1gLHpixbRjOnuyEHkV5obBVT
s0zRPo7DWaP1n7PWDkujEhNqcvOBsuDAd3WjAGdAXFqCgEU2wD/RAqx8T+PuA1bQtAvD3LFXW8FU
GFsk86fOfl50PRlpWhNDVbeeKiuOnylCnzkxW1Qi1mnxkI2ZyJTth9pesfP29CEF/e3XEDnZDmIh
jRdGU3oJzbsh9f1aPuBSJ4em87meE6kSmq/2P1cuOeDVp5W+4lpHXoX3KPXMvlmfOzC/fs/5vp2U
MU4MvN2XpaDTAo+wGio5OPN2U9AtAOX6UQkt/+RXn9tXSE0c4FHabzgrK2xPzLPQrFHM23SrVdvj
6gH80j7EbdruKkyhBPDOfSmQGe/rtHoSOU6j/Cd8e8Y5yyouDhGYEMca5AaceSAL8pp1mqbKiKLc
011H6UC6FeevPyM+DHUZp5N/udyHx12jB+TYI3nvLrW41z1b6UqbBE8yhJQ8S4Gw2FHPCylU/vFg
GZDyaeVqTUj5goGmnojkv/j7XZ/yyFz+2VWFwclbuo91AgYMLGLSqlpN2MWZYm+NiCuPDgZ/5UnL
+fRQGic/baL9ZX4rjfSmHDl+Z5ivoMWRGSdvFcjdvB2jBXjVkcsxJEBN/nT3rPQ3nUSFR1Ga20x2
Opk0OT9jG/odjbdqGDlu9AICmGbhZI6FYcQViyjH563aYLkqLOQdKeI0GJW6NX4bRoJS9k04aJfB
BK76E9xhlrKE0UMtKFlrFpX3M8xZVQBoZiR/rtksSX8h4g4d5iW/tZnCX5MkZpbUclIt2+b1JrBa
xDizUf1QipaM8J+GNblBTnoIhfvRFz71eUeVcBYswVaOGoV5YQu2JnLZrD1iKUnDQ9rSn6BBH3oU
5nfmaW2qka4jH/zU0WQi0R4L+SA5QtmjsMFp7/ltOkD7lkqNlKiBu25iNR1bOkCYyS9Me+I4NAMG
3xgtRlW26xkklyn/Bjrj2jtZ2rjflzdwGm127ZdNa5JWnHydnDBfW6wmLlCK+HZVQhYl6vn6vVdA
jrn7gN4SkZU4h8AE+sJhJwvstI29Y1hQEq8BsGznsmkbNA9vfAdwvXXdP3gSjAfFAM9990iA5Y1v
INYMq9ukvZAkjYMXiOp0LYcsa3GvBj9urGqIvM+G8cUEiTkOjplwNl/GV7Y5biXnncPYXdRCzpD1
E8RKV1Qj0M7ZYSajS7vGoNngeTxF2kdwxYJywhVmZjZGDq+Vl5ZQJDI8Buw6nEcQ0aJFz7C5k8bQ
iN2bLnd97xQqNpGoG8kb439lemz333QMy7r4u7HaCKhRFTUQFbXfHWMn64D/Wlw1FszLryLdw7D6
8Hb8J5k1/Xsx6ot0FTrot9IT1LsyBmUNd9sDVC7lVWpQNvrWJrvvz2M8qEakPyNw49C5zsljMSPV
VDojYdM0ONF6UxyqrhKgO9KieSkgDBxJtYEiGEHPDMofhxtqpOt3gaRhAaOW72zPHLG2/ZzBhpHr
0r6ATWA7xkjtQ9Hm25mn+n2ld6v/lXktkiGeh/e+DnFcHoFElleAi+jdqJtR0/yJd3QI8TDu+2Ea
VVSniBEhcHyvpsCBVf8FiX36LhOFbVeH49BXWYSHoieYjh34SYTccVefB8Yo5RpF148uIVtNorZv
VkazpFL+BmGHYmkPnTUp+3bxdH+110qkKbMTF0DgERoM2ZaSttWBJc1tXCmib9sD2KgE+Maz7dEN
+V8oZWWLyEulXi5X1WYtOmV5dyf84eCJS8vkWQ/eef2ofC2hwTPd4SwGbM1dHzz6s6+ek3XYugfU
VEF8tfUuCwKXZGumHl4QXJYXH+PMyZtCFaAjxv4Ucf2sGrqBz+K2+oq50ZsBzsmicmkvQypV+Kp5
RSHHF20mt3SJADrzmQblsxuC5RQmBaNEQ65n1cdy4EH3DSikV+OQvfetHcbDd3EG5myF6Aq1JJKH
LTBkv8GSEH6p5Iays+2HWqAsto8uZT6mlyOyef/T6xVfKd3b/GcF8s9hU7pzQC1Ow9ELkVpjt8T1
ZGtvM6mbbfWF/bp69y+sjjUwrplM2ENCE9Yes/tKRz7CvF+WGXRfEs34g/3FHm4+H3NXmk6t+/6M
uEVsX06gFVASFjBkatO8m+5NjuDpe+u4LamcF8LThRTpJTsM03xE1pVXyO1NCsoRkpPc0ZRvxz9L
0uMoHDTAuOq6HjZ6F01kF15n3LwYa7QLAl0LEsW2yQqcfmsaT2UqqY454j5VYojJihF5y8H6ijgl
7CeTpntg6Zi2NFaAUcZek3ga05ACGobxIo3MBpWvYKa72PIIBNZt4IvCnOOAh09zrHWdKk5wlRfw
QyzS1/vI2e59xZU5eXme/iFnFxWjZfGDNTe/m6s4/h2nQM40anLZXmMKxoeBm0uhUeWmULIsZIu1
WNe7wOwFuszHtyZjK3W7KkOOpweMxqAaY8r4W2UccvA0/ISBwJy4c+v+mz8JEUlmmN75fPTiI97J
xYO8pSkNJw/qcsAm8n2L3T1RYY8D6D+c05JGBHcLoQiXoMTenpt6HFTZVUrv4ayWl8XmKNH85iWG
yloDyuH3+W70Y9tavIh4VA9bwFQIUAOeLoyCjhVRRjUCGFVIjUXjszjmxyUmCE+gRKzLTwj4M/Ew
9RPH8B4ftyiydguloiwInE8A3+Loq3T7PYdiXwUMf55n2xUmCWMVNCwXaCJt/3fYJlZEOWLNZle7
lNiABbFcJWkAPOH6LLy/BIzNVdhsxdLSuPOZiipjHRcYnsudaIDSgl5+uR/PxbQLe2r74cbK4swG
QQzcFSo5rOtT79Ldhu+JwzBg9m7kyBNcExYOvD96ntx+SGlgeCVUiWnSoJaawln9cPLHOyq5C2mH
S4pzzge9Cvf9rsB/cy5efgPlT7+sc66qPWk/8RAH+yhL1nUxTt5SBzUDxPXEoUsMZ3ey6c+CzEXa
6OirjX0S/UiFoShIqJdcITG+1+Dl5Vp3YBLJByVoUhasaWIYcFfr5gERf2D0yVPQVT9U86zV3P3s
JRNyCY8OnE7/wkNAkV6JCtO4hjAkCFokV+5eW+NKyjyUYWCIu3JbHr2swOkkbGV+7vD5nZAdhmmW
kNo+P0fb0Z3Er/uah7BsmKDpzQBneDAZlea9cXqsWsU0TlCsvfoQkNwv2GMUX5iAW6PL1apexSc/
IEbbHtFWd3JdUJLjWRcS8ImEMGKIh32IotPt2ScKMitydVong6xZ1qZODTLn8+9J+751hplJ4JFF
GYXsYQrnDPMtBNJ9E64jD4khJ1TLC0e1NURqS2YI/PkKlCAYQ3MzwdJ/xToMvuopEfH3gQhsmXaK
8md8T5xNhTUAp0RTXc1gGO+GHOZtx0yjc2J3C/3/Vz8XUIMZECZGE32jYHAT/YtTRntLqO2QDtDa
+DT4ER/0jw48OzcQAFSJpIyG/I1z8CyVQynvpNuRBWCivEB2y/syW0VNkyyhddxPyQx/JdYVQAYt
ODhvxE+1YTuBewOMWReKQK1T09q5wzdifkeoEhCULnCB7o0FeiUFk0SggKYCmRjmcw08eq62mUxg
RJ2oH0uAkZlkjJWXPLBo9XC5cMgeg5kG4jHn+mjwKP+7bzVyEOYFgqrTzSlBiWuUdxs0vG5TZqBE
Cg0DQhqtVJymE3DrbhvovoCZNRJmt+HJcXiHvCzE7spjWxYEmjDNXnyqBZGicLdtHxEz7hF5ULKP
xHetwXvv8PKH7CO7ZkDLGfOA5sBxbnbNto3fKvZChydtiTL5ci2eAgT4ADkAcbb6BDufI+trWqsr
wbR3t6Sl7mJ0NLWZ3rjv2vXKaPjO7jXUX+oAPsmCKT2BxM7ruhxMOQQGPK/YH3RnrrMm+k0RFa7Z
1FoRJxj/BmsjnqPjG9rB6CskJn5JTkA6m2+6swO3ZenTNUbMKAA9fbIze4yDVku1p068pFCm2+0P
+54C1H+sWRQK94c3HnmYY+Hu/T639fW/ZU3luctrNXNa+h+QD1fW+yTsad5+CoPbd9SmE5Po7uZV
UsUMja9gUwg1C6dHR8/YePILWWTlKb8cmD4+sNt+j1iZQL2hLb9SooHEmj/ZoKBrHTVC4NKevvaR
NxgaMRHShXX611Uk3qmpmeCH1ee9S4LKuBFxWmh4+D+Q202jIZ0JRXz71DJPDg1JjZ8TlBjg4kI+
0g7YFRPhze2y7kPWKqYFuKD/vdW9OoEgWzafvMuIPzFCsre4LiSlnx0PMR3ZhEh7Kt9jBsc03lnr
QOqb94733JLF1ft/ZnD5X621PsPGZpKoJH7u1kC1O30sw5F74vwg1/sWJzBFneBZmNsxEoE0VcrJ
JH5GxSSccWVQpYQzpb0wVRQAzuskQnyBkXiSWQA15v1xQ2KADHN1M3hwBxecO23NVkrBqa33rwF4
pkSRt4e/z4KtQRkm1XJoC9KsyiEpkg/F/HPaxaqqpUaO8xLSG6xv3PFRDQegIba5aRTNPGD1bama
VomxMuGXl/1vCZN6nblAh5gC4KgzopZHTa2GFDFeWooxR9dOWwzzXbK7X1C+Del6OSumIbVZxtul
FzRV7spna/LiEchON38fyiclOhRC2sLQQI1WTWvjGTjLwBoYRCALyTZcUDwPo8uzrXtJQyI2Vfoz
llKSxnIqLflPy0H9JMX9g3p3qFsXLmvbKY9MWQSsoZ3rkWpWuArZUk2QTgLlNfiYuLDYb+oWmhSG
YPqIL46BN6P+OCTPphwiD8uObBmvbJLdGyZFCGuMlnSNDMId2y/JimdsYJX31kvaGUNGMuCAvSxb
eTBLY51Mr9rqrtmaM0ywEWupaNexg+cyVCSEEn2l1QqMopA7mG1Vce2LBftjFbZ4Kexpql4KBgeH
EeSyGlRVH7pi6rClMX4qEOi1wujviSjDoTrfZTS/UrM4a+ZNx8nMCd+xQka//1D7I31xj0HeFhLw
gIqUSH1xxmckxVvXYZbc3xuKHTRpmfd8LQXHIXdjaHDaYXFkkdDPL40grqiyg2tfaHLegzDHVScq
WDSN8pOC/H7U5pi75j41o9xFb79b+T0czYjJZEiLw+ny3Hc4GTKxMEe88SsJHxmn9x8v/oql5QaY
3upV0rGqxu5yT7hB2meosMd5DyGWgOKpfh8zstBaq0r0aWNpfP4f52XCFqMpOC91x8Aln4wU1kqH
nJ2nPZpeX76JzBuphUVOy52oXvg/vkl3OOtPpnyIxbx5g01SrJO2IWLm7VSjI84AuUzhWxKd/NJz
AGsXxXPSfqRP4pGL/+K/4KtzSXTRWi2BWvdBf1yVks800HSNggAq54eXuKBZsnfZ17i+b6pdxTjT
oBVFNb36hzs0fk15OOSQy/1RhK7lsFVyDu7MZ108ZyppKCaKKfEd79nLDGU3+T90T83p+o61IUzm
iN0jF7djONqX9lrJ4mUY7KD0I47csCIBOYmG8l3g/jHJA6hktp8B1I6py+jTm+gLu3DL8qqPPq+n
1QerSEHKQB/m0P/oWw90O8qGuZ4eyr6UgRTluMLs+W+ElKNV1TCupEL9MKjjibhyliF6DX5Jfuqt
la7GP0zwKMjf6h5gCtaBHa5Y5AdADCPBhQfCazQQIYd359ltcPPcIxfOjMX6PElAegSnNTPwzUhb
FhiGrCGwPXn1bCu6BEtu5ClgccYTUu5GkCiwBxV6bgR5zTNDMdb84O1W09P9vDW9FbADcViiFaZh
eotq1YDQEb7FdrqGOKFtvxgBf7frWvk/URkZCPbQ2EDAeucNvYOTTKvDbA6bvvPGwsyGGCNGSF80
+X6dC3Zszw/tzk675vaElAXzG9t2mUZWqNMQaA2hoUghDtXV3Ag2XpbzNx+AmgZ/qo9gN1qyIyhP
55/c0eDpuf9JZrDZeM6+KKQxxaTJkniOWpLerKu0qPdOYwg4mwb5TgLw3w5Wn+ShbHKVB69IRXPw
racXajFAwHyZSu7p7Ha5hAFGe2sbgfMyioI6EelAU5HxDsIFl9J8LJblZIn5Sj0bjBWG1ALhWAJW
1dYpEEsIBPMJhX2vH6bTbU9WLh+EmDA/9sykRYRhArDuWyWgkJSVslsmIp0NUx3FaAwe07zv+Zfw
ckomCMXuv8JqVb0v9GHxLuSH5o8pIemCP3h4yuYp9tqVG1QdCPaVIZECBrHdtF6N2e41CUgHC5sw
Fa/gh06qhKkxIf3S1iUkRZOuLIhavB8VRn/SJp8LvuAhvf4c1eqfMJgB0dW4NDSIKEhOlSRnCxMZ
HwQRge41b0TAHYM8PQVWUhOzkQolyC80cIlYHRU4VuNZWko49qFO+16tjQsaYz89s95DqNjEXdbr
GMYkdbKBAf0D/XdYmsQbhNVDOrGPxzRSa0HaRxKX1QVTlefBWUgi2PEs2gg2c4yHO3qfT43VK/gn
Tlb4i2PS1oaqNjNexsGXihv0TlGWOg6VMBAqzQ4=
`protect end_protected
